PK   +��X�2�]  ��    cirkitFile.json�]��6�}�����"���gƵ��Įd*���RQ$ekG�z$u���/�ϴ �vKئxf�N��q�//qI���l_��l�n�,~o���n;�aj>{W������|v��.����}y�nv������k��)����,*.$�%�*ɊL.�Uf+�d\��RŲ2j�/������tFF��́��/8�!_2*B��dT�|����B�9P�!s�"�K�@E����(z�$C8�PI���,��=\�!z�$C8���B<��>4�l_�7�w�M�_�ȶ������X�Cp�P�����������k���ԙ����ʪL
�����|Y/DA�#=��$e�Ge���3���n�H��!����X Ϝ�1Α��{±��[����B�p,��2�cA��!zL'C8�8@\{��˞D��Bb�C0f���4)̂�1��,� Zo���`p݉��eǰ�\����c}eǰ����N`}eǰ����Nb}eǰ����Na}eǰ����Nc}eǰ�����`}eǰ�����b}eǰ��E��]���ò��F���  g������:�@������0������8���c`~� ��Lˏ���o!�gX~����\�^���W8a��c`~�%1��ˏ�����a$�?��t�����>X~��� ?�g?X~���a ���`�10�<���ă�/�G�(��q?8y���	ˏ���I.`���',?����N������X�8���c`~~J���ˏ����\`���,?�秡��N_B~�hWN�ԡOpj��\>sz4��Kn�3�W�ͤ�uf�g���s��2+��Ҽ?a�J��d�+���z����rYe�)}/,mf�k�S	!�Rȧ�}�����oeN��aϏ[A3����L�B]jӿ�	T�s��4�Of�Ҽ?�J����k�L���C��Z{�,<�־?��Z{����Y���,#�6�,ݹ֞��`�˵�D��J��'�/X�q�=Q��ko�D�	��u@@ԟ �O�'��D�	��DA}f(CI��$�W�+�Z�|%Q��(_I��$�Wç"�O����SD�)��Q��?Eԟ"�O�����D�i��4Q��?Mԟ&�O�����D���Q��?Cԟ!���g��n��3D���,Q��?Kԟ%���g[�}n|9�j�����g��?��t �j�b���R�F ��� ��-C�aj�b����F ��`!��-_�aj�b���҆���ڸ����QH]D'X�f���B�
$�8�H��?�DN� �B�
�8�HE��!r������`a�ԕ$,aq���8
�+W��Qz�8�B���8��8��qRW��	�9,������ N��8���!$zI�X���#��a�\�2��a	?Lo�Ws!PÂ~pTװ���\Ú�n�Q�~M�5���@A��\�Z��z�Q�~M�5�#��@��\�����Q�~M�5�?��@���\�ڄ���Q�~M�5�[��I��`�irB��+Q֕(�J�we�HߦI�����D��"}�&�J�6R.��m�,	�H)E<,ҷiҰ[���4�XP��4�X���xX�oӤcI�F�+�a���"^)$a)���E�6MZ��m��"�f!M^��m��"��4yY����xX�oC��x��m��"��4yY��J�xX�o��eI�F�4�a��M��%a����E�6M^��m��#��4yY��ʏxX�oӼ*K�6R��m�2ن�����;��K8P�q__��+(#�:P�ꗱU(._��(2~a]_����hl�E��;�
# e`�󄚌�z��M(Ԉ�XF1�l##�gj9"`0*Z@5��#�⡕E�>"`0*Zr3�$�⡵(�C"`0*��F��b�Q���X`T,0*�����D"�K��%hD�Q�ĨXbT,1*�KL,V+��F�
�b�Q�¨XaT�0*V+��5F��b�Q�ƨXcT�1*�k��5F��b�Q����`Tl0*6���1F��b�Q�Ũ�bTl1*�[���m����6��}�9'8��& �+�	a�
mB���B�F ���&��+�	a�
mB���B�F ���&��+�	a:�ĄH\�ƅmX�f���B:��p��n�(�S�M'X�f� �B:��p��p�(�S�M'X�8�B:��p�qpX�8�B:��p��q��(�S�M'X�8�B:��p��q��CH�B�h�n�- 5Rh�
�)��F�5�H�M���zhT�_Sp�ڄx X��F�5�H�M��zhT�_Sp�ڄx X��F�5�H�M���yhT�_Sp�ڄx X��F�5�H�M��yhT�_Sp�ڄx X��F�5�H�M�>M���Č�Ӥ\I��
m�a��M�v�ɻ�ҕpX�oӤ^I��
m�a��M�~%a+�	�E�6M
��m��&��4iX��B�pX�oӤbI��
m�a��M��%a+�	�E�6MJ��m��&��4iY��B�pX䛅4yY��B�pX�o��eI��
m�a��M�J,M^����"}�&/K�6Vh��m��,	�X�M8,ҷi�$lc�6�Hߦ�˒��ڄ�"}�&/K�6Vh��m��,	�X�M8,ҷi�Ql'ڤ���Ph��20_zB�M:�W�2��&��}4��&e`��B�t����
m�QfSO(�	PH��-ԛRh ���
�)�60-�Rh�0*Z�4��& ���@S
m`0*Z%3��& �b�Q���X����F��b�Q���X`T,1*�K��%hD�Q�ĨXbT,1*�K��F�
�b�Q�¨X�;��F�
�b�Q�¨XcT�1*�k��5F��|�b�Q�ƨXcTl0*6��F��b�Q�=fè�`Tl0*�[��-F��b�Q�=W�������mv�ź�8���ه��9,�6e�ԋ�v����~v��u�K���z)�L��d��ܗJk3+�zYp]J)|�}u;'pa�7X\��*H��'�D�x�b�lR�3R�'�S�X"�D�M� �}G���G�Q�����o�҅z䠼�K�)c���>�&������>Qn��-�#��7n=%��#B�ۺ��	�o&�[�$+���_�K��K�����K7:%�� ���j�:�7�� �!�,iT?�c1������2���[�:x�����l��8�;mD�}���2�Ȃ�m�AdA��� � Ct�aY�!�-0�,�ݶDd�n�"2D���ⴥ5l!�'"|�'P:�i�
*@e� J�8mKA��1��?�HW���(�<L�C��-F��"��^:�i
�h|9 ��1N�MPy�P.�H���m&�< ��b1㴝� �r@�c����� �l9 ���WAX =ύ�у�GMI�Gv�@��l!A�ˠ 	/�m�/�U�?,��������� ���l A<ߠf�?,��F������ ���l�@<ߠ��?,�������� ���l�@<ߠ��?,��F����� ���l�@��  f�e�X�z��$����tnF �����ƶH b|�NG�c[! 1>D�$`��-���Ӓ��S��&x ����P=��T�c; 1>Dg+`������z�K�Ǹ����.E'1`���	������,�0��Ctf�h ��a��94|�K�IMX���RtRf�G ��!:�3�� ���Ԁ�� b|��b�c������0�X�  Ƈ��.`��z�@@����pEe������	U��`��J��`����'�t�~�=��������{���eB��qW��Z���&�N��O�&�N��O��3\{4�?	 �a>��>	�*�p5͔�$ ��e!S*� �J�LL��O�*1\]0�Z>	���p"����$ ���MU��*QP�(�JT%
��*���
�L��
SR�)���$U��*LI��
SR�)�!RQ���JTT%*�U���DEU��*QQ���J�T%j�5U���DMU��*QS���J�T%j�U���DCU��*�P�h�J4�':T%�U���DKU��*�R�h�J��?�g�����s�_ n��������Q���bv;��y��h���i>�sE�,5?�'��i�۴}K�2ߖ��m�U曷��ڲ��[po�[lo����[po����[o!��h�x�-���Bx�-��hS�� ����x�-����Bz�-��P�By�-T{��By�-��P�B{�-����B{���[ho�����[oa����[oaZ�z�-�����z�-�����I���龓Ѷ9z-\ǹ.�p�����W����+��o���CEe��N�1ė�_1�|;%Wv�x�`+��������b}��G��ʦ\6*�9��9~��F�����!R�C*<�O�tx(?��C�t������#�r�Y��y�]�����;�*Xa�ɥs:�W�҈<cR4MQ976����/�͡Y�<v��������.��5�Q��kƲ2gu�u)�eyY.�V��ҋ��>n�F�A�B��wXj�	-�_���wG��ʍe63B6�4%�
Ɩ��F+]75���q�x�cNx�;p��A���ߞ�
)�����~�j��k��u㇈�k] X׻�k�s���m��u_�S�s��_0?���V,k�+�5\�Y��U-���Q�
ю�p����/a���m����g��ڡ��Y׽�}�iN���Y�̱��3���v���s�g�V�Xݶ_������}��}9�{&�	w�D�<��9�����y7�s��/7�;�m���~�h>���ܻy��`�];]�����w�/�?�o��]��g����}S?��,��/���3��w-���J������o�M��q��݇�#��V_��ԟ}o���8�#�g��(ƺ����s���5��W�9���~������/��w/W�=/���I~��g,/Hʹ��Q�y=0ݏTs�..�D�t�,K��1�R�r��cHS�J��.�1טˀ��h�:��E��$1��۞���_o�>��?��߷!��pO"�E�����[��z���r{�*�����93L����T:�I?j�gF�y��L����J�3�4"+gY�*ˬj�=���\�qB�i�J����K#7���g���������s{�y��y=/�v: ��ճ�8`/-��s����쑟m���f໊x{���˾J>��@{���b�^�0��,���s��
=m�/�*�~����p�U��X�Pi�V�P��B�G��J�Yx�E��Qh�%=b��e���A>hÆl�!;d��,Ԑ�����B΅Px>p ��ŀ��e�!�.�,�@;��k�.��m-ڮ���cv3#��H<9���c���qpQ��1^��Et���,N��0Cz�"��H���"����j.l�\�]Ts�vQ�E�E5i�\�]Tsa����f��ڧu�@)3_�6u��z����n���h�ջ7���ٺn?�EU��.�����e��i�xT��eYi^7m����f�F��q|����]�j%�R�ƕ�Q�xV��K���Un��nm����ɼ*�2w�T�̍������,/���]�r����w��3c��e]����gR�:[��,E^Xmܥ�V�	~���x��v�N�����n��ϐ���v�z���L��"�BW����+ɗ�������wǗw����K�����;ە2n��K!r���2����ݡ9g#��vU[����x��\fK�r�Ty!��<�����ύ�k� �y�V�4���m�x���}�y[���-~����W������7�C{쇗?�7.�dsn�|��4�=s��*3:_٥-3Úe��MfUd��fYr��Y=����En��V�8���zɪҩ������A�T&���K�,�˯�4Y!�S��]��^	.Ԡ�\:i7M�\^�ɒ��ta#sL�VM]ڪ~ZeU��ə�ïͦ��_:��<�Ϻ��?���WAB��(�t��H����\J<���V�]�f������>���;��~Ժ��5�#H��}l��o��%��]V����g�������o�������i�'����c���7m��2����z{r?�eb'�m���l���_SRw�M��n��_��w-��7o���#엫W����s������y��.2~q�-����ϕ;����g�����FN���b����L'�m�6���SI�?��ЩҺ�~���Ȗ�6���}c��dYMy��R���״��7;�/3��_$�J���RJ���~��D��?�5e6���Uw)B���!e�3�Gt����Jp@o�J:�/� F�Z�Q�p�\ l�Wu�$���н��/��">"�*��2&�4�2�h�z��d
1���5��&(���_W�e+�Dv��ql��7N�M��=�1O(���y	G,�kl�k�T���Z9t׿���z�y���<6�u��Ń\��_����?���r�|���c��?�{}�eq���WS������4�`��� PK   @��Xw�'<�  �  /   images/0df5ba52-08e8-487a-a0bb-947223afc81d.png�YeTг�%�nda	�E��kI��^b%��K�������.i�F:������9g�3�a��7w��U��qipQPP�d4�I�?����w�U��8.
n((H��0�o��?%5\V��l��p�F����9ٻYY�Xs9��f�Ҡ��~T�����:21�B����l�1*�(WH���bZQ#�,Q�Q���C��T��DA������I��׃q�t�}��1X���PRj$�km@���1qd�j9r��YG��]�~�Y���WX�z=[��5ҵ�� �G�2Ǧ&��PI�c ��p2���*t���7F���3�7!���X �R�Q�n���aI�2v�̩���A����99��}�w�ܦ;9�l>`�E��8�������Yz��a��O��W�q��O����:3(a�{4
�u��Wᵋ&̪���F<{�j��kr���[���mUY��KR�x�P?�%�^T�H�m�^����?�`�D���Fm��H�w�⡂s��&L��B;�Ґ��oԒc�MR\���������![����Mb�'�o^u��O0��'� LP7���9X{^�=��c��m�(SL�clv=���п�-o�I���QRּXI�)��A2�v�����?�jj��G"�Z�\.gۻ�)F}{��J��� RΥ��b�zL(�;1.��>	���Y����^��cD>�A"��f����Sz]w�m��a����8cAeE�ʽ��8�+0��Q�
A��*2�<Q�b0Rz8�$5�9ˣ�U����t��/a���F�$���>��ăU��VD��aa�}>	v��
E��幫������m%���iW�:��	o=�{m��ڜ��X�z��T(�^�xPG1�36WA�h^����aqly���RY�?�����Q�1�LFv/(]��|=��jg��X��\V#s1π��ļ�*�D�]v�o:��K�<h�^�Ә��nO�[��
�X���Ɏ4pc�8K�S�p�[���*�>�;$	j#C�0�'�,I��3gIi��F�U�E�k]wS/c]p�ܜn�:P��8�cn�0�_�ު�T�1�Sa���)ۻG8�,:�e�PQ�ƛ�Pd�:q����B����U{`u�g�`�Oq>29�h�6����%��9�4HO���7�(�_%)#U'b�GY�O�:�9�W�ܥ�7��,�]	��S
�2l��|��z���]���^��^��Xß3����f>�(M�r�|�5�K�&`�|�v���Vz�Ԫ�^m�y^�
��U;�&�����&�U�S�'jϧd��=�ڔřQEh�%�Zfp*q�TTg�`͂��K.]��ǭQ����1���䦭|��&�Y�o�HĈ2�$�ѽ�嘅*�<MJI89���9�ֿˏ�X��͗5�������Q���Pl����}Fn����Y�w����雅&�|*�V��ee\������#`K�7���di�/@�H�ᶗc����� �2f�qp vug��>�V��u$�*H����Қɕ�����n]��5��*�Lb@*~�Q�Ah� V��9`�j{��
��@N<4���p��*0�r�y�J۰�1� �Ef�pZ�4d�f�5�L��F/�V�@�z�.�SLeC1a�H�ڍ�B�������~���ݠ|A�� L�Tx'l*��GG�]�!�3}��+Ղ�[����<�s�<w��4�-F���"w�J�\\�!����Js��x�;�t��e����O^�皈����w�f�d��/8β	{ύ�IXh<Aͧ]�"��[՘��Y��n�?�c��ގ'�����$Q���k�u��J'z�5����'\�/��}M��[!����@��my�w�v,�d8��t���zrH!J��/�8�9ɯ�smdN��<وD�a+E��x�0���8f�����c_����n:c}��4�``b�z�
���b�D�P���L���@j�R��k��q-�O[:?�)��+�MD)����tG�X㾕�D�]��2ڟ�*)�Z�dxy۾���(v4==�,���o[�T���QbE`TfD1�Lfm�p��8��/{;��Ze�u�s4~���ī�������uO��cno��o�OX˙,p"�m~��496lNRU-��go�`�[�G�j��3�az�|1��6 1����t��M�+���s���Sh��5�?O�~'�v!L�n�p|�c���@��ޠԟ�g��P��7�aY��]��"�P���[f_���7H�\'�2�y������pM��d�v��NKѾ���<��$��6E��#�|o�t�7������v�?�N�򕋑)������(��̑�{�K��V������1bM~$�ل�*A+6=�͑u���6@gN�ԑ!��g�"����Nh��b�4��r�5#P�>���g�4�ӛ�q�ַ/B�z�a`o�6<J��*�mt��"6����N���ö_��|q��/g�1��M��l���5f�n�Vs14X�,,�l��F·����S��})�v������Ppy�X�:�N�E����%��&/�i�l�����؝>�~��{�=W]㉞a;2S�1x�G�y�M��|���U6�-�H���]��ơ4<+v4�ae�1e'Z8�Ύ����~ȿ�3M6&��t���$k��
K{tg�X�l��o�!Fd��Ż$	6丌iho��7�����cO�P����J %炏�{ 6��Z����dSk�W�qO|�:U�̇�	�߹N:g<�JO�g�e߁�{��Jݦ��UBD�'������T�������䆘,aI*է���^��Cn�<� Oj��;Қ���bU���/����WE�t�M[aam�����޴QY�v�ɧ��8|~�L��6kI�&�|��݄��ز
�[����4�l�۸��9/o���Q&�ox,bOK!:�ՔzX<c��IB`	����Ѧk�q�����N�|�Ƕ�]|����4�����jx�=���G�݇��_ϐHU'���j|��Sdot>n��Zg7Wl�룳@��n��`.wR�vA�gwRs�m���
�E���~��2UDMjH�2:x�Cӵ����*�9���E����dɐC�S�K,66d�!�1���Xp�qS�#��8����1!^�,�̞�)��+�0GX�`Do��[�w�k���*�Ŀ�v�����o��*��7�R�-���v��gj��e��#Q!~��?yxW����}�����&��֪����CA�U�%O��F���-�E��a���K��Ծi�q�uS�f���G�h>�*�1i���
C��L��&����zz��O�+�/�]}p��m<<�XfRX��'j)QL�3��	������:^tű�q�*�PQ�I�0^B��l"pp@P���,��-Y�죷$�7+���Î���a��SЉ�vb\7���a�#f�.N���e�G��L]��$7��Z�m���2���Y����Xf��^��2�hT���(��O�)�%ԊL��W>,
��&��dm�{�ew�>��� ��e������ǅ�m�qF����{f:���l2�$�vf"kb�C�`&;`%�����"��:��c
by��C��g�����´<�]��~2�o{ ]�/�(u��<*��~ �e5��D��6�ng��}�~�p�D� ��+Z��N�f�>b�F(qGg*շ���s�$n��5/�������Z� ����҉�ٜ¥2���1�E�����pW��,��ߠ���n���[�p�Mx>��f���xd���$P�a�q��Y��{�#���M����oi@LnU�U�b)��՘��_lm��q00tX�z��JU�6��[c8��\r�U}{�y6�awp�P�Q9���eCe�F
xD K&Q�'}!TϦg�����2��o������ٚT�u�G��ő��/"�2�5�F�e2�,Ww4b��e��k-K��7,�BM-s5�/�&d�Kͧ7�\��c���ù��v
�޺�iI�.��Z3��E-'���_����'ٔU���*�� 3�{��!�
��w�L��X��
Ņ�!8xO>]�ԛ@��_o�=<0���%������P�ph�H[��]k�9�:'X��r��l(N�J�l���AQ�Jd�qjQ���YT	�M>��>V'Ts?ܫ�\T�s�H�Ǻ��"vʛ) ibF,�1}�NR ��c�}I�L�C�Z�P��P�MR-?=�qP ʕM��*P�����}5��TG'�9�J��ᐒ��ˢq}V��6܇蓜�C�aT&5��2��Ut���-�#�8�m�؛�)
�|zMP^ݤ�;�+���ZI}�������)�u�,�3{��{uE���6^���p����d'�	n�X�e�~Y�GT�b4y���y��4�@D�e�6b��%����r[hH��7�����4J�67�D� �;���� 
�G�xBm��z�o����8�vp�s^���U�"���!}�%KL��c)d��YЄ�����6�.?G9|��0� ���f���ޜ���u)��ڤ��G,U�:n�T��@4Ck�.��b��#��D
��EA�s�s%(��B6G�s��o�x$�!�!�*eO)Y��N�٧`⛉(>��W�F ��A����M��G�f�+�J��ƥl)~~�g��J2C	vh�n�?0���Y�Z�㢾r��?�5]Ei)�0`1{����u3��O�xF;|xE3��a�w�t�7)!"�R��`x[P�^�]������"2�v��Vd�"���=����i���'<��MQ�Lh�11��Hb8fc�3D�j�,UM��1$�f #�t��1��>��P��|�oZp�����|����Z��@&����\^����j����F��a�+N��aq��%jm�Pt���p,��@���)�)�ʳ��戟6���I�s[s"�E�t=쁮7�{��X_����1������O��I#���k�W!�^���
#�j�c&�Qq�I�ʳP}��C3e~�dZ��E���}LH��	�΃��O`�j��*�MA�߿��"�r�I�CzS�~Y6M�
�7�J����n�*�Y""�3�L��K;�V�(����M{+����)Z�%�Jy�ȣ����T�M��{�ai3�Ǵ"今K�^@����V��(�����/�-@�5���5�a���CD&#�'Zkn��Ԓ�jf�z(�E���o�wH��=�RJ^��������V�9�h�7^Znt7�"/����F�6�o)WlH�*���Vx�3���%>l�W_�@Y��$8N���e�Sw21E52��g]/v�	hy����c$�9{�r-4�7���[zw��:7��7/�c��,e=9L���Eyx���{��ũY�H|h/�
��0]f�(��|�PX;�����zU���w�%�}<IZ��d��0�;�me�z� ��/��̈�2,�n�3����ǟ�ا��:}�E��a��1��*���������,*���cĦ�ȋ�ʩ3������S�T_�l�p=*�UjY�J<SI���p��yZ�5�����W{|�\	✡�o��i����>6�����a�W{��UB�H�C�i�� 0�Eg҆�rԼtf�h�V3	���P ��?����0�D�#V%��0����~@���R���ՠ��b�v����w-|���Y�l�D�@i;� �C�;W�T��c-��H�&Aެ���6[�f*��}�Tj�7/K�S��~������yI@�<�^*�y3���8ա�^�r�\s�w�z�I���&��T2�ۓ����7�����2��`�=^�X�&a'�^��𼓻S�p��/�n��v���ˠT��H�qi��#�l�ŝ��ܰ8��X.gr]i\����E�~��z|���	����l}
N�	����Ki����V���u�hV���^�wv�	����~sCM���
cb.�����"���(����n�ޢ2Ck��l0��5��Bt*n-I��CFR��9�i`���C���,f@��'�C�̲= ��į1�$���Aπ�(�y`��OJdD�q���zO�b�Ot���,��=�-��EO�޹1��qa)�򞑧�)w���ٍI1O�d�##����rcǑy�u$�6����)퍭:F�5��и�|�=��8�դ�^�~�К�!%�IZ�$ �ز�W���52��sm��fx�#.MKw<�ǓwT66����0E\�k2w�r�$%{�p�B|������b�>9��i�nI��j]�K�}0ߍU���[�yTήzM=�y='�� `�ӕI	u`�r*�[�R�I����ߟ|)@Eirx��4 �я39¡ۻ6�.((2�;Ȣ�3kO_~��i�:��e��u<��u��b1���+��V�$�hUh�gB%�B��ߙ��ǧ�6�}4$Y�9j{1*��m��c�@���&��,��u˱K(tqbV(�6��������Υ|���]r��[Wtaq��Z�d��ی� ��9�U��N��,����uy��-���ȸ�����E@5_?b��A��'��eun����}��;� M%�9��k���z�:�h+�̟�w+�-��t]vh��UN}�X�f��P����Xn��UZ�M/�F��fn���9G8Y��PЋK�]�G�oւ~�8;e,�=�>�Y-����3�l�/Q��Y��I0K�mL8�ķ��W�{��^��L�A��&���u��k�:V�k�@	s��2�-�hm�rO�Zܺ�q1�=��`�HkL������=�D￫�#nk��f�7?�ͤ�|���/��6Z ��g�y�1
�ތ���J�_����u���Υe�T�Q|x~�ՙvm���})����H������qڑ,(r��Y�Q�R�>�lrϋ`Sg�}��Z���+���o���ׯ9B��V��2;|=�|���m����0��7��V��d~��]�)��V�˥�0��/4�e�BF�� 3o���C�~��'&�����������=Oѹ�_���<�h�xh9w���A/ٿ�ޚȟ��7�)���ş��G}P(qt-���uB9#�-3i"V_c�"�S�V��%�C�)�����J�V쀵Þ�Є2�If��Qt��]Hn|0��e��r�c��#���5I�L�����Tn�)[�o��]Ჲ��f�X��)b�3q��T�#~��[�*T~�1���=n)7R������ë->�R3>5��(�*S%m�?PK   @��X`�/��1  �P  /   images/4cf22100-3898-4fbb-b8e4-32284cc8d12d.png�zwT����ke�ā�AADz���F�P�B��5�Q�T�P"��@@�@t�^BK"Aj !-�=�o�[��w�u��ho8����9g?ϳ�w����/��� h���!h�$my��V���vI�����KA4�*����8>T
�s����C�U(44T���~A�?ܸ��Der-�!ht��{簬F��١�+��
�폌�TtXjC����ѷ������o���n�щ}��M�^x�}�uWͶ�ߔ��f�Ǵ�;n�~�Q��W��z�4���xŏ�C������W^�MZEǰ�1�{^��9���Yne[7�A� &��{.���u��}[bwI=�"�<n�l�lܨv��~�i#A77o6���ɆL�1����'MR�%j�&����!�4�UF�u���a��U�(��HNU/�"4���`G��dN������z��7T���9��\Č�ق�=eOu�Z	���Rl�ƚlGXYQ)��oVu����k"qz�g9P�4��x�T�ͳ�5!�U��i����#�-s�.�	�n�#�o�P$|Ek웅ĊKoE���K�-;᫞��H���f���0V^Ϟ
���J~��d�5ۙH�^��Qɿ=�Ƕ�%��V�._�|ǽ*?ͩl���-$n)����.mY�3���j�q�0�6��Ŭ儁��HSH$����m�ȥ�Tխ�'9��U���`�J�G���
w�(S/E�4��j��,�/��ˠl�����1��P//+n@�:�TБjgP1y�q�A�m�Zhs�03S��k~ק���SM����~���)ű��ٕi�A�rr������a��Vi�Y�v�iy-L�KTD0��B ,a<g��~oBnr���`[�R�2|�vQ�%��[��f��x�ӳ�/�D]q���;3�P����̿����b���0�jy>i�N����OX%���D��5�Բ���F���SI;s��Mv�qV��.mۘ�/"�,'��ʸ�\h�.C]�����i�ײ�ͼ�P�x�|FeS���K�f��(
� T#'9��(ٚ#uΈ^M��C6��c�?��1�4b���?/��V�*�c�h����x9�Hˈ2�l�1:f�C��ժ	t.�`���8'rVs��ޱ-x�%�X�_��ZA��>x���5i��©LU�
�{}��X|�H�뾒,���%�U�K���s(�������2}����:Z�+
����*s��,
���Yl�$��F�~۹	�2��	v^׮�s�ά���;5���&�0�+"ѥ+rm�ӑ��1�^J$i��1g��1�n���i=�)�T\?�V5�ęU����(��������öfo��dG�%��mmsk�KW�dii.����N���^�5�x�$���5�Hx7Eֵ��<�w	u2YxC=�~��%���F����	��e)�I��~�w�#"[�u;[g�C��z��ZL^4��Z�V��v�w�㬚{{ Q��/��5�p��_gp�0a��9����b�4S$C2^�x'��DbNg��e�w��I<���I����n�p���ˢ��hsl�W����!o��s�����)|�OѢ�t��؛�a��ţ��U��y�>�GzEN!q��\Z1L���|�O�`$�I�BɆ�������{&T����$x�*����V�dڄ5$�M��Dko�tD��)C����!�5ʘ�@aK|�ׇݓo��.�'�񓪮j�1��6|�x�F����G[C��&e�~�]�R��R�l2��};�b{Q��d<:J��Q�}3����mk�
���8���9��<���~��������o1ϊ6C�n�2g�!E>�GsD�?u�mN�|�1;8����jc֭�p�����Kn|�{�3f�<�SD�7�J�jPZI�Sќ%h�ED�M��+똢��[���,���� t| imj��".�_�iܔ������c��㪐J/��ƻ{m%,�̉Hw`n6+�G�:�NJD�t�U}B�0��Z}#ҍ���q޹y(��!H�'s�6�L
^�zc�#���^	�n�Q'���_�+��W�kƌ��cf����,\�����p��N�[�����I���Ss�?ݵN�I�o��I�I������j#ꪸ����&�m�?�y��)g���|�|?:�+���*�/���8�6�?���J4����SS��5���x�N$V�Q��q�!���s�dǒ1%�48����t���J��0Z�PfbvD�Q����M�"bմG�2R��#R^D��+刾E�Um������uA}�I��
�~�Շ��S�u0�u������!��d�n�Q���7����x�|��r�|�ST��kO�d��pf�G����c�'F��adyH+y;]�Q���$F"���o�ܟ�Y�����ck[\;3�*x�X�d��VDVQ��mz��4����A���0����> Ph#M�h�ī����t��[�pQ}���YY�H��EN�����n�p9�l�Q�t�sݦPM'fc�)@bc�R<�@9�?x-e)^
��-e�^�)մ�{���4� ]y1����"2o�@`7���xZ��R^y����olP��_@[I�W�K�y�)ZNx�����^�W�c�(�����Ʈ�'6�Rf����.�o��
�5!�e(:J���׳��VK�;��`�;0�[�x�aҊKG�V��\p���n[����1z	���z���i����/�Vqke0�J!!⮬�r���CJ2	��QNG�E�_J��l@#��^}���C�]�k[�2����6��]隙�x_��`��$�ʿ�\G$�����X�f��I������Lq�H7�>�D9A��-�G�ٺ�g��Zi㣊�� �3�[5�P'I>�ּ-�s��ӯ'$��0�ϓ���quwg�����j|=g��!��iy�bf|�m��/#��f����M��*	�c�-�=�v�_�R�\�@�+ŧӳ#���=���Zq���#{��	o)

��YK3`G%	�<��2	�6(݋���|tߦHs=��L|��N�>9e-�M�&3���4�C_��쭪
-+���rc(�^$?�Ɵ7w��l��$�T:��{�=G����Ҁ��ŝ�Hn�@·[
_w<��]���%�65פ'��oA��1�&�.E@P��#�ed�u,sǚi4G'�����oWL���}r�Ї;w6ut��R���������T�HGC�_�g�����ltԱZ\�>�tHH�Nir���tq���gE�t���~�������/�o�hfn��~VT gj�������Q��m�����������QGY�S5�z͏b��8�흧���QȂ�/r$����|�x�%7��cR:;��O�<�o����C��jb���y��N���B'?t�Ė]]Jq�R�Ħ�`��_�?���+����b��q������;[��ߚ���*�:g��[��(EB��f���dXF�iA_mT�w�ؙ�&~,�p����	^�8a���^��뿽ɥ�X��(�;�`l�-匬�O�X�H*|�������[��~�S�b0�{�g�ϸ����%3˧��wZ�U_�ѵ��df��pE�����K��e�]c��>��N�2e~�B	��,�Z��ב�2�����쮦�K0E�3���/�D2��������/�w���>ы���˾�j֮[:^�����9�~�{f��d��������A�����wj~Y6��-�jlg�[/,���覹�<ԛ�U.��V�t��W�(ڱ�
LyP�N�����H:�`W�?Om^5=Ë�P粤U�
�JŷJ��4¥�)޶TbK饇�⏌��h��ԔR@P���w������k�[oę��R�8;��+Vѣ��?VYG,Q[���ϟ?G�]�啜CU>\��͢5��S	����LϺ��U��uz;a?�Ϩ���L�Is :j���c�SzM����`xDطXJ��J���J�\"�
�
�ʋ�C�#k��FY~��v��k4�p���ƛU�¬v]w�IVV����Wf�/��������t�ʼ;���ã�-;���|	�OXg��r��9^^�d�Ou\�6О\S�=j�.ѻ���B�ط$n�9ԫ�ѝ*���B
������H�ۙ�vmrM�k?�L����[��k�}Q2����i%�����������A����L8&�Kg�f$�4��2n^�'�\]�z��q�ODw����vd�eK��t�ҵ����l����o����)��̋I9�sM�&'�$<�����F6z�.l�|V$s�2Z����u�k[��6�u��ٳ�S"C1h�����_t��A,n����Ξ�R��Wk��<�_����r�y#m��� �:��2^GHq�ձ�y��H*9-9E���:�ʚKM�VH�J\t��N�#Cflo;<ߐ�r��Z��~3�e���i�u�C�+����a�^&��@���c���4�'������nW7hx��I�*�ek�p1�y\ޣ�Zrڥ����SW9�fy�{���#l�	�a���ʍGV�Ը�m��T��jL�O��4f����w`���4���'"���S��B%׵	�j����{���J	O��:'6�|�|*���h	̧��o�c�I}�֥1��*a=�?�#�}7=5�1���f��v���h�0��1��t�_'�5��jd[�^g����N�H%W���D�U��=�=�S6A7�\@�S^��I����X�5�u��.'\�G=���x"��w��n9�|��-j����ʫOfٝ�3Q#�l�9DW��	J�lX�����'�N��7|L���K���)5*��S��蜜����$؛�ܹ6�A'�ezx���Z�m-��z-;�&G-`�A����� ��*�Ls�M�����U�cA7߸��R8�Jyl�B��Cc̺�W�r@���/���G��FKo	�<���? ��N�E��H��E!��V�XZ���<ҏ	\Y��x<j?�n�ˠ�	A1��BZر�y���ň�	Y��<�%	)i�w؉z��B@؉)�����W	5���@�*n��@m�@t��%>pu��Z+��ɐ�����Y�G��t�Z.s�5�I�Þ�/�{%�h���ex�Y���cd��w@�$&'[E��a�*H��fyT~.P��" 3��"e׷��PE��J�eI=�{t�r��'�Z8$.����!�^��Ō4a��&"��d��if/L��h���W���8��9��݂9���0�)(�r׏��?m�v�ݲ��E��_�f԰D.�g�;E�z]��w^
�u�W�'�=0M/D���%����э�v�y5Ń�p�	�'�WVW�Y�R�GF`?�SޖLXP$|�2��%ZWO���C��6����.KKyM����[S��t�];lj�rkm������K�RX�Yʪ�oR���,���Z}�'���RO�ϕ^�I���s�;���.�ai��A�LJ�)����%��[��T��QG��z�)ޗ2�>�c�.�.El�>��;T.��=IaHlfȒX�賌\J%�|�ر2?zi���t��홨��G�����s;��ǉ����d �w��R �DDKaYʨk!R�蚋nM��q�vOI��`�IE��דR�p�X�p���)�-����B �{!<�yƯ�;#�H�aEP�tU>�{�	�i=[n,�n{�0�5��4������Ŗ�8#T���;?<�Q����{P�3h`:l�񢽓ࣝ
��"���J��W|��K����O�!g�9I�^M��s�h/�|c-սz���;"Pc�ia��x‒Zk[W��wQ�fۧ��h=� ȣ��h<���lA7ԱjF5�a�O}�x��@u=��س���@�(W}ҧ�U����?선,��a܈�^��� �J85sc6���[�*�D�nw�1�wow".CMA�q�I��'O�Վ��i��Lt
����h %��M��`���o�N��c"��;� ��:1Y0q���gtw�6X��]ǖ��ɹ���e�g���\�{������+
����2��o��,���9���z3V����VB��sf'��p�L�����b[� �U�iX��u�X�ɓ�+���Q<���O�RY����<P,�>�X�Щou���_��Ck��.KY��ڠ�sM##�X����b�?��yJ	�{`E�/��w���X�D�X�����U��w�{�ck<%4�V
K�י^-E8酿�yȾI�5@Ғ��8�]���R5&
����A -%��bK\�����|�SL���Fe��Wn�c���� �{��+v�1ɝ�2�Sz�/�X���i?>sʲ*+V�/�$*rXK]t�O8vD���X�z&;�7��!���f��.�����k��,ż�lj�\;��x0f�X�+a�{�$��Bҁ �������@	*q��ɤ�t������l�~K�r9�4��*0ˁ� ���%i9�,<���p������[�1��S���^_\21�&���a+��)�y�;��]����(�'?7�R���]��&BL�N��e���K��x�����O8]^]k5V�����U2����N:���չ�yف9k��)H|l�;�H>���%�ef�`Z���9���3�����X7G�����9]ζ�J?�X*�}|&�N�)��7�bvqq@4ڍ���ݤP�����;�j�S ~�@QUUZ�&HV�*�][��u�D_y�@f0�B���'���T�'F?_H�ZX�Y�t�\8��R���u,o��U�p���t���U�cj6���ܖ���V5�1+��C߂i�.%��%����n���E�	�t�[,�s:��'�� e۪fJ�KV�&��Z1R��T�}�Դa^�r����7����҃r�:��X�R3i*��d��vRZ
[g6�Q���5���D����޽����u����6���|�ٲ�G�Q:Z��^�����eC�7Mͱ�a�K� �� ��	x����,\]�r��/�ݪ�9��e,v�����^���R,sY/E5�<lAa�f ��@�u&G�gG,��`O '���ݍ��x��b�~2I���?Q��M}��8e����'۽�J�h�������-!f���*���ˮ�bl�����(��=}�
װN�5��r��l�ky�HHb~8���
A:O.�|+�a��I~�����&��[{��B��u.�3��j��+f<�\և�Ù���έ�G|�yWu
h)I�sO��$Өw��C����;����ѡ�{c���;'����uc�5)��Vs53������\X�y�HZ@������:!�����5v;�L�I6Y�u+�9ft�̦\s��\��잘l�*�T��>�	-���B �����#�&G��>�������v�l̮xR��ǆ����K_Ձ�}+���W�U�������@�NYQ��k�j`E�WZK�1=i��q:RN)n����H�tiJ:P�zᣑ/P�y�G7����u�ER���I�N,E�Geh�/R�~��v�����P�S���h��	����*}��Q� ��I�̉���2u�ku�O�e��6�ͫ�/���I��O���{���Ԍf�ϥ��D�$y6y�G\A0������ӧ��"b<r���^��J������aAu���8H@NZ��+���� �4��Ҥ�ZM�2�K��-���:iR�n�4v@���˽�v��*���o~�0���%б'ݽ�/�[�&�o��������}19s0�+���@YSZ@�E�7��oR��Ջ9$��L�C��f
�'2������6�vxmM�vi�4�������%�H!\sŃ�.��f�M,|B�̶y��}���ie��>�{�.�|y��yـ���
�}�.)��w���������n��ݳq����P������$
�Zᦙ�HOOWR#�Ck��ټ�Pu�]܏3m-�j�9�,��\�]>�_����4���R��(�^,4G'�>15�1��p����\�n����?�y
w��O�a���rכ�G�7��-�?n�%k��-d����L�矒��w��t��y ��� /����3>\��4�����5<������r�o���+�w_sv/�/,,$�v��w�y�\�����/z}{�`���7C�A��w��őQ��R�B����O�U5.�*m��L��N\$M}j��i5�� �k׮�GԖi<�%b?�^�����.��'LMM�Q`ʣ_��˫��K[F�yuȃ�ѡ~����1/iSK��>}�Ժ�;<Mxu�c{;-NNk��#wi���� IÏ�*���T

¶+V�������g�AѬ��N9�F�8:������դ?��&�:l�mh����k,SX�ۧ/���iɽ��7�`��r�jK�̥d;�%v�_ĩ�Pa|�?sͅRр��PTJ��:t֏�@��嵐���$z���RU)w���|�Kr]�k��1v��,"����fP��B_�mM����R��r���ɨWI��T��Vg---�_"E>�K�*{�����i��(7%��`<�{���Ҿ����x�yf�'�O�0���?r�i�:�J��_Gg�C X��-T�ڰ�:/�q���tqk~���a�E�o�˫4�u�~�����d%uV�����z\�sx� ��Pf���SeQʴ>�x��ȣ'qu
��x��iuӣ��u��yt�/Ru;��0Am�[����蝣�(&�|�Ė�zV�'�y3"qwl[������VC��^�.�|�PVy鵵k�"_�~�S�Q���dy!lg~2���A��v]}b޸��D�L��7 Rs����@a�ֈb��Y�)���o�[�o��)C��1��kT�(_o�nn�;J�'u��v<v���Nm���Y���(iDl{U�]9�-ă%	���(48����W~a	���Qתr!��ƌ�8��'��a��/�3g����QC�ݸ�Z���Á��*��<�v�ك�bǢƧ	�͉ւ�V2���f�0^!�V�w ��~�k9��վ��n!K}d��+*��C�p@���L��Y�9b��+� ���)��i9f��rv�.ʔZ�`�3�+�E��l�Jw�^E���R�}�U�)X���:���c���؀3��8�/�`��d��{'�>��b��s�E���˴��V��XB
�͏t�6`fڭ@�M�q~Fz�<���2-V����5;),��K���Z^z��	�sj߱h�Tܝ��P�(����\���$�4x�}F�L�t8����=b*�޿Ֆw�����H��+'''u���à+3++ѥ�-�%��%w�{�'x�V���6<z�r!H={���~���#hgyo03�L-���@��������*�	5_3���:��dL h�O�Ȫ'R"�} g�*(lY5;u��L?m�`z�ժ�N����(<�<�i��XϮ��a��6���^q#�c���,u.E��A����R����;? 	y��sCS��v���k��ʾ��-�Z���9�RNHH���8t�;�G��0�2�^DzBJS��t�k�/��������GX�M�¡Y�ʡ�ȭ�=�E���:����h8���6��>�Z��l~5r(�~@���z(�/��HMi �j���K��̕3�c�w�O�TK�Ǻ�v冗���RPaNmS0��sr6���1��Ws��X����|Z�b��<8c�3B�@�^��M޿Ȥ�R/dG�Ǭ�?9�ә3M��hl�� �or��,���T;���|>�x�"\�\��C!Y�U�l-2����_|{������s'���.��`��*)ͮE�����~;w2xHp�d%!"!{�(�j����DZVا��h��ﶤ�X�-*��������U�a�t#��8�ؤ�ac��A���M��;����?b�P���k��{�2�O�c��J���P�.S�#:�Ԍ�XL���X�^`�]̈���~X�V����M�7=��3QD�Ejǌ�����������Ld�q�C0�D3�ٛ���!I�^薁��9  ��U�2�%pN1�o{~�1�K&�$d��k�m^]�����<Cty�����N������CX^܀!Z����%d�	X�e����4����@��9�S�@��I��7�y岄x�Y�p-��XC�-5ԩ�6r�����zf�3p? CF��G�&�������t�����6 ݳ�a�����/%Le�7����C��D^.�w�9�P����q-a�����+��Y9�\�+�뛱0#6$��M����f�L$� �h�0(��I��g�I� gdU9`���6�3�3�T�}�6�i�z�����YE?j��,���x�I�����N��y 0�	5�K�VaQV�ʠ�(�XRu~Nzhw|���Vlt2�b�J��o:�N�uБlI��s*Ɣ�?_<i�*bn!�2�d"����X�K�m-O>��1PPk��/? W��|�d����ڮ��Y�92)��lڿ{ҿG0��	',5�6{c��vO���\b_�KYf���DN�� ��S�fQ^����oVf<�II$� �T�bK(|��#���sY�¦P[R�Y�*���:f'�Dz�(K��ULx��Eu8ڮ�m�	�l�r���$|.FY�ʪ�n����\_�3��3/�'�V$u�B�M*{@���Y��$`,)����0N�j�
��s;���0�S�`n:Ժ�U�ܮE}�����/~�Y�i�2�d�����I}��V��n�bq�
~�=s�&M���`� �-4�r=]*�</Mb����$�h�uNZ����;9E�]C�&��e�*F�O�]��C脻�Nt�.�Db��D.�S.��Q��k�ǧ�V��,pN0~�N�@����b�I*VBsC��ЕϏ����K� ���Xz��
��dR��L��3M?+�x`�}���׾����C�J�$dΏH`��7.0�!�^Qꤐ|nU�ݲw�L��sC9��Q�;�^�uk�3���:=�/ǝ���Z��m6Έ�|X�-H�7�$��� rg���M/
B7�>�-9;Sw�0û�=�d��HR`�/
�?
�Փ�y�B��{ǆ�R�`�x����=<����fƎ��M���3 ����[4Z���HϟM�y@K\.2q3x����Q����������F��I���EL~��5l=źl����%�I�4ԕ��U`8�z�5w��d�&��S�%Xܳ�Q79}�js�5��h��U�aI�-:y-'����܃D��g�Y�����[�"j�s�|�Gm+��nH5���;D",���9JC���h����Kp���Hm���Ǟ¬��w�mB�����c� ��4[JFrl�e8��͒@�z�r�F�\XR���ӧ��K-$t]�	�P�hiJ�l��u�jz{\)�������q1ۂ�q���c�=�5!t�Е�,���f�ұ�R"�@�"i��_3��氊p��L��Ͻ\] ��t�֧^Z���mP-`����9�a���{l�����v�_�\�~[u7F�`�خ�3�b7�������� %D��;t��xy}�j
.
��Y�.�)$�D��	�s�޳=?��ޓ��M=C�7����F�-���̯)E��)��
�j����R�Y�Z!NE��?j�-�R�����6�� S��ݰ��;1+*83OIV㉹���)�v;g��ˢ� -�`h��al���X���Ě��o~��t�,Rrè����|7B�~^L7�/KV~�YՋY|^�eچ��h�[���`��������^�"���|*��V��l��R�a�W�\�mT[�A����y���ݓ=/��"Mv#�nq[�K�GӴ�Ն/u�������z���J��]ޭW�Z�_��K�6<�M��b�����>�#k�r�y����$8�f�M H%W�dns@?r��D�N�n���R���+#jX��\��� �lv �z���@}������a�X{"Iu_� 1�<0�<�7j�=�5�tr�z���|�6Qh%7,s�Z���?��/�k���c�Y�3de������-�^K<��\��s�-�M1F;P�5�t��h���p0�_�V���������}	ݜ%�R����QG4�\ON�ͷ�<�A�}�lk5ā��{`ƶT1�	�$9|�&dV��(s���	�/#��g�s����I��I|���y��p��+T;�O6.v�g�IۑC_w�8_�p��sM�$��ݻ7���4!����Mv�\;�_"8������f7��d�)��+�����NIJ�孫�e�1�h��"i���T���F��diV2#8;�)WF��x^/����d���%*%�B��}u� �y����>�1����L�1�����%#��r	r2��������}6�_���g�CohyyY��|�.��w�b��Ws�u�kM�3�Ctʆ�EҊ&��'���L�1�i�,q���&��O�	�3����r�PK   +��Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   +��X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   +��X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   +��Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   +��XA�r&�  y'     jsons/user_defined.json��[n�8@�b蟙�/�ʟ[w���H<�EPP�
�%W�A��̚����	��N?R�uH�ޣKZ~�V�K�D�^u�JUՍ*�qt���n} >����ӯssj�|}�m�˅�v�a����zQ���~$�r4S����jݩѥj��ӈB��M��kDt�,׫�z<4<ݶ{���j��S�&y�$E�a%RXT�<F�gR�g�eOݚ�����j�����Bo��"�1�"�Uy�r���V�Ĥ<Z67���h��EqY�\r�b��E"�H��ʌ��PY?^��7�c��o��\�+d�]�˺9m�6:y���bZ�˹���{s�G����z:t�ޙC8~<�	�q_7�����洼\u�n\�Ӝ���i����=$�\��x�'����)����z7�s�+s��t��������J��=�t2�x V������j5�_����z���H�6��՝�؟zW��T_Ճ���],�F5���C���2����e�[��ܻ�)@��s��\J�b�RĹ�ZZ1�����L�dE���	bRP�'��"#1͒J(Rl�����q����دd���l�&�l�VM��4��W�3��XW��E�讐!E,��vG�ɴhoe>WV:=��e�6�5h?dS�}�r��;��c3+}��_�濷w��w:w�֩�!o���ʺ��͍��k<N�}^���5�;S�w�Sóv����ڍ����g:�Kv�±�o�>�g��1�����>�d�7��E��ѧj�VW���O|�Cl��	���� h���T(V�!Vjo�d9��r��eBl�q8�
�aҕ�iGg�F�O������ZݷU��u�ҹ�������J(IQ�����JJT��Ld,���H2�*�#��X�A,Q�tY����"e,�|;
Տ���NN�mw��ws�2r�]���ʇ)��3=��8�t���W<���O�0�.s����/��^Q�p��+�2�������6S��C��@��64uL�@Ы�s/T�P�Nb/3�����M�t����NX�O�I�m�,�'��}"�ԟp?����r����P�������~�-�~��BQh���¶R����������~��ce�췊�VQ� د���@��+b{5� 9<[�||�οf$�]C�@���rX�:c@4Ύ/��a����,�v�F��t���3��@2;��P|2�g<uC�\��/uԶ�f����¥@t<����QG����G��Q���8�Ɏ����ɶ���sI�5<LvL(��$a�cZ	u%��c�&2Y�ɎE[
$ga�cݖ �8�k7E�0ڱ�cPtXC�X�Q(:�!s,�Z�1[B�a�IhE�lq����/R�L��Z*<��՚;栆�Te�9��&���q�sPCMT��;���* T�,�;f�����h9&�ۅ�al \�	�=�f��@��K X��^��_S�X�����%�0�0�Y�1#��%�0�1��1��B�,#��y,������-��*$�cR����Vl�B��]�چTHU�;��^j���۹��k�B���[���k�B�B Z�],�V�@�l�6XHU�˶k��T�@�<z��B b�@U�2�T�!�@U�2�QT�!�@U�2�T!�X�
��<�|�7m>�z_,�{��O &�C��� !r�n7o���6�e8���jQ6�J�7e�~ӛ���C������9�0�1��%F��$⢤�$�������?�PK
   +��X�2�]  ��                  cirkitFile.jsonPK
   @��Xw�'<�  �  /             �  images/0df5ba52-08e8-487a-a0bb-947223afc81d.pngPK
   @��X`�/��1  �P  /             f7  images/4cf22100-3898-4fbb-b8e4-32284cc8d12d.pngPK
   +��Xd��  �   /             Hi  images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   +��X�IM��  � /             ^�  images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK
   +��X	��#u } /             �� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   +��Xp>r�  �  /             !� images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK
   +��XA�r&�  y'               Z jsons/user_defined.jsonPK      �  {   