PK   %��X�M��i  �;    cirkitFile.json��%9r%�*��bH��7��O-�0�J�ƴ�Y���Ou�de�DF����ڗ�gZ�o�̸׿�ݎe���$tU�u�?47�F�?�yj�u���=>�:<}z���ͷڿ}���}��o��7?�������/O͏�{��˟��?�8T�����cn��$��>u�7i�\�UC]5:�V{?��~P�ͷ����y�mA=h6��`��ԃec�ZP���kA=x6�����C������������M�F�U*�T9�SUwuW���U�z�9�`���Ɵ�r-�������?<UO����?>~h��?�!7���*��m"� Dl~�ֆ�3�����8��}��@�G ����?�Md�Q�m"���lEd� ���4l�L���Fb���6�����F!=����[&�=�7q�O ����X�gX�g��%��&�=�s=�?��Md������p$}1q�3�3��!�DF���&ԃ�k����?�Md���m"� �L����������&2
�.a��(�q�m"���N����;�&ԃ��N����;�&2
~�d��(���m"� ���c���N����;�&2
~�d��(���m"���N�	�����m"���N����;�&2
~�d��(���߮;���!w�<`���=?�ۥ�/�=�I7�JU��X9[U탯�7�ru�U��si�p�����}�g­�'���8�b>@��$A�< m�R��P`��g]�|��e¶c����Ʀ�+��j۶�b�Eקa;��da3���a�+��6ӫ��}�1 b�Z�L�"b�Z�L�"b�Z�L�"b�ZP[	ND\�)RD\�)RD\�yM� ���Pɏ�[�DT�h��HDE���[�DT����HDE���[�DT�����CE���[�CT�ȹ��CE���[I7��?vn��PQ 晀��jZ)IS����z*i��j��yy<i5Ë���`2q�	V��O�K����	�	��/�'�.R��?��Ml��PQ�ǰ���8�a[	;T�1l+a��°<{u������ei�Tk�1˲ƬXs��?f��1���w���Y�>�j�+r2���D}���!d�W�?��Ml�cQQ����\*�z/Xs�� N�\~;��
��ќ�>��YVl�[~ԇ �n��9Px\$��X#������t3*
�ʟ�3.B_:�*�c!��)�v��	����K��3<�"u{�?dn��QQ����:*
�HY ���+�<P�mgR�d�_=8F}@>  !�?�meRQ�]1 �u�x遺l;Ր
�5^z�u+ӑ���\��}�{�r��4��@�7[��T@��7��P#o�k!��xy��N�u�F���w���3l�\'ܓ�����mĞՏ�Y���>�6^@T��Ǜ�v���ZPt�N=X,w��ƢS˝�rE����$˝�rE����
�]�rE����C�r��A�i,:����%,wPt�Nݗ0�Cp7C����Ƙ�M賕s�Y:Xza�i0�r��t����4�m�\3p�e�N�0����1�+�8X|����9X|��|��:X|�����;X|�O�ԭ���<X|�:���1r����I�U��]���VNX|�O�'�,���߼;��7����x2`�ŧ��n�B�Co�ww�����)��?����c������œ�',>�WN	���',>Ƨn>3 �,����U`��������k/,>�W�w���',>�W����',>�W�ԃ�c��	�O��b `����O��2`����O���0���NoC緁�~,X�X�|���`|�`�?�|���`|�:H{�����*�?�����`|��?�����`|���?�����`|��	�?�X|�o^ti�X`��K� �A��,�R��X`�i0�R�����X8����-�~^����+E�������W+Bڃ��X|���?�����`|���?�����`|�5� �4���O��X`���c�/�:RLM�ĶJ��U��j�*�ޫ>�q�x�2�hjVsiB=X����J��z�`�s_��MX�`�هJ�� ���O������@�G�&@�&@' ���
pH{���	��d�?�h���`|��C����	�o��`f8N�������k�9���������r�z�O�񕲉`��z�O�񕂏=��4�1��5����T�tc[�J�z�<h�@�C$(�3`�
WeYY�A��H��mz�Z�+���H+�y��#�����jp:nѣPt���O�a��.VQ�N����^��9wPt��ԏ_`��.�P������^��9wPt�����X�K0���X���%,��CpEG/aI|X���qs���%,�K]89n��%u2�;�"���,߁"���E���@��� Wi<a�Xb`��"y��?����;PE�=`���w���	{��r��@�� ��%߁*�'�A��,��2��e|��򁊒T��*��@Eɓ���u-wE�@q�� ��`UD.NI]��",��%O؃�VEX|�K�����C}Z���'�A蟉]���'�@��ɰ��<a�X�a�(Ny��?�&��;P��=`M��w���	{�����@u�� ���߁�'�A��,��%O؃d���߁�'�A��,��%O؃��/X|�K���W��'��<aB?X���?R�,_���<a�X�`�-�d���gN���V?X|j[������# �O�ғ'�A�,�����<a�X<a�(�y�$u,����Jc�w�s�"W����^X|K�5Y�s�_R�K7,��_�}9Y;�>�U��X����M]Su)�*���.=���?B=X�a���y����VRWr�l�G;P�JX���m���j! *]`�H�&J}@�~�Z'�y���o��(��xo��b�T�����@1�� ��߁b�'�A�+>,��HO��^~�J�.���eJ}@�n��'�y����@A�� �i��}���\��=@��n�a�@MS��U��'�y����@Q�� ���M�����	{�������x��)�.�fݼf(+�r~��w�$*��ҍ\���`��w���	{ ����V~䒭�$�=aR.h�Z����J�x��������������A�o�m�;\|�W���B�?�}��*�1���dŭ����qƌU�*c�����*�]g�f���'Wc4׼����3����<�'^��6\�c��f:�fz�f��^�=R��u�I���'5_'��|�{�V�%�|3���XS�q�Q{u�G���R�C]��Ξsgù�z�!5_�5���܊���a��������l�)Z{櫲�h�aJ3�V3W�����L�3L�3�@��?��?��I��c�j��I�fk��z��z��z��z��z��z˝�0���z���Y���Σw���ϖ�ޞ��6r�e�;��f�%|�|���s�W�q�s���K��,�a�1_�F<ӗ=ӗ=ӗ�]�����Y3�6�"ݚ����Cަe�>po�X�g�s���y�;��\`�s���˜=h���̯Ԋdݞ;�3,�������o`�{������^Ԝ�o9�Gù5����Oޘfݞ9��	g�3_��|i"O/�3��K�{{��$ͼ=/b&ý}`ݞ��ڞ�ۯ����\o��'�0>ڽ6�!�q>ι��0Cܽ[�3iAx}l&.e3���q)�ski�,���Q(���{��kC�c�^��3����И��6&l�����2u;��o�A��r��U=h�������7�ݸ;����Ӧ�������X5]�V��ɗ��a��[ 4_��6Q����f09|ľ�Z�6Uj����!��b��|��e��k��θL�rU��X�w��A�i����wo��ꌰ�q����RH}�c����h�a���w���mԕ�%p�:���۴u���z_oݝ�|��N��6*�
]^~��+㚾�v���*䠰qwR����І<�JY*�\�_�`����m�5���Aiμ���
���z���Gcm�>�>sfl�:wW��6o�n�[�;����29Ӆ�Q��i��k���r�y�u �"���H�^����qR�uN��2;9YN�%q�Xʜ�e}=��
�Z��w8��s1�Vʖ�ٌe�P��]��d��&
��k�0�֬�H��ä[��^��ܚ��j���k#E�/L���E��x���>��y�)W�Zu���
yǘs��(���V��/	g�x�ω/	��k~N|I8�^�s�K¹��:�%��zm�F��Z)�єIl}�>�Щ�5[��|C}P����I��g����"R��y������|}s��|}o��|}�As��1�n#��֞�y���뾗Ê�/K�AW�!�>V�ml���Ö�&5�Xg�4�8�����z���䉴�c����l�G�ζqT[�t��ǫ(͙����uB
�m�1�*LSխ5Ul�:����u���|��I�ן��|c���3��C������R�L�[��u!�[&��K�����Nj���5�f��������V7���,r�!�ik���|��I�ן��|��cgR�t[���6\�pN}�:��Rfkq��|��ck�ɮڎC�����`UVZ�j���ꨶ�8R�e���ϫq�����Q2�j��u�vAjkY��|��CʓOe�ri�T���y������ڎ!5���������C�����ͷ<��&>��5����yCeh��dH���dH� �A2����dH5�A2��@� *��!?6�x�"
QBq2��2� ����"$,h�,�I@�0�⶞�N�_��11�"���n�%5�g&X�ְ������ L��#��a1\Â��R%]=21��8ʒ�N�c���⸁��R���	7��qca}���/�B�L蘘`qeIM5@}��}�gK�o=,��,��^,�[�|eIMu-@�`�q��(Kj������Q��T��	�-l>�����" L�����q�%5�.a��q��(K�wcQ�`q���8ʒ����0���q��8�`qeIM�l@�`q���8��T�	�	�,��,M_�Cm��⸇�q�%5a��q��(KS�&����MX��8~���m����(KS�)��Yɚ>���4YGeꞹ_��K����LL�8�bI+",�,�f�w���%���d��WD-�B�?dRKՠ��ԏ-���ԏ���������DD C��"""�!J^�)��"qQ�aq��D��܄l *&X�&dQ1��7!��	�	�@TL�N��b��pB^,�����`q��D�X��8!���	7��M��3M��`q�bis���	�/�Ʊ	��b���R���,�_,���d��`q�j�E��qXGY"�Q1��8!�*�aq��D���l z��)>�zuM��	����iJ���K�Wj\�˦b���Əcό��l *���	�@TL�'��`qe��WD���l �"&,�_����I�+�b20L�u�K6?�����0o0)���	�Q�HyETL�u�K6��a�*�l���mm��`q��D���~��u��	�@TL�8N��b�׼"H����5�(�,ZS2���pۛ�8N�+�b���=hM�+��n�4�]`b���K6�'X'�Q7�ʟyETL�8^VC��<L+#��oc��7��gY-%�!X�V��u�vg@ϰ"zK`�"X�VF�W#�X�V�`Ex�"�J`�"X���Չ�*�U�`�� ^��X��<G�5��*�U�`UQ��(«V-�U=$^��X�V�P��Z��:Ǌ�XKN��0�Q\"h�ڒ�,í���2h�ڒ�-��\�@���Z@!AF|i�%�Vˠ-9�2��(0�Zm����VF����2h�ne��Z-���Ő�VF����Kh!��2�L�(2�Zm9#í�*A�eЖ3>22�L�^B��	FF�]&�Vˠ-g�d�����eFF�]&�V/���]fdt�Z-�����VF����2h˙Dnet�Z��dt���e"h��rFT�[]&�Vˠ-g]e���e"h��rfW&1IF����2h��cnet�Z-������VF����2h�Ypn����e�ˬ�.�2�L��A[���p+��D�j��ƀ�2�L��A[j%�p+��D�j����2�L��A[jW�p+��D�j����NF����2hK-net�Z-���D��VF����2hKmnet�Z-��Ԩ��V�$��Q2]�dt���e"h��R3H�[]&�Vˠ-��d���e"h��R�I�[]&�Vˠ-��d���e"h��RSK�[/��D�j��6��2�l-�X��R�L�[]&�V/�E��x]�et�Z-��Ԝ��VF�-����BE>��|����e^F�y]&�Vˠ-�e���e"h��R�Q�[]&�V/���dt���e"h�Z�AF�]&�Vˠ-�>e���e"h��R�T`�xkX�C�>���M�c�p�*����>F�q�@^�`ǭy��z��*��^"�\��~5L�W	��k��
�U��ګ�o^��zp���U^%���z�*�W	��k�R�Ë�zp��Z�^�W	��k��
�U��ګD.n�
�U��ګD.l�
�U��ګ����:Z͔:��@{��*�!�%���d���:Z��Y$�2�K��ګ'�"���_"h��^=aɭ�A{���	�Hned���WO�Er+#�D���z�,�[9&�v��*��x�U*	2�L��ګ'��v@��^=a�� �ˎ�^����2��k��0��VF���=^{��Y`LA{��*����A�eGk�RI��e"h��^=aɭ�.A{���	�Hnet���WO�Er+��D���z�,�[]&��x��f����2��k��0��VF���=^{��Ydf��.A{���	�Hnet���WO�Er+��D���z�,P�=^{�J��.;Z͔J��.A{���	�Hnet���ګ�����L�$��2��k��0���2��h�U*	2��h5S*	2�L��ګ'�"���e"h��^=ay�AF���]���ˎV3�� ��D�.�^�p+�ˎ�^=aɭ�~��j�Tdt���WO���D���J%AF�-T3�p+�ˎ�^�� �_v��)�]&�v��*$�����z�,�[]v��)�]&��x��f����2��k��0�D���J%Af��h5S*	2�L��ګ'�"��P���W!$��-T3��]v��*�]v��)�]&��x��f��
����eG���0��Vbw�x�U*	2�e�L!�VF���J%AF���J%AF���=^{��Y���貣�b�$�fz�,���L�E��k��0��VF���]���6��Vf����{���Ǐ���Χq�)V�I�j�T�tc[�J�z�<��8xЊ^~5Z1,���lk�1c�*7DS���U������_�e[�+b�B�`��+b%B�$���u ��x�Ƹ�����8����6�j]W��S�NU��]���Vu�u��~�!Y��'���n"Y��%���N�V�>��R�aXٍ2$+�Q�de�2�X�80��F�ׁ���Q�f��Q�fe4ƅ5Ƈ��PI3��b��b��/6/6�׺W]�1���ڻu@3��b��b��b��b��b��b�J`��N^�Ǧw�A�^f�R�e�����Z�9f0^l'/n��֖3��x��x��x�͈13
��Q����C3������=Ƌ=Ƌ=Ƌ���m������j��/�.p̼��Ƒc������������a��Τ��txx��e-�cf���$:�������xq�xq�xq�xq��8f��j�s�&u�x'/�08̌"bf�̆����x��2RqV�ԥ�[͚짗X�#s�L^�1�L^��y+���؄��Ӯ6�fLق��r�PW�8����P��n�ϒ������7���M[��)��ob[�a�*gu]��u��m�U��n��dE�-$����u$���]f��'�t,B�c�^WnPcv;�UqhL���!&�K��;�2u;��o�A��ʃX��A�J����z3�},$+���6}�\��d�M�j����O|��Ҿ��.m���f0�=�}_��m���Cߍyz�:BQ��b��ܿC�w�ev��Rg�j��S]��N�XHVv�4~Lu�]�8��dV)���1�F�q�ð��deK�tl���-���Cն��^��}[�_�P��bq���Q�ju�&��5}��}�U�c��.��0����u�r���m�
*�޶�Y��7�
ˮ�#Y�]M�1;|�mէ��ΌmU���tۦ�mݍ�_HVvy�]�v}��޵1Go��<uMեЫ����wzkI�dE�I����C�b���ʮ<!Yٝב�����7g YI{���]}M���fF_���5+�43�)oH͐8f&���8��C339p}t,n.��qM��<j�<��z������WΛN�:֪���D��gX��)$���JU�b~�,;Jo�2+*���Σm��e��IV�^g�����&Y�{]M���zڍ�F����zM!������N��!̅HV��B+�c>���O��;����'$+��	���Z���R���xB�:��b�w?��f��9e43��#��/kJAW�!Ǫ>V�ml���AY���\P��'gə�𐕨��VǪ�}_�.�j�m�>%�����LS�`�h��X�!�P٦+W���۬�c���]�X�I��]^HVvy!Y�אM����P�R]�~0Uꓩ|�㐺.����!)V�ׅ(Vvy!Y�奷�غw�Sy��z�Z�تU=t��DX1&Y��de���]^bgR�t[��˦\�ڦ�J�I�V)CX�#Y��%������8��{�}��e�+��������N��쯯v�P�q�ʓ��6���M5z�:m��EX_�X��2�<�Vf�Rۤ�Dm���k�`��{���$+���i2������y�|��/fۧ�����h�JC��ʛ4���;�!{:�V{?d|�p�q�������QCe��;Ȑ��y"�!5�"�!5i!"�!5�*"�!5i4"�!5�="�!5iG"�!5�P"�!uѴ���ڸ����Q��E�c0�b��o�%uYT�`��o�(K�r��	�5,��,���>&X7�8���.�1�p�o��,��,���J&X7�8���.�>1�`q���8ʒ��H�`��q��(K�rV#�aq���8ʒ����`­���R`q���8ʒ�V�`��q��(K�r��	�-,��,��o&Xw�8���.G�1�`q���8ʒ���`­���aq���8ʒ����`��q��(K�R� �	�,��,�K���,�{XGYR�JL�8�aqeI]jL`0�v7qۛ�8�aqeI]Ji`0�⸇�q�%u)�����Q�ԥ�,�X'X"VS�'�X�d��WDD2D�+""�����I��;
���I��!
��pI��
��`I�� 
��PID2D�+""�����!�qa�	�@TL��M��b��nB6,z����`�D����l *&X'dQ1��8!��	�	�@ԉ%,�����p�o��	�@TL�8N��b��qB6,�����`q��D���l *&X'dQ1��8!�*�aq��D���l *&�J
n)�	�@TL�8N��b��qB6,�����`q��D���l *&X'dQ1aq��D���l *&X'dQ1���q��8N��b��qB6,�����`q��D���l *&X'dQ�~`q��D���l *&X'dQ1��8!��	����ބ�qB6,�����`q��D���l *&X'dQ7�aq��D���l����?<UO���zE?>~h��?�!7�$`���/�Z����]	^��X�V�`Dx5"�J`�"XՃ�Պ�*�U�`ͺK�W'«V-�5σDx�"�J`�"X�E�� «V-�U=D^��X�V��DxM"�J`�"X�C-�k-«V-�����%�Vˠ-��2�
�.!�%������2�K��A[r�e��Q_"h�ڒ3/í�A�eЖ�neT�Z-���a��VF����2h�YneԘZ-���)��VF����2h��neT�Z-�����X��e"h��rVI�[]&�Vˠ-g�d�����eFF�]&�Vˠ-g�d���e"h��r�O�[]&�Vˠ-ge���e"h��r�R�[]&�Vˠ-gDe���e"h��r�U�[]&�Vˠ-gve�dt�Z-���=��VF����2h�jnet�Z-�����V([Q(]QF�Y]fet�Z-���͗�VF����2hK�net�Z-���J��VF����2hK�net�Z-��Ԯ��VF����2hKn��.A�eЖZ"2���2�Zm��"í�.A�eЖ�.2���2�Zm�Q#í�I2��d2����2'��D�j��f��2�L��A[j�p+��D�j�����2�L��A[jQ�p+��D�j�����^F����2hKm0net�Z-���8��VF����2hK�6net�Z-��Ԝ��VF����2hK�<n��|����e^F�y]&�Vˠ-�e���e"h��R�Q�[]&�Vˠ-�%e���e"h��R#S�� ��D�j��֧�2�L��A[j��p+��D���h��t>��U�õW�[�z�;nȫ�õW����U��:\{��U �<�[�*��p�U�7/Dx=��A����X�^=nȫ�õW���Ex=��A�@/«�õW�[�*��p�U"7�[�*��p�U"6�[�*��p�U�^Fp�fJ���H.��k��0��VHv�讣�LO�Er+#�D���z�,�[�%��x��f���H0��k��0��VF���=^{��Y$�2RL��ګ'�"���c"h��^=aɭ�$A{���	�Hned���WO�E�,��2��k��0��VF���=^{��Y$�B[b2��h5�f����2��k��0��VF���=^{��Y$�2�L��ګ'�"���e"h��^=aɭ�.A{���	�Hnet���WO�Er+��D���z�,23IF���=^{��Y$�2�L��ګ'�"���e"h��^=aɭP���.;Z��Y$�2�L��ګ'�"���e"h��^=aɭ�.A{���	�Hnet���WO�Er+��D���z�,�[]&��x��f�'dt���WO�Er+��D���z�,�[]&��x��f����2��k��0��V�(��.;Z��Y$�2�L��ګ'�"���e"h��^=aɭ�.A{���	�Hnet���WO�Er+��D���z�,�d��.A{���	�Hnet���WO�Er+��D���z�,�[]&��x��f����2��k��0��V�̇�.;Z��Y$�2�L��ګ'�"���e"h��^=aɭ�.A{���	�Hnet���WO�EVV��e"h��^=aɭ�.A{���	�Hnet	m��Ï�����O�S�\���Ʃ��ƶ�6��:4�yP+b�@�X��gE��8c�*x5Tn��j{k�8v���!��g�de�]��]vIVv�%Y���!V�J�XI+5��@΋�^�q_��_�q`���mj�0��Rѧ�)�������]����Ι�(C���O$+��D���K$+��D����(C��eHVv���n��y�y1޻ehf0��ehf0�1.�1>�1N�1^l0^l@1��������������������4��x��x��x��x��x��x��x��x��x��x�͈1^�0^�0^�0^�0^�0^�1^�1^�1^�1^�A����������������������>���������������������Zf�xq�xq�xq�xq�xq�xq�xq�xq����&ߌ)[0�Tn�G]���]�bj®!��n?���vS����Vi��Y]Wmc]eb�{Շl��"���'"Y�<Ѯߑ�캝v���U�{]�A���TWš1]mL�g�de�]S�co��t�*��XՃ6���E��f��XHV1F�>t�j�o��X5]�V��ɗ��a ���b�&����j�ߣ��U�ڦJm?��8ġu�>�X�ŒԹ�����*W�Ό�P{���t������bi�����q�=�ɬRH}�c����h�a��>����F][b����m�����6F�����be��}��JU�Kd0)����+o��;�B��XHV�#fh�Ч�Rօ�%W�1�*��{�:gMO��+,�ћbe7z��>ֶ�S�dgƶ�s�V�mS��FM�/$+���΄��uջ6��ms�����z�z�tGx�IV0Xv��de��HVvGX���y�ʮ8!Y��&$+�҄deW�м���������~ �̮�<j�<��z������WΛN�:֪#��$+�#��:�#)eKo�2+*���Σm���K����?*Q��k
��]�q���Ѫ<�*�^SF�>�*�}��Sck=M��?�X�e�de�]���o#���xB��;����'$+��	��@΋����f���	�̮爤|�˚RЕsCȱ��Uk�nl�@P$+�++�	�Yrf-<d%j�<�ձjz�W�ˣZg۬O	�$+�9�+�'�?O�>�*۴c�j�Tu��ql�:���KX�$Y�?gB��΄be_C6]r&�C�Ku���T�O��C꺐�/���X�_�X��de���c��UN剢�juc�zT��5CaŘde���]^HVvy��I��m��.�r��j��*u:$�[�A瓬��[[�M��v��=�>G̲�T��MWGEx�IV��W�~��S�c�o��}��T�w�ӶjP��U���=�����Uj�T���V:]uM��xoa=�d�5�?����o90=~x|zx��ۛo�}���O?~h�<~������Oo���o��8�+��N(6I��O]�MrD�3�1�U��j����)�{��A)g09P���&��A��r��}�W�ڧ����橧��s�B�s_��'2�D(��z��'ƹ�8&;
疝��6�o�8��k1���q_����+��V�n�j�Y����4���Z�c�ju�7Bc����~ fl�wǺ�a�y����.�t��;s/xNOԉ�$<([��pv���0��@L�a��q�{��}{ǹ�gߞC~`�����w���[�x�!Zng�D�|5�MK�'P@BT93̂�����t&;�.5M�F������zkX=�ԭ��c�pW�l�b�*�7��t�qdz��~N��/�3�L�mE����g[2���r�D��slx�h5��y��*h9=��/έW&�Ԕ1έW45͌sk˹��1O��ζrkb�,c�c�����oW݌���x�U7#��2�z��&�˲"����8P���ԉ�Y����L�
gMTQ�`ٱL���N/��
���R��W\�&����F����OZrᬭ&��H�e�&���<��=����y�ۯl�P&so�YtH�*���W��p8�k��9�����H.5�S���pV$N~ ����߿bq������(N~ �1�clv8/������s4�g�7<'�G�6uo~IT�u���y^Tk�L�����_�c�s��OXX�:����������q���͏#?s�5(^������XO_���k�������C�_J��m������a!B����3���Љ�WD����Y���~i��_�����CP�S�1\�3��w�����^��s`PpOul�~���`���`�<y"0�?���2_�
 �8
 �T�&���p
��
��
���/b�����=��A�=��A�=�A�>�@!p��C��=��b����W����+�ɣ_D`�
��9APq�;5eO=��?��f�#��lF�|͇��(�J��u�����d�.�Y�Ev��7 @�oh��#p�uB�rb������_�L �h�����8!�G�=(�G�=/�G�=6�G�==���"�#��%�#�)�#��,�#@0�#B�3�����\���:ΉA�>�	A?܉A�>�	@�9��s�X?�)pB�
}P&��U1(��V1(��W1(��X1!}���{���{��玮�����BP���bP���BFD���T��ÿ��&��4
�Qc
��	�/��1-Q��:}»�S��Ї��~��6wz�Z���`��{��?שvLTDn�Հ3�6�qO���o�Ǎ[����>�G� ��횈��0����7���o�z�����s�<������b��������o�x>�����^F��僁Llj�@%ۄ�>p�D�6��t3Q�M���Llj�@8ۄ�>0�n�1�*�A%>5lj��9E=g70c ��m���׹8 �u���ő	n5 ��m���8 !Wb.�F���|�	���:&,@�Հ�;ٸ{4VvjI��bۘN��m-�|@ �'w��Jl��1�ab���G[Su�z X��<ٸ}4���M���|�	�Y�q��aGY}�q�k�Iw��| R�md��&�md��̷�J>
b��|�6TI��� D[��m��] �D��)߆*�|�x� �oc��� �S��|S8ba����O�6T)�����O�6�>@<u�xʷ1�5��  ���)߆*٧|�x��oc�E��/(�Ҹ*��|X������4s���-�Ɣt��1_�U��)=�k���X�y������W�sI' Bs���*�d D�M�JL\�)&��*|l�)&�#e|[������ID�6��bB=P�G�5JR�@�QlhDl�9%Dl�9%Dl;I$԰�����	���T����A����T�(���A����T�H���A����i"T�h���A����I�	 �n&�Pq 棈	�<�ϭ�Or� �y2�c�L��踇�ג��� �w�qk-��
�rK<���N^�������oc'/���7s:�"�7s:�8 �z3��^�d�k����0 X�H�=̵��A�O3���$G���v���&�� �<R;�o"��Gj��D@�����8�� D��l�B R��z`y�N
����U�b'�
kaz�
#;�)TXAwm��
����iB�X���4�� �o�yX,����B��2�Ŋ�;�,TX�Hͷ��rGK{Pa��|;�-T�hX��%���$���f���s �̥��Bl�"�f�������_�,���C/�1�Ŝ$m��Pa�sXk�Go��Pw�3�<ϔ��y0TX�8�182��<�Ǵfg�X��} �	w�U�{�����g�f����Q"ߣgv�ށ���&���c��7`:�Y��4�z�`�,�?,>Ɨ�?��O����?��O���)�� ��O���/�����`|�!��K`���4����5����;m��!���!t�8 �
F��KJ-�C�_�j4��Ͽc8�M��^ĵ
�T�Be�� Z�h�V#�h�%+�!Z��j4Q���Y�5aɆGs��-`���d�9Dk0B���n\��!����h9F��ˁ
4�hIF���a��6Zŀ��w��ڗ"��E�A�0B�Fx�	i����vZ���j�!Z��޽ڞ� Z���#�h���C��#�h��X�C��#��^mV.F9���q�5a9���-j�5a9{��-j�5a97�N5A�0B�FX�|�9D�0B�FXΫ�9D�0B�FXע9�����{1-[,Z��j4�rl�!Z��j4�r��!Z��j4�r �!Z��j4�rz�!Z��j4�r��!Z��j4�R5 ̡C�0B�FX*�9D�0B�FX�3�9D�0B�FXjI�9D�0B�FX
_�9��q�rA���)�S�5a�0���S�5a�����S�5a)���S�5a�;���S�5a���Уu
�F#,~��u����f%�h4�R�M)Z����w}�LK�h��*�P���Ph�*f��֋�p)h��~x~z-j<Z�x��#�h��r�C��#�h����C��#���-w�Fk��8`�z���Jb-yZ�j4�R�!Z�j4�R�og�Ƭv�bu���:l��񯥅S?�Iu�������U�mzW*7����X`v�o�s[P|JR?T揼�A��?,�%	�ۃ���w�$!��;�?��`<�?,�%	�ۃ���w�$!��1�?�z�d2�?,�%	�ۃ���w�$!�y���A���;P�����U��� �a��AH���	��uƋEx�!���"�B�2�C�%�N�p��"`�G��0��-G��<a�!Z��):x� �C�,#<Rt��A�hiFx���	����p�����-su�^ҏ� Z��):x���������� ��:�U�!u��b��<a�!Zŀ):x��ҫ���>���WТf^�����1^��8`�Gj�0���q��� <a�!Z��Ax� �C��#<Rt��A�h�Fx���	�Ѣ��H��1�Uᑢ�'b�I�*��H��1�Uᑢ�'b8D�0�#EO\R������ <aC)Z��+�Q-[��� <a�!Z��.� �[�X;�x�>�R��#<R�����u��O�R@�z�B*hQC��G}d��#<R���A�hQFx�B�	��o��#\�Px�sġ��2��8`�K�ֱ�#���%�R��;J�ꝰ��-y���3<apq^�J�8R���A�h4�x'�Y'�;<aC)z�^J���hF�T��n�g�Y�+R@+ 0�#�O�p�V@`�Gj�0�������><api�	�|?0�#���wy����V@`�Gj�0��pG���
�H���t��:R
�A�hD�,H}d��#<R���A��2h�C�,x� �Ým)�,�|��	��ђ�E|�2"���WF�>2Z�)�x��[2s����*#2�<aSfe�
�O8�J�
�^w���hF�Th�!z�ga��Ï�����O�S�\���Ʃ��ƶ�6��:4�yP�����AsznN3̙�9�0g��,Ü[�^��8c�*x5Tn��j{k�8v���!����������2�s������>2�'f���?l�z�溠����:����6�j]W��S�NU��]���Vu�u��V ���R��. ���R{7�ze� ��ss+C��F� �߈��i�8+C��FȠ9�[��2h��2h�!Cs�Rs�Ro�]4\O4\O4����D��D�;#��B�{\?5\?5\?5\?�\?�\?����v�&q���T��q���9 ΋c�nk��%��z��z��z�cOT����.�ݬ���W��S���똞똞�~�,�V��h����r���G���:?������b��b������������0�b���aa��y+��ܖ��a�Ś�Ł�Ł�Ł�ő��q�}�8>�����q��㓑;���Ed�oq�6r�6Χ��3�M�-1��i���q�͝�s��ܩ=g�4����i���|3���XS�q��fu��w]�u�����*�ܼ;�֫I�潹�^�bj�&�UƮrV�U�XW���^�!ߠ��M �_x��'�[x��w�dnߣ?hna�l���ε!��
u�+7�1{��84�k���	[ܓ�o��Lݎ���jЭ�\�cU�T:�>}P֛�nݟ�~s�M:W5�7ٕS���i����˦�0��d�o�_��GL~�b�W�j�*���w���m�Oi�q�ܴν6T}g\�O�*uf���;��ݠ�uR���7~LuY�8���tU)���1�F�q�ðuR����N�6����l=Tm;��?mݷ1��כ���߸��}��JU���lR~\�Wގ�w:�aܺ?����Sh�Ч�Rօ�%W��'�*��{�:gM�{)��ߐp��d>fw������Ι����k�n����Qo�����_;�>�U�ژ��=����R�U��]Z���=H��C�x ���k�<$s�F+���%Bj�1I#���!���x�2�"��o���9#�܆����ƫE3��̜��ze�D�7wg�2���[X]�x���W��ʼ8�N��&�c�u��r�t�ձV]��v��$s���ؒFչ�����f,S�����<'k�銳��-�ފ���-�ޚ��[�5�B1��x+��FS�UyV�Ħ��}�U��`C���lΩH��T��s
R��9��ƸDj�1.��o�K���c���c��#�������/��n%|�lxa�׾,]97�T�X���a����ʂ�~ke��~+M7KȬg��,M�G�:+���������6��͕	R��<cJ{.��b݇�Be�v�\m��n�ƍmSG?t]c73�I�7���~��I�a�%g��.Օ�S�>�ʷ>��B~/6�!���������o<o��u�*��$��X���U=�z�!�isU��~��I�7���~��cgR�t[���F\�ڦ�J�I���zm=?�������c����<+���1��u��Qm���[+�]?�9�W���3x�Cg4��]�����$������g��Uj�T�}������\�&����Oo�|i��x~|�?����o(��|��7E��e��͋�po���r�b���7e�_��e�]{�
ͤ}�M�i+e����8�oG�uB�.�O�|�C�����)�aʎ0��)-LiaJSZ��bJ�4��--�� N_k���$�&�3	�IfL^�2մ�4-	M!�������k[S��ʵ+-�R�S��i�n���6��ʩ.���:m�Ni�RS���T�T�l*e2����O	�S]�)�g����ciK�XZ��"�q�����E,-Ri�J�TZ��"�i�L��mg�F�͡Uo�l�|i�}�������͒��ݍ��툛�����������%�y'��'�E�܉�B�O��[&���L0���ȍ��J��/v5er��#�Y�bC�tj�!et�딉�m� �4nP�����O�Y���L
����)M�����I̫��MR)���&�w��3�1d/�q�:��L����9:�A�V���R*`��pЭ�%������tke�N�[��ݠ;~��*5��OCӷ��SO7��0� <at�
�����0p��w�(qq�7�_@T��$��5�va��� G�};O�[ �ψ�s��,t�^_�$CF�������s��H�=3�ߗe��t�2Kn9h8/�Yz���pR�CX@Tsq���B��E�<�2G���x'S�"�BT��̋�_a�#�\�,���=���P�}3��q��rȌ���!��H�*�R��E�7�W���J�=y#�z�v)��,����@.�G,��v��*&X�**Y`��j�V0������58�L?�hӞ4^��y�	�¼jm���P��0ѳk�����J~��YX��FV��ͪ��%D�o�hV-����;G�*�h阬��9����xB��d����b��y4q���Z�!��`p���nm��x����B�qkK]������|stk��xX���nU('F���5�7�v�B����aM���P"ݚ�����s��R��Is&°��T"{�ʴ����[]?#��������4r�b"�;��W�ר�/������W�ר�V��PKB����Q��r,L7<{X`���#��9ؽ�2�8�t�g�}V���������_2�#���I����j�0�b~كd"��/�Ox����/j��ƀ��`��8\[(�-�֜�P���"^4Qn-���~���q��AI�K�9����,曱�4x�l��ម	\��*���XyI�3�l�]�\]8#��3V��{~�дÇ�����y���:<S��/��'=�ɼ�d�?ٗ���'���_~����Oa�Sz�)��_~�g?���50}}0=2}}2=4}}4=�������v}8=:}�D�I��'��G��G��g7��6��6W^̜��缘+/f΋��b漘+/f΋��b漘+/f΋��b漘+/f΋��b��+/v΋��bބ��-t��vz�v�_�9��J���i������+�vN���i�t�+�vN���i�t�����+�nN�����t�+/n΋�Y漸+/n΋���漸+/n΋���漸+/n΋�����+/~΋�����+/~΋�������9��_y�s^��?��_y�s^��?�%\y	s^�0�%\y	s^��qc���a���g���|�9���g�����9/��K��������y���ë������Ç����T��y�y�����c���?���)�k�����3(Ҕ��T�k��O?N����<���7�s9���~�������~(g�sgd������|Ae�z�c�ɿ�y�z��s!]z�d�e&�w}�Q��ԭmh����c~��o��}7M>�����t'������������d��7�Oﳕ��͕���S�axy��V&�w�5����˿x���[_��MZ�,h3�̹�ο�ɼ��?�����S���3o�;���a�S�������s�������EB~l~(.��}�͇�ʟ����o���>���_�~��������o��ç!��ix����޷���4�ϟ�?��|��w�#��|�il�矞���ۿ������?���C�����}�	 ��=���^�c�f�_��1��}4�q]S�Wp�>���k��X��+�}R��$����O~����-����*:��_�j��F��Qkm�Z��z���8�W�����i��̟����i��̟���Ӽ�0�����W�f���s��������#��t�]�oS�{kW���P�a�U퍮��i�n赮S�Z�kH*q��p�x��d)��o�D�Ͽ�ۀ^�Ͽ�������F�:}nu�vy&t��ι�,��r�Bd�s����R�����>۪_=�Vw������m��/~���(��>��/��/�����>殫^�^���^w�I�#��te�D�?�z���_~��|�a�\��x�!������ü�^~�w��sO��Py�K]�~�w+�/x��4{3._�ٻ��ѳ��{��z���5c!����I��P��'��^�3ǅ�����~X'���a�z�r�]�ެ\���O���)�\V�w+�ە����j������q�z�r�[���_�,�������~�z�r�Y�^-_��_�+ׇ�����v�z�r�Z�����W��+׻���eZ�ؗY�����������i��ݛo�{�����{���7���o� �m]7U=&�'}V���U�}V��Q1�����~��V����wi۶u�e�T��}���C�T�I�]ۗ����څ��󅽯�=[��۶R�vCg����s�����Oϯ�1�4_����;6�J6�jU�
�]n����}�oC1���﮳�/O�׿{��e�w�B�q��K�v��'�*��牥m�jo��������>��Ҹ���+�J&�Vy&�*�m��m�+�����Mj���v�bJ�r]���J�:���V������c�J�2Q��\&��*�6�?ۏd�����קo���Z���^���/�~|z���>}z��Oo�[g�����a����F�=ll��O�V�ؗ�8�g���,f��7���ެy�UHm)mS�jHY�T��yJ��D����,zXRٷ���y�d��T��Mq0v̓��ac?6C=�j�IU.��j�.+����g�)�m�.��Ϳ>���4<�����|������7��?}�o��z���M����O��o��y���7�Y|������˿&C���м��`�i�qh����^� �ʹ`1�̄�Oo��7����e���wJ�n&S���%䝂zu�j��9i���:x��⍴�1e����Ͻ��v��b���̵KY���,EZ�Or��Kk� t�?�_f��]~��fZ����xߌO?����>�?�6��z�����sٔy��7�9�6v�J����mM5x+�e-�7}m��z�g�j��s�C�������/��Y_^$�������)��{����u~�i�����_==6}~������PG��j���&ެ%�G��<�尕��`�J�35$�w�hZ#Uz$1g�����em	N��ǯ�N�����ڙ;\Ǆ�n�5�1և<5�s�8湧n���j]��7�@rR=O�[�qu뾾[x�KX<�s�䶢����ꬬ:�Y�t�h�\��8���"��Rܡ,�]ݡ��}]w��_E_����W�K��:��)>/ތ!Y�&KӺ<u�ݘJ��4*�������Ji^��x�K\��oç����������o^]��g�R������:eR�w�O-������/�@�z[g�u]��Bյ.I����ax�G������ϗ��8�����o��R����WꝾ�k���ߦ����?�$������vx���o~����M|�׾Byҽ�o��wm
����v�,ˢ�y\k��V���͗��X�Ȧ�Ӷ�HE�i3�������kv����_<���s����璪�=�����_<���s/�M�s)e�i����cj�<W��q�|7�NH�k :n�2Y��7�q�h�_��o���{�*�����o~"�������h�BA�w��~�stu�]CK~�!k���%8��,VeY쇱�k��!}����e\�vl�ڸ�R�.S��̣��_��\�|F�޳_ѷ� ��5v��*��Ʀ�-��Zk��i僽}ݻ�����mե�UI���4I��B�N��B�T�u�/ivӋ�m�T���/��]����8���m������#��M�%9.���Sr��d��ܧ����3mB��vN�k�o�(�r]���KG�t�7�v͐�.�j�l��e� G��j�o}�lP�~NZ�کw9l�d/\��˲�џc,_fC��ė;��ˌ.7���g�L��7�.S�5]�ۛ�\&>�G�K��:{�*�~y�#�����/n�^������_�������Ӑ��.�a��Ϊ�H��"�ƪ$��׻�>?D��Z~1��d��������j[�ϯ��{����^9��wyV��KH�o���1�y���&��!t�̌R��X��A��&����j��e��3yNu�]�_R�>�wep�S
���a��[���������z��%r���2�K
��߻���6Q/����!n?O����ti'����I������^�Y�fƷoO�;��cf]��a���W����]e󜨪Ƕ��7U�!����DzmH_ޣ)��dX��#�SZs�����t��C��.����W�����+�D�y�+3�:+:S~����'}���Mw�>���LS^Ł��k}�ַv�ܚ�$k����_�a��pXҧ@O;�v4[�l���Y�]����E�WpX�'h�G�@��K�-X�4k����\u�d��rD3\�qݼcbhs �b5�W��|v�-�F�&K���j4�C���V�^��,4�0[�v�U�D���y�;\�/Ǎ��'�Ep�W�����N^��H�`���s��4���G؅���iu�W_q/L�^~2������6^}) q_Aƫu�u��A����}�f�^�޵N�.�AQ�����ꗟ���/^�g��JI%�փ2C��&���fO�t�5}0C�Q�Y[�|��p�=�r�U�e{Z羪H��;g���_s��6:�m���d����VQ���Ƶѐ8�|m����y����eT�_�j�l/?�r�VN���Y�a���{���ջ,���.�J���x�}S��J�E���}���r]�]�J/���ar��yX��O����n�����wC�����4<?�������]�^�?��������!�e��Wn:�{�����?��_�ZM)T��.��?���|4�~�j�����7H���������Ͽn�7��w�}��T�������LKH���~���S��/�־.�W�x{�̞�̫��tm�/��O߽�Sv�[��ۿ�~��s����%��
��>+N���ݻ��e��Gt-}�}��2ݧT��~��˂!E��e_+�X1��G+�>���!��2E�>��NG�ߕNP��P�����S[�?p#�v�%�G�B�+�JE�.�.�E�8X �"���%�
� ak{�#@6�ux�{~��w<F�;~{Yp��F0�/���,��2�hg��G���΢����9K�w~��o��Q�吶!�v\�O��#`�C�ޣ�sS�x�+�.\�Y��g.#�L�򣭡�C�3���_>P�B,��+7oy���ܝw��E�{⢒cHq�:7��1<�1�1<�1�� ���Eaq�q�mF����X۸=79����=H��E���:���wWiE
*�ˈ�qh&B)^�9���Ϯ����� VYo��>D���~��J�,���XgN\%�K�7�R��'�b`E����>vS�w�y�.ae���hWQa�������5fWS�R�朊�-������8e1���IW�]t�����9��α��|�a爴�q{YH�S㻅Y�UT�P*���ș�s�������`wy{�]���^�Z�)�w&<�n�dB�vڂ	�Y��Y��npjH�w��+np{U��W靫֢A�0)���E�.n��npj�x���wW�H����ݠ3��G�h�r�Y+�:����r�@�wW�D����Zz�z0�=�JzG��O7[tи�q�2���� �3��k9�p��Gㄥ8��K#������qu�J�ow�%�G ��S��2 �2i�׊ V ,�?:��b�ǧ�5��믔�W��+,B?���(j�1�7�Q�	�b�k��?�����Ea��Ds�t���a�����@+��a�mJ��z���]�s˫~�N��
iq�R�WQ��	�ɫ�ȶc���WcS����U�m�J���\��E�<���˂�g�@����O+�Y��ˌ[�,�W�±���aסq9r�.�n%ɪk�^f�ӕ�9qup���B6.jJ|lM�8-毊$��v�"P��4I�bk���˸��a,�;i5��@TI�L݃%����_f��"��ɣ�o����é玲Yr̕x��Oػ�n>F�p��V{���N�9�.[�*�`�l�]�]N�T -�T��T�W}���r��ek�%��Rs��6��|1E��σ>p�� 6�o�wt=�6��-Z\P�����9_.{�V�[�l%g/�fH�~�%aЈ=pH� 6X��:����f��]���׏/������d��yi��f]����Sy������~����ߛ�#g�S���c;J�]:6X��ZX�-\���w��~���e�?��t�Z��q���H��r.i�Iܧc����,�ۺ���~w�Z�_�wg���8��|ڇ���?����H�����y�ZN����^^8�K��_���m߅q;���;���x`Vw ���Y��gE�{����5�;W�8G�6$ �p�S��`!�����Ӳ�~{Y��Oq��V�;�jd��&~�w��?��	�������ek�~��K��$1K̩$.�;w�@����s�.B4/^q��/��f���夜�M��U���!V\���=yR� V��,�=�<�w_T���z�� ��z���ݖ��*DJ1��S��=b�)}d�R���S}WymY��oqϮB$�R�$ftS9<A`�O���W}�`���>�Aƍw�%�<H���E��U_1X�>*��+E�|#�,�g:@\NX�� �V6�8�ۛL'`��QseV&��~���ڞf���"�;|9��Z���8|D�rf	�@�}6����%�G����'��
�8��?�u �U�����3`e��~Kd�c�-캖�Ԅ���JXS&�9=D�	��J�v��Ĳ#ܗ ]�V�h�L��:xt=^��
�������	�9�<g������j�L�ݹj�Yz�Y��(��{�g�U,��2�e���M!^�U+ŌX�H)=|�x�5�I�&�D;˩=�{gY:�?s�J�#�s��\î�Zv�2n��~��{�<+⽸8F,���6;):' 8i��`��'�/`��|L�n��x�����5��j����� L�Ig�~�q���Sg��e��o�?����;�쪯�����g�ñ���g�[X��Ϥ�׆V�`ắ���������K��	��s�@/�̜`~��t���7:d�`�X <�	�����"��9s_i=��4����?'l���l��(6e������km�	db,������^��ek'Bz[o��>��J�VLn�`aO��Y/�U�UO#^���Bږ9�E���u��ċy�cR�Q��i��������o��U��Y`�0��YÜn��Y��0�c��K��3�O� �l/���r�Z���R�w���u��˾�`'����N7» ?�wHy���~�k��	 �e�3��"�D;?�m�Y/oS�� ����𻣨Լ����� ��?�02N����N1�+��s'^V/_ur�\�0n���qw	�ͯ(��Up�wJOel��e9�7��hQ/[s��Tw�������8�C�<<�o>|z�m�O���?C��ǟ��z��>�G��xُO����=���{z����Ǐ��?��PK   ���X`�/��1  �P  /   images/05f650cb-cb4a-4256-a168-b327b67eb2f6.png�zwT����ke�ā�AADz���F�P�B��5�Q�T�P"��@@�@t�^BK"Aj !-�=�o�[��w�u��ho8����9g?ϳ�w����/��� h���!h�$my��V���vI�����KA4�*����8>T
�s����C�U(44T���~A�?ܸ��Der-�!ht��{簬F��١�+��
�폌�TtXjC����ѷ������o���n�щ}��M�^x�}�uWͶ�ߔ��f�Ǵ�;n�~�Q��W��z�4���xŏ�C������W^�MZEǰ�1�{^��9���Yne[7�A� &��{.���u��}[bwI=�"�<n�l�lܨv��~�i#A77o6���ɆL�1����'MR�%j�&����!�4�UF�u���a��U�(��HNU/�"4���`G��dN������z��7T���9��\Č�ق�=eOu�Z	���Rl�ƚlGXYQ)��oVu����k"qz�g9P�4��x�T�ͳ�5!�U��i����#�-s�.�	�n�#�o�P$|Ek웅ĊKoE���K�-;᫞��H���f���0V^Ϟ
���J~��d�5ۙH�^��Qɿ=�Ƕ�%��V�._�|ǽ*?ͩl���-$n)����.mY�3���j�q�0�6��Ŭ儁��HSH$����m�ȥ�Tխ�'9��U���`�J�G���
w�(S/E�4��j��,�/��ˠl�����1��P//+n@�:�TБjgP1y�q�A�m�Zhs�03S��k~ק���SM����~���)ű��ٕi�A�rr������a��Vi�Y�v�iy-L�KTD0��B ,a<g��~oBnr���`[�R�2|�vQ�%��[��f��x�ӳ�/�D]q���;3�P����̿����b���0�jy>i�N����OX%���D��5�Բ���F���SI;s��Mv�qV��.mۘ�/"�,'��ʸ�\h�.C]�����i�ײ�ͼ�P�x�|FeS���K�f��(
� T#'9��(ٚ#uΈ^M��C6��c�?��1�4b���?/��V�*�c�h����x9�Hˈ2�l�1:f�C��ժ	t.�`���8'rVs��ޱ-x�%�X�_��ZA��>x���5i��©LU�
�{}��X|�H�뾒,���%�U�K���s(�������2}����:Z�+
����*s��,
���Yl�$��F�~۹	�2��	v^׮�s�ά���;5���&�0�+"ѥ+rm�ӑ��1�^J$i��1g��1�n���i=�)�T\?�V5�ęU����(��������öfo��dG�%��mmsk�KW�dii.����N���^�5�x�$���5�Hx7Eֵ��<�w	u2YxC=�~��%���F����	��e)�I��~�w�#"[�u;[g�C��z��ZL^4��Z�V��v�w�㬚{{ Q��/��5�p��_gp�0a��9����b�4S$C2^�x'��DbNg��e�w��I<���I����n�p���ˢ��hsl�W����!o��s�����)|�OѢ�t��؛�a��ţ��U��y�>�GzEN!q��\Z1L���|�O�`$�I�BɆ�������{&T����$x�*����V�dڄ5$�M��Dko�tD��)C����!�5ʘ�@aK|�ׇݓo��.�'�񓪮j�1��6|�x�F����G[C��&e�~�]�R��R�l2��};�b{Q��d<:J��Q�}3����mk�
���8���9��<���~��������o1ϊ6C�n�2g�!E>�GsD�?u�mN�|�1;8����jc֭�p�����Kn|�{�3f�<�SD�7�J�jPZI�Sќ%h�ED�M��+똢��[���,���� t| imj��".�_�iܔ������c��㪐J/��ƻ{m%,�̉Hw`n6+�G�:�NJD�t�U}B�0��Z}#ҍ���q޹y(��!H�'s�6�L
^�zc�#���^	�n�Q'���_�+��W�kƌ��cf����,\�����p��N�[�����I���Ss�?ݵN�I�o��I�I������j#ꪸ����&�m�?�y��)g���|�|?:�+���*�/���8�6�?���J4����SS��5���x�N$V�Q��q�!���s�dǒ1%�48����t���J��0Z�PfbvD�Q����M�"bմG�2R��#R^D��+刾E�Um������uA}�I��
�~�Շ��S�u0�u������!��d�n�Q���7����x�|��r�|�ST��kO�d��pf�G����c�'F��adyH+y;]�Q���$F"���o�ܟ�Y�����ck[\;3�*x�X�d��VDVQ��mz��4����A���0����> Ph#M�h�ī����t��[�pQ}���YY�H��EN�����n�p9�l�Q�t�sݦPM'fc�)@bc�R<�@9�?x-e)^
��-e�^�)մ�{���4� ]y1����"2o�@`7���xZ��R^y����olP��_@[I�W�K�y�)ZNx�����^�W�c�(�����Ʈ�'6�Rf����.�o��
�5!�e(:J���׳��VK�;��`�;0�[�x�aҊKG�V��\p���n[����1z	���z���i����/�Vqke0�J!!⮬�r���CJ2	��QNG�E�_J��l@#��^}���C�]�k[�2����6��]隙�x_��`��$�ʿ�\G$�����X�f��I������Lq�H7�>�D9A��-�G�ٺ�g��Zi㣊�� �3�[5�P'I>�ּ-�s��ӯ'$��0�ϓ���quwg�����j|=g��!��iy�bf|�m��/#��f����M��*	�c�-�=�v�_�R�\�@�+ŧӳ#���=���Zq���#{��	o)

��YK3`G%	�<��2	�6(݋���|tߦHs=��L|��N�>9e-�M�&3���4�C_��쭪
-+���rc(�^$?�Ɵ7w��l��$�T:��{�=G����Ҁ��ŝ�Hn�@·[
_w<��]���%�65פ'��oA��1�&�.E@P��#�ed�u,sǚi4G'�����oWL���}r�Ї;w6ut��R���������T�HGC�_�g�����ltԱZ\�>�tHH�Nir���tq���gE�t���~�������/�o�hfn��~VT gj�������Q��m�����������QGY�S5�z͏b��8�흧���QȂ�/r$����|�x�%7��cR:;��O�<�o����C��jb���y��N���B'?t�Ė]]Jq�R�Ħ�`��_�?���+����b��q������;[��ߚ���*�:g��[��(EB��f���dXF�iA_mT�w�ؙ�&~,�p����	^�8a���^��뿽ɥ�X��(�;�`l�-匬�O�X�H*|�������[��~�S�b0�{�g�ϸ����%3˧��wZ�U_�ѵ��df��pE�����K��e�]c��>��N�2e~�B	��,�Z��ב�2�����쮦�K0E�3���/�D2��������/�w���>ы���˾�j֮[:^�����9�~�{f��d��������A�����wj~Y6��-�jlg�[/,���覹�<ԛ�U.��V�t��W�(ڱ�
LyP�N�����H:�`W�?Om^5=Ë�P粤U�
�JŷJ��4¥�)޶TbK饇�⏌��h��ԔR@P���w������k�[oę��R�8;��+Vѣ��?VYG,Q[���ϟ?G�]�啜CU>\��͢5��S	����LϺ��U��uz;a?�Ϩ���L�Is :j���c�SzM����`xDطXJ��J���J�\"�
�
�ʋ�C�#k��FY~��v��k4�p���ƛU�¬v]w�IVV����Wf�/��������t�ʼ;���ã�-;���|	�OXg��r��9^^�d�Ou\�6О\S�=j�.ѻ���B�ط$n�9ԫ�ѝ*���B
������H�ۙ�vmrM�k?�L����[��k�}Q2����i%�����������A����L8&�Kg�f$�4��2n^�'�\]�z��q�ODw����vd�eK��t�ҵ����l����o����)��̋I9�sM�&'�$<�����F6z�.l�|V$s�2Z����u�k[��6�u��ٳ�S"C1h�����_t��A,n����Ξ�R��Wk��<�_����r�y#m��� �:��2^GHq�ձ�y��H*9-9E���:�ʚKM�VH�J\t��N�#Cflo;<ߐ�r��Z��~3�e���i�u�C�+����a�^&��@���c���4�'������nW7hx��I�*�ek�p1�y\ޣ�Zrڥ����SW9�fy�{���#l�	�a���ʍGV�Ը�m��T��jL�O��4f����w`���4���'"���S��B%׵	�j����{���J	O��:'6�|�|*���h	̧��o�c�I}�֥1��*a=�?�#�}7=5�1���f��v���h�0��1��t�_'�5��jd[�^g����N�H%W���D�U��=�=�S6A7�\@�S^��I����X�5�u��.'\�G=���x"��w��n9�|��-j����ʫOfٝ�3Q#�l�9DW��	J�lX�����'�N��7|L���K���)5*��S��蜜����$؛�ܹ6�A'�ezx���Z�m-��z-;�&G-`�A����� ��*�Ls�M�����U�cA7߸��R8�Jyl�B��Cc̺�W�r@���/���G��FKo	�<���? ��N�E��H��E!��V�XZ���<ҏ	\Y��x<j?�n�ˠ�	A1��BZر�y���ň�	Y��<�%	)i�w؉z��B@؉)�����W	5���@�*n��@m�@t��%>pu��Z+��ɐ�����Y�G��t�Z.s�5�I�Þ�/�{%�h���ex�Y���cd��w@�$&'[E��a�*H��fyT~.P��" 3��"e׷��PE��J�eI=�{t�r��'�Z8$.����!�^��Ō4a��&"��d��if/L��h���W���8��9��݂9���0�)(�r׏��?m�v�ݲ��E��_�f԰D.�g�;E�z]��w^
�u�W�'�=0M/D���%����э�v�y5Ń�p�	�'�WVW�Y�R�GF`?�SޖLXP$|�2��%ZWO���C��6����.KKyM����[S��t�];lj�rkm������K�RX�Yʪ�oR���,���Z}�'���RO�ϕ^�I���s�;���.�ai��A�LJ�)����%��[��T��QG��z�)ޗ2�>�c�.�.El�>��;T.��=IaHlfȒX�賌\J%�|�ر2?zi���t��홨��G�����s;��ǉ����d �w��R �DDKaYʨk!R�蚋nM��q�vOI��`�IE��דR�p�X�p���)�-����B �{!<�yƯ�;#�H�aEP�tU>�{�	�i=[n,�n{�0�5��4������Ŗ�8#T���;?<�Q����{P�3h`:l�񢽓ࣝ
��"���J��W|��K����O�!g�9I�^M��s�h/�|c-սz���;"Pc�ia��x‒Zk[W��wQ�fۧ��h=� ȣ��h<���lA7ԱjF5�a�O}�x��@u=��س���@�(W}ҧ�U����?선,��a܈�^��� �J85sc6���[�*�D�nw�1�wow".CMA�q�I��'O�Վ��i��Lt
����h %��M��`���o�N��c"��;� ��:1Y0q���gtw�6X��]ǖ��ɹ���e�g���\�{������+
����2��o��,���9���z3V����VB��sf'��p�L�����b[� �U�iX��u�X�ɓ�+���Q<���O�RY����<P,�>�X�Щou���_��Ck��.KY��ڠ�sM##�X����b�?��yJ	�{`E�/��w���X�D�X�����U��w�{�ck<%4�V
K�י^-E8酿�yȾI�5@Ғ��8�]���R5&
����A -%��bK\�����|�SL���Fe��Wn�c���� �{��+v�1ɝ�2�Sz�/�X���i?>sʲ*+V�/�$*rXK]t�O8vD���X�z&;�7��!���f��.�����k��,ż�lj�\;��x0f�X�+a�{�$��Bҁ �������@	*q��ɤ�t������l�~K�r9�4��*0ˁ� ���%i9�,<���p������[�1��S���^_\21�&���a+��)�y�;��]����(�'?7�R���]��&BL�N��e���K��x�����O8]^]k5V�����U2����N:���չ�yف9k��)H|l�;�H>���%�ef�`Z���9���3�����X7G�����9]ζ�J?�X*�}|&�N�)��7�bvqq@4ڍ���ݤP�����;�j�S ~�@QUUZ�&HV�*�][��u�D_y�@f0�B���'���T�'F?_H�ZX�Y�t�\8��R���u,o��U�p���t���U�cj6���ܖ���V5�1+��C߂i�.%��%����n���E�	�t�[,�s:��'�� e۪fJ�KV�&��Z1R��T�}�Դa^�r����7����҃r�:��X�R3i*��d��vRZ
[g6�Q���5���D����޽����u����6���|�ٲ�G�Q:Z��^�����eC�7Mͱ�a�K� �� ��	x����,\]�r��/�ݪ�9��e,v�����^���R,sY/E5�<lAa�f ��@�u&G�gG,��`O '���ݍ��x��b�~2I���?Q��M}��8e����'۽�J�h�������-!f���*���ˮ�bl�����(��=}�
װN�5��r��l�ky�HHb~8���
A:O.�|+�a��I~�����&��[{��B��u.�3��j��+f<�\և�Ù���έ�G|�yWu
h)I�sO��$Өw��C����;����ѡ�{c���;'����uc�5)��Vs53������\X�y�HZ@������:!�����5v;�L�I6Y�u+�9ft�̦\s��\��잘l�*�T��>�	-���B �����#�&G��>�������v�l̮xR��ǆ����K_Ձ�}+���W�U�������@�NYQ��k�j`E�WZK�1=i��q:RN)n����H�tiJ:P�zᣑ/P�y�G7����u�ER���I�N,E�Geh�/R�~��v�����P�S���h��	����*}��Q� ��I�̉���2u�ku�O�e��6�ͫ�/���I��O���{���Ԍf�ϥ��D�$y6y�G\A0������ӧ��"b<r���^��J������aAu���8H@NZ��+���� �4��Ҥ�ZM�2�K��-���:iR�n�4v@���˽�v��*���o~�0���%б'ݽ�/�[�&�o��������}19s0�+���@YSZ@�E�7��oR��Ջ9$��L�C��f
�'2������6�vxmM�vi�4�������%�H!\sŃ�.��f�M,|B�̶y��}���ie��>�{�.�|y��yـ���
�}�.)��w���������n��ݳq����P������$
�Zᦙ�HOOWR#�Ck��ټ�Pu�]܏3m-�j�9�,��\�]>�_����4���R��(�^,4G'�>15�1��p����\�n����?�y
w��O�a���rכ�G�7��-�?n�%k��-d����L�矒��w��t��y ��� /����3>\��4�����5<������r�o���+�w_sv/�/,,$�v��w�y�\�����/z}{�`���7C�A��w��őQ��R�B����O�U5.�*m��L��N\$M}j��i5�� �k׮�GԖi<�%b?�^�����.��'LMM�Q`ʣ_��˫��K[F�yuȃ�ѡ~����1/iSK��>}�Ժ�;<Mxu�c{;-NNk��#wi���� IÏ�*���T

¶+V�������g�AѬ��N9�F�8:������դ?��&�:l�mh����k,SX�ۧ/���iɽ��7�`��r�jK�̥d;�%v�_ĩ�Pa|�?sͅRр��PTJ��:t֏�@��嵐���$z���RU)w���|�Kr]�k��1v��,"����fP��B_�mM����R��r���ɨWI��T��Vg---�_"E>�K�*{�����i��(7%��`<�{���Ҿ����x�yf�'�O�0���?r�i�:�J��_Gg�C X��-T�ڰ�:/�q���tqk~���a�E�o�˫4�u�~�����d%uV�����z\�sx� ��Pf���SeQʴ>�x��ȣ'qu
��x��iuӣ��u��yt�/Ru;��0Am�[����蝣�(&�|�Ė�zV�'�y3"qwl[������VC��^�.�|�PVy鵵k�"_�~�S�Q���dy!lg~2���A��v]}b޸��D�L��7 Rs����@a�ֈb��Y�)���o�[�o��)C��1��kT�(_o�nn�;J�'u��v<v���Nm���Y���(iDl{U�]9�-ă%	���(48����W~a	���Qתr!��ƌ�8��'��a��/�3g����QC�ݸ�Z���Á��*��<�v�ك�bǢƧ	�͉ւ�V2���f�0^!�V�w ��~�k9��վ��n!K}d��+*��C�p@���L��Y�9b��+� ���)��i9f��rv�.ʔZ�`�3�+�E��l�Jw�^E���R�}�U�)X���:���c���؀3��8�/�`��d��{'�>��b��s�E���˴��V��XB
�͏t�6`fڭ@�M�q~Fz�<���2-V����5;),��K���Z^z��	�sj߱h�Tܝ��P�(����\���$�4x�}F�L�t8����=b*�޿Ֆw�����H��+'''u���à+3++ѥ�-�%��%w�{�'x�V���6<z�r!H={���~���#hgyo03�L-���@��������*�	5_3���:��dL h�O�Ȫ'R"�} g�*(lY5;u��L?m�`z�ժ�N����(<�<�i��XϮ��a��6���^q#�c���,u.E��A����R����;? 	y��sCS��v���k��ʾ��-�Z���9�RNHH���8t�;�G��0�2�^DzBJS��t�k�/��������GX�M�¡Y�ʡ�ȭ�=�E���:����h8���6��>�Z��l~5r(�~@���z(�/��HMi �j���K��̕3�c�w�O�TK�Ǻ�v冗���RPaNmS0��sr6���1��Ws��X����|Z�b��<8c�3B�@�^��M޿Ȥ�R/dG�Ǭ�?9�ә3M��hl�� �or��,���T;���|>�x�"\�\��C!Y�U�l-2����_|{������s'���.��`��*)ͮE�����~;w2xHp�d%!"!{�(�j����DZVا��h��ﶤ�X�-*��������U�a�t#��8�ؤ�ac��A���M��;����?b�P���k��{�2�O�c��J���P�.S�#:�Ԍ�XL���X�^`�]̈���~X�V����M�7=��3QD�Ejǌ�����������Ld�q�C0�D3�ٛ���!I�^薁��9  ��U�2�%pN1�o{~�1�K&�$d��k�m^]�����<Cty�����N������CX^܀!Z����%d�	X�e����4����@��9�S�@��I��7�y岄x�Y�p-��XC�-5ԩ�6r�����zf�3p? CF��G�&�������t�����6 ݳ�a�����/%Le�7����C��D^.�w�9�P����q-a�����+��Y9�\�+�뛱0#6$��M����f�L$� �h�0(��I��g�I� gdU9`���6�3�3�T�}�6�i�z�����YE?j��,���x�I�����N��y 0�	5�K�VaQV�ʠ�(�XRu~Nzhw|���Vlt2�b�J��o:�N�uБlI��s*Ɣ�?_<i�*bn!�2�d"����X�K�m-O>��1PPk��/? W��|�d����ڮ��Y�92)��lڿ{ҿG0��	',5�6{c��vO���\b_�KYf���DN�� ��S�fQ^����oVf<�II$� �T�bK(|��#���sY�¦P[R�Y�*���:f'�Dz�(K��ULx��Eu8ڮ�m�	�l�r���$|.FY�ʪ�n����\_�3��3/�'�V$u�B�M*{@���Y��$`,)����0N�j�
��s;���0�S�`n:Ժ�U�ܮE}�����/~�Y�i�2�d�����I}��V��n�bq�
~�=s�&M���`� �-4�r=]*�</Mb����$�h�uNZ����;9E�]C�&��e�*F�O�]��C脻�Nt�.�Db��D.�S.��Q��k�ǧ�V��,pN0~�N�@����b�I*VBsC��ЕϏ����K� ���Xz��
��dR��L��3M?+�x`�}���׾����C�J�$dΏH`��7.0�!�^Qꤐ|nU�ݲw�L��sC9��Q�;�^�uk�3���:=�/ǝ���Z��m6Έ�|X�-H�7�$��� rg���M/
B7�>�-9;Sw�0û�=�d��HR`�/
�?
�Փ�y�B��{ǆ�R�`�x����=<����fƎ��M���3 ����[4Z���HϟM�y@K\.2q3x����Q����������F��I���EL~��5l=źl����%�I�4ԕ��U`8�z�5w��d�&��S�%Xܳ�Q79}�js�5��h��U�aI�-:y-'����܃D��g�Y�����[�"j�s�|�Gm+��nH5���;D",���9JC���h����Kp���Hm���Ǟ¬��w�mB�����c� ��4[JFrl�e8��͒@�z�r�F�\XR���ӧ��K-$t]�	�P�hiJ�l��u�jz{\)�������q1ۂ�q���c�=�5!t�Е�,���f�ұ�R"�@�"i��_3��氊p��L��Ͻ\] ��t�֧^Z���mP-`����9�a���{l�����v�_�\�~[u7F�`�خ�3�b7�������� %D��;t��xy}�j
.
��Y�.�)$�D��	�s�޳=?��ޓ��M=C�7����F�-���̯)E��)��
�j����R�Y�Z!NE��?j�-�R�����6�� S��ݰ��;1+*83OIV㉹���)�v;g��ˢ� -�`h��al���X���Ě��o~��t�,Rrè����|7B�~^L7�/KV~�YՋY|^�eچ��h�[���`��������^�"���|*��V��l��R�a�W�\�mT[�A����y���ݓ=/��"Mv#�nq[�K�GӴ�Ն/u�������z���J��]ޭW�Z�_��K�6<�M��b�����>�#k�r�y����$8�f�M H%W�dns@?r��D�N�n���R���+#jX��\��� �lv �z���@}������a�X{"Iu_� 1�<0�<�7j�=�5�tr�z���|�6Qh%7,s�Z���?��/�k���c�Y�3de������-�^K<��\��s�-�M1F;P�5�t��h���p0�_�V���������}	ݜ%�R����QG4�\ON�ͷ�<�A�}�lk5ā��{`ƶT1�	�$9|�&dV��(s���	�/#��g�s����I��I|���y��p��+T;�O6.v�g�IۑC_w�8_�p��sM�$��ݻ7���4!����Mv�\;�_"8������f7��d�)��+�����NIJ�孫�e�1�h��"i���T���F��diV2#8;�)WF��x^/����d���%*%�B��}u� �y����>�1����L�1�����%#��r	r2��������}6�_���g�CohyyY��|�.��w�b��Ws�u�kM�3�Ctʆ�EҊ&��'���L�1�i�,q���&��O�	�3����r�PK   ���XG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   ���XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   ���Xw�'<�  �  /   images/0ac982bd-8891-43e7-be61-3976077ece17.png�YeTг�%�nda	�E��kI��^b%��K�������.i�F:������9g�3�a��7w��U��qipQPP�d4�I�?����w�U��8.
n((H��0�o��?%5\V��l��p�F����9ٻYY�Xs9��f�Ҡ��~T�����:21�B����l�1*�(WH���bZQ#�,Q�Q���C��T��DA������I��׃q�t�}��1X���PRj$�km@���1qd�j9r��YG��]�~�Y���WX�z=[��5ҵ�� �G�2Ǧ&��PI�c ��p2���*t���7F���3�7!���X �R�Q�n���aI�2v�̩���A����99��}�w�ܦ;9�l>`�E��8�������Yz��a��O��W�q��O����:3(a�{4
�u��Wᵋ&̪���F<{�j��kr���[���mUY��KR�x�P?�%�^T�H�m�^����?�`�D���Fm��H�w�⡂s��&L��B;�Ґ��oԒc�MR\���������![����Mb�'�o^u��O0��'� LP7���9X{^�=��c��m�(SL�clv=���п�-o�I���QRּXI�)��A2�v�����?�jj��G"�Z�\.gۻ�)F}{��J��� RΥ��b�zL(�;1.��>	���Y����^��cD>�A"��f����Sz]w�m��a����8cAeE�ʽ��8�+0��Q�
A��*2�<Q�b0Rz8�$5�9ˣ�U����t��/a���F�$���>��ăU��VD��aa�}>	v��
E��幫������m%���iW�:��	o=�{m��ڜ��X�z��T(�^�xPG1�36WA�h^����aqly���RY�?�����Q�1�LFv/(]��|=��jg��X��\V#s1π��ļ�*�D�]v�o:��K�<h�^�Ә��nO�[��
�X���Ɏ4pc�8K�S�p�[���*�>�;$	j#C�0�'�,I��3gIi��F�U�E�k]wS/c]p�ܜn�:P��8�cn�0�_�ު�T�1�Sa���)ۻG8�,:�e�PQ�ƛ�Pd�:q����B����U{`u�g�`�Oq>29�h�6����%��9�4HO���7�(�_%)#U'b�GY�O�:�9�W�ܥ�7��,�]	��S
�2l��|��z���]���^��^��Xß3����f>�(M�r�|�5�K�&`�|�v���Vz�Ԫ�^m�y^�
��U;�&�����&�U�S�'jϧd��=�ڔřQEh�%�Zfp*q�TTg�`͂��K.]��ǭQ����1���䦭|��&�Y�o�HĈ2�$�ѽ�嘅*�<MJI89���9�ֿˏ�X��͗5�������Q���Pl����}Fn����Y�w����雅&�|*�V��ee\������#`K�7���di�/@�H�ᶗc����� �2f�qp vug��>�V��u$�*H����Қɕ�����n]��5��*�Lb@*~�Q�Ah� V��9`�j{��
��@N<4���p��*0�r�y�J۰�1� �Ef�pZ�4d�f�5�L��F/�V�@�z�.�SLeC1a�H�ڍ�B�������~���ݠ|A�� L�Tx'l*��GG�]�!�3}��+Ղ�[����<�s�<w��4�-F���"w�J�\\�!����Js��x�;�t��e����O^�皈����w�f�d��/8β	{ύ�IXh<Aͧ]�"��[՘��Y��n�?�c��ގ'�����$Q���k�u��J'z�5����'\�/��}M��[!����@��my�w�v,�d8��t���zrH!J��/�8�9ɯ�smdN��<وD�a+E��x�0���8f�����c_����n:c}��4�``b�z�
���b�D�P���L���@j�R��k��q-�O[:?�)��+�MD)����tG�X㾕�D�]��2ڟ�*)�Z�dxy۾���(v4==�,���o[�T���QbE`TfD1�Lfm�p��8��/{;��Ze�u�s4~���ī�������uO��cno��o�OX˙,p"�m~��496lNRU-��go�`�[�G�j��3�az�|1��6 1����t��M�+���s���Sh��5�?O�~'�v!L�n�p|�c���@��ޠԟ�g��P��7�aY��]��"�P���[f_���7H�\'�2�y������pM��d�v��NKѾ���<��$��6E��#�|o�t�7������v�?�N�򕋑)������(��̑�{�K��V������1bM~$�ل�*A+6=�͑u���6@gN�ԑ!��g�"����Nh��b�4��r�5#P�>���g�4�ӛ�q�ַ/B�z�a`o�6<J��*�mt��"6����N���ö_��|q��/g�1��M��l���5f�n�Vs14X�,,�l��F·����S��})�v������Ppy�X�:�N�E����%��&/�i�l�����؝>�~��{�=W]㉞a;2S�1x�G�y�M��|���U6�-�H���]��ơ4<+v4�ae�1e'Z8�Ύ����~ȿ�3M6&��t���$k��
K{tg�X�l��o�!Fd��Ż$	6丌iho��7�����cO�P����J %炏�{ 6��Z����dSk�W�qO|�:U�̇�	�߹N:g<�JO�g�e߁�{��Jݦ��UBD�'������T�������䆘,aI*է���^��Cn�<� Oj��;Қ���bU���/����WE�t�M[aam�����޴QY�v�ɧ��8|~�L��6kI�&�|��݄��ز
�[����4�l�۸��9/o���Q&�ox,bOK!:�ՔzX<c��IB`	����Ѧk�q�����N�|�Ƕ�]|����4�����jx�=���G�݇��_ϐHU'���j|��Sdot>n��Zg7Wl�룳@��n��`.wR�vA�gwRs�m���
�E���~��2UDMjH�2:x�Cӵ����*�9���E����dɐC�S�K,66d�!�1���Xp�qS�#��8����1!^�,�̞�)��+�0GX�`Do��[�w�k���*�Ŀ�v�����o��*��7�R�-���v��gj��e��#Q!~��?yxW����}�����&��֪����CA�U�%O��F���-�E��a���K��Ծi�q�uS�f���G�h>�*�1i���
C��L��&����zz��O�+�/�]}p��m<<�XfRX��'j)QL�3��	������:^tű�q�*�PQ�I�0^B��l"pp@P���,��-Y�죷$�7+���Î���a��SЉ�vb\7���a�#f�.N���e�G��L]��$7��Z�m���2���Y����Xf��^��2�hT���(��O�)�%ԊL��W>,
��&��dm�{�ew�>��� ��e������ǅ�m�qF����{f:���l2�$�vf"kb�C�`&;`%�����"��:��c
by��C��g�����´<�]��~2�o{ ]�/�(u��<*��~ �e5��D��6�ng��}�~�p�D� ��+Z��N�f�>b�F(qGg*շ���s�$n��5/�������Z� ����҉�ٜ¥2���1�E�����pW��,��ߠ���n���[�p�Mx>��f���xd���$P�a�q��Y��{�#���M����oi@LnU�U�b)��՘��_lm��q00tX�z��JU�6��[c8��\r�U}{�y6�awp�P�Q9���eCe�F
xD K&Q�'}!TϦg�����2��o������ٚT�u�G��ő��/"�2�5�F�e2�,Ww4b��e��k-K��7,�BM-s5�/�&d�Kͧ7�\��c���ù��v
�޺�iI�.��Z3��E-'���_����'ٔU���*�� 3�{��!�
��w�L��X��
Ņ�!8xO>]�ԛ@��_o�=<0���%������P�ph�H[��]k�9�:'X��r��l(N�J�l���AQ�Jd�qjQ���YT	�M>��>V'Ts?ܫ�\T�s�H�Ǻ��"vʛ) ibF,�1}�NR ��c�}I�L�C�Z�P��P�MR-?=�qP ʕM��*P�����}5��TG'�9�J��ᐒ��ˢq}V��6܇蓜�C�aT&5��2��Ut���-�#�8�m�؛�)
�|zMP^ݤ�;�+���ZI}�������)�u�,�3{��{uE���6^���p����d'�	n�X�e�~Y�GT�b4y���y��4�@D�e�6b��%����r[hH��7�����4J�67�D� �;���� 
�G�xBm��z�o����8�vp�s^���U�"���!}�%KL��c)d��YЄ�����6�.?G9|��0� ���f���ޜ���u)��ڤ��G,U�:n�T��@4Ck�.��b��#��D
��EA�s�s%(��B6G�s��o�x$�!�!�*eO)Y��N�٧`⛉(>��W�F ��A����M��G�f�+�J��ƥl)~~�g��J2C	vh�n�?0���Y�Z�㢾r��?�5]Ei)�0`1{����u3��O�xF;|xE3��a�w�t�7)!"�R��`x[P�^�]������"2�v��Vd�"���=����i���'<��MQ�Lh�11��Hb8fc�3D�j�,UM��1$�f #�t��1��>��P��|�oZp�����|����Z��@&����\^����j����F��a�+N��aq��%jm�Pt���p,��@���)�)�ʳ��戟6���I�s[s"�E�t=쁮7�{��X_����1������O��I#���k�W!�^���
#�j�c&�Qq�I�ʳP}��C3e~�dZ��E���}LH��	�΃��O`�j��*�MA�߿��"�r�I�CzS�~Y6M�
�7�J����n�*�Y""�3�L��K;�V�(����M{+����)Z�%�Jy�ȣ����T�M��{�ai3�Ǵ"今K�^@����V��(�����/�-@�5���5�a���CD&#�'Zkn��Ԓ�jf�z(�E���o�wH��=�RJ^��������V�9�h�7^Znt7�"/����F�6�o)WlH�*���Vx�3���%>l�W_�@Y��$8N���e�Sw21E52��g]/v�	hy����c$�9{�r-4�7���[zw��:7��7/�c��,e=9L���Eyx���{��ũY�H|h/�
��0]f�(��|�PX;�����zU���w�%�}<IZ��d��0�;�me�z� ��/��̈�2,�n�3����ǟ�ا��:}�E��a��1��*���������,*���cĦ�ȋ�ʩ3������S�T_�l�p=*�UjY�J<SI���p��yZ�5�����W{|�\	✡�o��i����>6�����a�W{��UB�H�C�i�� 0�Eg҆�rԼtf�h�V3	���P ��?����0�D�#V%��0����~@���R���ՠ��b�v����w-|���Y�l�D�@i;� �C�;W�T��c-��H�&Aެ���6[�f*��}�Tj�7/K�S��~������yI@�<�^*�y3���8ա�^�r�\s�w�z�I���&��T2�ۓ����7�����2��`�=^�X�&a'�^��𼓻S�p��/�n��v���ˠT��H�qi��#�l�ŝ��ܰ8��X.gr]i\����E�~��z|���	����l}
N�	����Ki����V���u�hV���^�wv�	����~sCM���
cb.�����"���(����n�ޢ2Ck��l0��5��Bt*n-I��CFR��9�i`���C���,f@��'�C�̲= ��į1�$���Aπ�(�y`��OJdD�q���zO�b�Ot���,��=�-��EO�޹1��qa)�򞑧�)w���ٍI1O�d�##����rcǑy�u$�6����)퍭:F�5��и�|�=��8�դ�^�~�К�!%�IZ�$ �ز�W���52��sm��fx�#.MKw<�ǓwT66����0E\�k2w�r�$%{�p�B|������b�>9��i�nI��j]�K�}0ߍU���[�yTήzM=�y='�� `�ӕI	u`�r*�[�R�I����ߟ|)@Eirx��4 �я39¡ۻ6�.((2�;Ȣ�3kO_~��i�:��e��u<��u��b1���+��V�$�hUh�gB%�B��ߙ��ǧ�6�}4$Y�9j{1*��m��c�@���&��,��u˱K(tqbV(�6��������Υ|���]r��[Wtaq��Z�d��ی� ��9�U��N��,����uy��-���ȸ�����E@5_?b��A��'��eun����}��;� M%�9��k���z�:�h+�̟�w+�-��t]vh��UN}�X�f��P����Xn��UZ�M/�F��fn���9G8Y��PЋK�]�G�oւ~�8;e,�=�>�Y-����3�l�/Q��Y��I0K�mL8�ķ��W�{��^��L�A��&���u��k�:V�k�@	s��2�-�hm�rO�Zܺ�q1�=��`�HkL������=�D￫�#nk��f�7?�ͤ�|���/��6Z ��g�y�1
�ތ���J�_����u���Υe�T�Q|x~�ՙvm���})����H������qڑ,(r��Y�Q�R�>�lrϋ`Sg�}��Z���+���o���ׯ9B��V��2;|=�|���m����0��7��V��d~��]�)��V�˥�0��/4�e�BF�� 3o���C�~��'&�����������=Oѹ�_���<�h�xh9w���A/ٿ�ޚȟ��7�)���ş��G}P(qt-���uB9#�-3i"V_c�"�S�V��%�C�)�����J�V쀵Þ�Є2�If��Qt��]Hn|0��e��r�c��#���5I�L�����Tn�)[�o��]Ჲ��f�X��)b�3q��T�#~��[�*T~�1���=n)7R������ë->�R3>5��(�*S%m�?PK   ���Xyɜ��  �  /   images/110f4c69-ce42-4daf-8800-65b9db14e3fe.png�y�3���tQ����F���E'Z!����� !8D/�[⢝Nѻ��{��|g޿��wgv��}vv�_vgg6�P_�����DKS�:��� ��bJ*�����K�����������I:_5sߗ�N��0(F@@����[���^PAO�s��=c����q���W�AO�]{����s�|ǋ5���5$��/�}�6�av�B��0��Ѷ���*��� �mik��Tr���ArlIڥ�z�!��lS�I_������i�|�J��?��!�����"L�L�f�>M�8�~SP��v"p�_��b��*�i��:�����X*������#�F&~x������NG�2Jr3��?�P�sH�{�>7��<X�̠��A8po���k	l�ʸ�x�cu�����[o�Y|��r��q~>௳ .��P�m�^��H������e�/�����$��4i�80�o���j��C��ޒ�<�M0Н7!���[v\T���D��As  ����؎>��8;E*F�Z'�"�o��x+�G���Ǫ���8�i*7ls���Ef�;��&�f�o.)j(kX��㉉�4��`=M�¬�x�W��Z�Qj�5��.'%lNVi�����ZᏱZ>�O�.��鶭LP4�0��F�}�P{�����m�9��#e�I�NRۯї&G���k���ֈ�h�54�
��ܳ�=ӄNzۆI�<��ΰ �8�Ż&���B�/h�;ykm�|���ks�_T4�-:���Zt]:�U�QL��X�d�M�P"{L��<�8t=�º#�QR����{B�hh�-��j�>�
�V=��d����~�?}���Ԉ��˽���[PUS��H���,WkD |��k]��!��8ex�y!}:f� �TP�#�x��(�l��e.��9�.�G����qy���{�0�8�����y�VN� �t<x;:[_��E׫���O/(�����C ��/�D%��{�&���R�����Ȏ����l�	��q��9�g��0}�)���$+���<�����?��tl�3j�2�I'����ȭ�7�5zW��=��!HG=o�_��b-R������1ߧ?W�c?�&����l���'u��ٕi����QMrˏ�}�)8!�T�����_����������ƅ �fO����1���dG��
Y�jƁf�?
��"���F���3G����G��e�>2g-%�4����!�c��)��rB�Ƕ� �v��G��%G�a��PD�F�/�	̈́Xbz������?���-(�� O�vA��a�{�nq�iGᅂ�_�"m�j�$^�p!ZVgL���T������Nv[|�}NY��(�mFz�׃u�Ѝצ� >��,���svSBy�:�K����e���vx_�JX���k�|-�[��NZ$>����gR!;g��<��6�
���ei_(l�����9�LV3�֜2Q{�(�~[�蕇�Ld�"�gttE\ݞ���mS��bt;�f�&�P�c@NjB��aa~�y�&�����Q�X�
p���S�L�n\�f�3�E���s���'�쬨t�؛r�O�u�f�֩��	��t��:�Ȼ�V�����-��!:�	�P3Fo���I� ��cd 3�Q>��k54Kl�xg���sI�o	%������lJT�'����:�6Yd�7��e��|t-i"a9u��Z�������#�����_Y��W������P>�ɥ�פ}P�;�_)Tu����O;��Kw

%��,�%��yܔ����nH�ʇ=���Ҫ��p���O��,��Sf�F5��T��NOF��NKv22bh�p!q�ؓ�����I�%R�O��Mw��h;���i����Seͯ;� Hզ���Z��N��W�:iֱ��wy%�7q��>du)��b;a��3�y�0۞*�h�������`��V�}�0~��g�E��&�>�vR�_��=PΆ��W�4hiŦ�W��<�̿*�0��e��Vt����aG���.]Rdİ�p��b�]d����&O��U����@*��r��o��G���}~9͂T�.?�0�y��[�v�xc�>�sc�o;sӉa��1������6"?��[m���%�/��1�Xs:o��%a���2��D�w�~�S.Q[���?�=
�KE����� �$P�"j�8��v<~{dR�����j��l<1�T3�d��%~#�`>ߒ���IҙK�q�l�TS<֯x�po���\���׀l�ʡ��D���
R��A|2�jB<�τRX���� 1Rc��R,�mq���@Y1����ݞ/o�?a��c�2�.Q�t{�D�-k.C[������U��.D�,Z�3��Ge����x�\i�OWZ�	|�#�b�@��^���%�,_t8�|]���t-%�1�y��V�qC����T��žډx?�}Y�[>;*nn?ˌW��̡TO����fOM_l3�eg�K,WddW[�~Q�EZ�����FS��,c���g���ɭ	#�F�c�k���-3�����S!n���T��11v�՚�
�T�����O�480��X���S�]�`�X�RU�6ŘF�&^u�	J��1_)�@��$Ĕc�t�P�^$�%ETZ2�O��E�`�iN?$�֖f\Ծ��n�������Xd�hO����!�=�֊B� �>;�2������&M��4�J�
�4n���d)ЧO[����7]�$��tO28��@<FӦ�,&u�������DӺ��F��*?��#��ٌ�%f}ƚ����G�垛�@��pi(���L����@ӀT����5+�mA�ؗ��"t�RCR�o�1�n�Օ���A��_��ӵ���}i.(��M��`ܖ�	�ʦ�S��N�Ԩ��X@��r�ݨ�+|��mg��&'|�D�����l�LW�h�_ז�+&�`�C��gx�;�H��ӥ�v�~�L���k�x0j��8"��>�����;s��,	�w�ѫ9L�vE;��c���n-M�g�O�#�@�k�r�_�φ��1���w�/�~��N���S�f�u���X��[��N��%�DjK�r��9����� C�R��xtMM�Jfm#^��1/\�n�
�Η�jra�\h�1u�F=��O��9
�ʄ��h���~�>os�߫~�'Fw��D�����}\&eE�Ϳ
B%�ڰgF�F�j4���J7����s��sY3/����]��@)_r�T�Ǧ"�7��+`�R���dǚ�$[Tt�II{�\���Æ��n�n��q�^.�E0G���#��u���"z$1�p�а=��-Tf
�v$�&*VKN��Ɛׯg̋��ʹ�o��b�Y���������:K$��@t���P��E��h�+��,� ��P��z"5R�dEm�^�|����;�Io�G�&T�%7k�rĩs��^���j|!p۫��!�`Dn�f�%D'Ѹ����v�	w�� ��o��r�� FT
���7TTj;�@+	9��c�<ϟl��V�W*��U�����M�F���|o���6�b#���T��htl쮏�����2�`@9���<D�U���+o)�b�r��2pV������D^�O%��.�W]�����V�XDu#la���|k�Mr�����j�sG������P@�g�'#[�D��sWR tO�y���d��
�M�Ϗ��(���$+7�i���DmNß#_ah�o�~��h�c`8%���s��?�X�*���	�6�_~SxX�9>ZD(V�J�
�z�`6d!hN_�0�z_"*�� ��#�僖e��
󜳨���Q���C�k�'k�A�N�m8i�����QAW���V�ҷPH �@�\�Z�����v��a<�,A��T�I	h��߸V�87� �:M��N��͹Ji<|�kމ������sI̺��lE�����h,?�ܗ�Ӓ�m�?��t��a�!w�rJŀ�8��Kt�B�A䇋��x/�j�	L%kb}��/# _�7�օi�*[Z�� ���6����辧���������w�맛ʭ ���K11 G�M��G�2���O�Av���Ozy�8�l�\�z�Z~c4`&Tl���/Hs�^*�5xw��R�т���[Ű�n�-6�e�!�Y����z�a��NͰ�A��&��a��-���ZOR�;0�$n1��-��L��!^�)s��b�4�������Ϥ���`)�9z��k���8��⭍���
M��(��_}�ȅ�/OG;$�]����*>R��s
���1�ثq��(߬�SϿ��|���Q���<�T��dǡN�v���O�xQ���n�Y	cx_��utd������ϑ����|�#nd»�����b����r�Fs����J,�WV�v�������fs������f��n�{z���jꂕ�.񾾘Q"j
Z��d*4Sm"J9�[����>�zӜ2�]�R�S_�|��n�I7M$�{�(�M#��X�����]�T�ک��1�UP/t��&��^P3)�%Σ�~��~Y�.e�I���a���|��h�׉s�,� �̅{T!fg���|<����vC�4^y-����@���#1�1z&L�-ZH�<�x�TŽ�����#^h�����Ogs�;Ӫ�Ѷ}��f �CXmos��7�Jk� ��3u��r_�/gz����@�j��s6/�1��^~s�bٷ߿n1x�ɚH�c���$"����N��r�=�.�mYQ@f�lt,=��z��pm�(�x^�*�q�sG��<�Xϑ^zv'|4�+�[��-5����e[HaZ�E���)�*H1�LXpND~A%}�"�H�.u���]�����([��aT䝌�y,4q�@F�m!���<e �S>�=��c��Ml���p�p��~���Ώ�٧ѽA_���"�:'6h"7��]��>�����)�Y,��!x��E���2D�C |�3�������}3bFꢌ
Y]�p�qJh7gC�ʳL�2J��>2$Qk�7��*����V�݉5��	G\N)����p�rU�/��.,g��t��yM���n������Ȇ�
�kp��T(�MRS����+��jo�z'����"?4]��%��Y��N� �a�����}3İ���p�Nd��]�AH�fԋ��p���T�T�������C��Y��F��e�9Õ-a97�����|���ß�p��#n)y �d"uO��R��g�q��اv�_*�_��J/y�k��+�Y
���H��P��'ݞw%������զ<~qhzqzǋXÒ�j�R/�A�W�۔3�x����Wb#K&W����ښ��#L݌�ԛ1d:0�Ov����l'ں���s���g�eM���{4�?�'��Gڅ|P�%��s���T�_�V+�g�-��4�*�q-�8�{��s~l����R�jv\��y���;럘g��|�XZ���z����Cqfo��+�eG5��ځR���K>�m�Ic����_��P<����~�w}����B77�2&5�{���2SY�ONp��Yp�4����VI8Yd�T��Cq��I��1I�� ���ӭ����m 4�(�J3;Ml��o^� YMz����*~[�1���Y���b<o�wZ%�<Î�o�u�󪴩71��tsmO��$ٲ�U�8����\x�b�cWl<��T"T�����+R��"�]&i<���-a�ŮՕ��U��3���`�`�P��8�\
j6�����o���4���S�.�SƌK0���~��/q�>w
�q��I�@�7�y0=~��X�����i5=�%MI�P^���=��Za=�~�����dk`�Q^��$����ft2#/T��_���ihD�<�����y
[,�������T��o��sm2�b�#_^�l�ݞ���U���=���|���3�&���B�H���ľ���':���j�M�����~����k=�Ĝ�Xkt��������̈́��������a��K��On7�6�ӡZ��:s��D�=���������m�A�R3�{�Ղd@d��"����O�!|JY��6����(}�F՝����C�Q~�2j��z.06��A�o@�$^,������t'��Qw�X�^zY#s�;{t7�y�'��s��H��VʗlHEXJ4�-�O���jO�?P�_!Z�%[T!<z��VQ��.Y79��$��{�٤Ԩ�Ι��K�*�*̖pf^�,= �g^�^�f��̜U"3Ъti���Km�B+�?��8�����3�j*$˧��C�ϰ�y�]�����*�'d�V���h�v�2�h�uY�p���H�B/��Y?-^�i��uf�B�q���*��ƽ��e��Λ�j?�]��nD#�K���d�=�W�L4���1��������td�����3���0m5��XB�$KU*���>^$�֫�2�æ���U���+�߻}k۞���w�~ó�O���Yq٨摆M��|������/b��i����8jL�X�)��0S�;4��6����f��|�D����V��7�Y�؟�kk���&m=��� ���� ��2�T��J��fQ�Blՠg'ٜe?��|gF��%���eo�2�W�$y�^���U��n婎J�d����N���|M��D)4P }���F���u����M�=���� s�LN�#F<�\h.��fY��>/��6����%J�+w����"G:Ӣi����,�Aj5����IO�$P`�o�DZE�:��q%�W����W����bV� ?��m���C�@�f��@����4�Jr�^iSt:�Y�X\+�)�]�s7���&W'�!c�I��^�|>��`oْ�J�S�?NQ-��I|��b�]5.��b�l�D��Y��U�w|�_�D+vE}�u70e&�C�3u�&O��ڙ�1f����5�`Z	�)}������
�u8��io�(P��1{m_	\p��*X�RTX���U��i���z�m7�t�:�5mSy qR�����,n�J��3{�X�Do[��p��6�|�j�P�Z@�8�CpVKL�9@��|i��F�jL+$D�^�݈�0����j�^+�?��1
?Q��<����,]���c���V[��/�!%f����Di��;���o����V/{@O�����e�����:؜	�����Z���?PK   0��X�r��}� �� /   images/1235872f-9927-4bec-a0e7-84fb82154d9a.pngD�eX\K�5<����!X�ݝ`���0���%��a��������{�y~��W�?��zU���ՑT�0�H�   ����: ��  SP���a���B��P�  j�џL���Q����  \��=�uK*o ��EAZB�;���*�\Ε�T봟���5�>΍��mќ����3๣�O�D�ENnz�>-�b=+���'2S|�G���17����H`���22q���mD�-�۴�:����V�,��e�wg������rܯ��sڼSTr��G��D��K?���J���P�G����%����(�Y �^Qm���(�?�[]��^�ѣ�u�/GL�m=_w:�jƧ���a,�uXn�ht\z
��QͰ�ߝ���yN�Q��8;'Lȭ\k�'������ɋGG�F��[�������9�.I�>ag�1����KGa8�M���ڑ��5q��_���:�x�ek�΋OX8�Us,8`xJ �h���U�Cl-�i4 �G�{�%�$��*��4}�����:N�/>`��� k��O@� ��YUx=�B̯z��\%�j}6��l����\e����6
�U<!��琮��F�/���,!��'w7]33��q��-�������**Sr��0f���,w�풕��	��C[Ppg �*[0�3WŘ��Z�xdK#8S$�&����/�/��T"�'zd��#_�A?^{c�ڬ��̐���w<$vsy�zF���4,��s��p������|֐������Ӂ�>y�.��;p�!CA�@����E��n�o��Z�S�h`�� !�
 2[J~{;�S$<A�>�@Nq.1���y�b``<�	g����}s":::xUej��������H����< �ns�F=���x:���	��6ZՌM1A�M��C^k�z@����d4��f����H�� �MN�v��y�h !@H���
m&g^��MƏś�����p	���WL�3%��>����|?�Ɩ������H,�z�9,u�q���H#�����\����'��h���yR�ُR�	����}c@�Wغ����TR� �{���� Yפ�G
*�����Vf��*[$�(
��x��Y��s݆N�_�)����׾p`��X��=����O�_��?訲U��Vת�Z<1�,��q��Dl2r���}Y4
�^�60�cr��R�%J��r(�K��a+�.�H�����nm!����X�s���g��O��z�"S���O���Z[���@�W�E�m�&b��tC]��]��7����:��Dp(��4Y=Z��9V9S�i6$��֖蒱���+�o>R+��J�~r]�&����:Z�!�.�q�Z��e�/)a�oH��/t��@��,^���839��73�Kn����Y$/������	���ƃ��G0(��7Ōr�[�߽}Zmvؽ`}S*C���e��㢡}�=6�]6������vzr��RD������:+|��B�C���T���Cͩ��.q��<6��C��;v��7��W-�A�eb�F�%r管�j`PؒS����i���:k�/�H���ܨ���t
�w%x�s���6�W"�R��ɾg��Ϻj���?���0+'���*3����}���[�f�`���H��⺲���I�V$4��6�VKA�ȤN�>"x9x��Y$&��Җ�QN�L'�N"9��*윷�Z�%��������WGgg�^�gk�F{\sp��{�/����^����#e�gs�AB)�9C�_�����T��f\������j쑋���0��R7�C�^,��L���S�׿�ť[XΧ͸��}�l����`�����nn��:�^�@���xCd���p`�D
������<Y��:ǜi���z>=� dC.��a�.S�U��p�	ȍ�$�M��@�C Tazy�
aN=��Lr�=v�3� ��i�E�	��oB�VN]����
%�[�0ү��v�kK0�7�Y_�� ���MP��5M}w;����9��Q�����uss����t�z>C�u�d����)n+i[ �o��J`"�n	���8,.�� �2!M~-'q6������ꋫ�Z��B�};��i�������t�l��Q�d�b(_�[�a<m���<\�[�n쑻�4:�N����os��U�~�8��R�z�*�(Q�Ag�;�_>"��Y��؟Cb����,�Z�"���1r��}R��t�q�3��w��o �t0����'j�:575eژ�~�#�z��<N�/��}�ԉ����������u�(����N-ɔ�i����j?��WL?�w�u<�b�+��$�nO��z�M�ԫ�����4� �^��c��%�Dl�Ԛ�h�l�HH�%�0��iQ�ԧ�z@��1螓�X7oE9�6�@�}�-b~�K��ZG�.Ĕ3�!�������'�-?k��F;}���sR��P�V�mp�En�&2��U*Q��u��t¿��مxDz�4��nΖθ?����-���ǰ� ��4�6m7�������������<����u��b�x�M�����'e�Tgc�ׯ��&ї��N��y�NawS�?�ڀYD�k�\3�)~��8�ߟM_�u��h�`"��}aztv�_�L:�_�Ua��{�
�tA�|��~s���ß����+�q b� EKu3�F�ڌqGG�\�t�6o��ŧnԫ�H�e|u��aNZ�Zh=����8�Y��{�_ګ�+Mo���6>��q��~?LO���ᕁ��u>��SA
����M�@% �r�"š���-nD��1S�#:/�A3���b�|�=$D���r�����[b>`\�훑�I���=�Ӛ'��,q�j�%�!�acO�E��(*6��:s�c ��ܔZ1��L����k���v��u�
Ǩ<x5|�,�\�3	i ���rB���ū�ʪ:߃�xg�]�R1Ύ��Laq�%T�A���*!���J��RY�E�R;�<�M����y|��2���o�R�9Q��.�է����p�I/�V��D�"��ˋQ�r�d��������+�*����\3��>@u_��Q���v7V�B��g�RX��B�F���m&jG���p1N���X���X|Ŕ}�m�ã���!<��1���hK[g���B����u�<r>D:�=`R�7��ݒ�8�
��@�ˀ\@�m.k���i'?xD�)}H W��u��@�籛W$v��2TR9��p�v~����2�Z#��V�Ͳ%����"=3���:��d������|h�@��1^O���~5��w�@m��9�<_Lp��W����<WF�/�k�[ $���W��u=b6�׏��+SHr�F�U_&<Q�x��F�H�k�b�=� :�h�\�(>��k����aH5a���!#tַ�Z�C#)�l��k�%�ƳS����7�6�B�1Ψ
��cYۋ��DJo	����O�ܷfQ�6�, �oH�A����i��e�y53PE�:�A�dwH�A�~n����e�2P���:��Ps
�Q|���3���h�'-�$��Y��nz�B�'�bZ��Jk�T��h�:�ұ	4�-d�e?}�eǼ+���o�`��o["�q�t�����w�'�lj�m�N\���32�a�@[�S%Y<���Ѻ7�CP.Y.(f��N�[7�����.u�+RC�\={1���QЀ���N��V ���ʑA�-�B^#��]Y��	V��&��fdc3���� K������O��{��<�=閄���Z_��F��~
�� �8r@��z�?������ȱĘZؘ��n��|��=d�5����F��DLV�2('H����	��J��1F�m�Y�n�+��Q��j W�cl�t���ʺ<�w�b���[����&Ay�\�AlJQ{�pˆV�j���t�z��e{��2�H�3����S��
fz`Lޟ)�&��N�_Kb����S�j�$>Jn��<���]/��;I��w����ߩwu*�!�T�ޑ�bp�C�M�Ux�����9J�x�VB{��l�@�޴�1J���.�!�w�����㯢��c�&JwR�lC?��l[G�b6�.J,�z:�䈚3��>\H�wd�����ӏO'p����!�r��GG'E�wr�l�3�:6��}V��I����P�D�E��ҽ�7���UW[�~����[�Uvo���(vDg�Rj�88��C3;S�Nߧ/����$��KZ�I�!W5Iƌ�	��>aޡ�͈}�����.�w�%�ȷj^N|2�\���fg�׊gJT��	�1�*45V����^Inm������MTh���cL&6%ǋ�u���͝R.����N��G9`���+x��}6��4V#3��%��6)\�Fijn���8uM�f'��E�������Dy�66"E~�O,a��gG��)�7$�c�r'K]o�%g�
~�."O�~��n)���#i^�=�U���-����46���f[���Z`k<U|]Z����dUL�
=���d��#л����/k�x{�yx?Q�����ˁ5Q��ox�*#lZ�IylyD	�����z�C��8 �MM3K����&^(U�$'�Y���� ��V��נ\ѧ��9|�� � ��A�u�g�ӵ�,,J�����12n.��9���ٴ�B.y�@j1UJ'����A��%Ӳ��oRr�B
��������TF�j�W��1s�@��"bl�0'�s��Vl\�cvh(���cv6{�Z�\.� >;�31o�zD� ����!z�_�t���'2	�R�������/i�O�_s2�#$�U�V2��o�J�Zk?ew*/�Z0�_�q�[�l�Ecļ�DM׿%N�f8N���'������,؇Ъ ��L%�544����h��^2�|vl��{�є��`m|uU��J����2�����8ׅ��.5L��联���ј���Z���}������V�K���>m;+�>l6�'�)jSSL&h7j��Z�VNLS9�$+���� �Y����`E�����
?��Z��hw�VGN Z��G�'e���L�%���c�X�um��l�)á�ي5om�����v�U@�T���&���M>D*�3�ղJ�{BҐ����(L��.�賳0;�a��w�~�4 ��I�3K��ZӨ����E�~a�����J�v����W�\��r���~{�~�]�^b�0�I�7-�ױ��'��d&�R�R�4<������'�>�YekC�;��I7���.�N�t���h�p93BAj}!���j@2=z�ab�ޘ� V�z��G��Ep�c$`[\ �s�z��%:9=[k�Bh��!���:�#���X�Q�|���S�a����"*Fq7��,P���qQ��C������=jb1v>���Y-k��O�j��H)��F5�c?�u�O�X�h��?�����,m5����5�J��"D7�M���w�k�s������<K�r4VM�t=�|��zAaL�yC�����O�tΖ�/S}��g�Ѱt��qfRb��D�:����=v�	T��G1�غ`D�ӱ;����$��7��R{�a�x�`��Z�O�&���c>��	;D�
�2b���0?%#$]�h������!H�wft��� 8�P�}Ȋb�qJ)�Kx�8�s��}���������Rm�*��u�ӆ�t"�r�a��s��V>�oV49��NrX!��z�w.����<Xzf\�{�q*���J������G����,rAil9J֕s�&�G�G�I�<���-No���"6��W _;KW���m--N8���Ϫ���M:�'���F	� �Ǉ���f\��W�|aY��1�xec��#�BP�>��F���ٜ�����ݣ�/b�0�Gv�8���4^�4�0TQ�	�tYj��
��z2����u6VEP^��o��.2���Z-}��?��W������(�+�P/��S��V���̜5 ���ޤGt4�?��e�A��t�̵2!����i��&e�_\��Bʖp;�$ke]d�S�
	/���	i��U�q��6���J����� ��~a:�������_� n>�^vµR:3��l�i.��{� :5�t���=:mp��z����z����yVy�7#�r<��.����e��d>����~쥾��R�����N�+��m���(�F�ۦ����"�|)��G�KX
�;i��o%��V��OW���W:��īʙ�"�y'X�pa9�nXʔ�ރ�� N�[��������oQ��]w�g�U�~hY>Ye�Lr3��Z__�~�$�k#0���9!��?��#D�zol��皐��S���~VEe�e]`#�L�*���0V�V$e���P� ݠ�3��8O���+�J�n�l�e�	��ͮ�	�/:�0����u��w=G�ls�ᎂ?��¼�tu?�!81v L�����X�w;�������Ⱥk��z �!�p.���z�~=�C\��k����d85A�[u��Sh47_��5z49�n>k@���b�ol����~��Z7� Ff^�JK�#8��#�ո��Q��u�*R��L=�Ǩ�pQP�YZ�k2��z��5v�*��Ŭ��Ñ�ɩ=�;q���^ٱ!+ss#H��g����&A9���1@��=�
|� �}��w�#�lUT��*��f���D��e�@%�c���:�͘����5��뾻�����y��?G����������<5�rP	�)�\�#\el� (CX�+%��Z���Y������,�Jዜ?�A��o��H?&����C�]�*-SR�Nt��[�jA�r��F��/}Z�zMG5�-�B!�u��}n�s�5���T��oÐsjs \���XP^:Hz=��s�\56�Û~��w���W\���D�2���"�9��u������QZ���e&��_F���:�f7�B��Y���r�΋���VT��{���ۉQ��[�0��Onob�kVd��fhpȂe�1oo�ݠr<Q�� ��7���*�� ��$ &�G3��7�������0�<�@(a���a����w���A�|�c-n��n���ku�ד��a�g����_��{4)��R������jԢ�{~o��螄h�����H��f�!�Xc٫E~-�籄�ρ��4:6vݘ��̓�x
VQ��X� :�SZ���`��z�	U5�\3�A��]��$��Y�2K_7|ܪfq�08��\E��&��zws����}<��/����' &�)�ax�bt�s@�m�M��J�O��G�Jna�Մ+�+��\�<��A��b$)�eL��D�ڏ���]��(&�]\I	f����OF)>6�)).#�^�W4u�Fyyzei@�l'*��9aQ�D��%���O���A�r�>ym�gLB<�IX��՚�*��عcԇ��\ς
/Wl/=o�ѱ럡��u{���rc�M>����`e���T�;�������%���<�_��Y�`���F>�zI�F]fl�A�_K9�M'v#�^3��޶J9�I�"�1�f�����+�h��:F����ӗ��n�I*�c��z*0�̟뛙f��M�e�SO����$��ML�v���> �9��pf#`��;v{�Y���G*��O�_$�ϧnQ���L%!«�>t�Õ��".�B�k/f� 
��
L�������;�Zj.��ߠ����&�tbo�,�飋���KN��
#:wXjM��tEp�,ޟ����hLҗHzC� �c�3֢���#�D�f�]�-�	G3q8�%���q�����.ծ{��owA�qh9�b~�/�'K9v�	�r�PV�����Q���pt�.]�*0[ �!�c�E���=Ow��_^h��Q�t�7�XW�EВO*�(T�`dߥ�j4�L��G�����W1��T[�8�6O|vx_���	�1���o�%m�>�Ư����-�}��;v��u���n�U��J@ `�=B��%�E��ƞYr��c'��<[UP�ξ&>�q	b_�J|+H �k>�q��Y%�H���(â�,�i�9�.\�Q��M�w��ɽӡ�P����;�:��(�0��)��k�/ɨ�$L����+��{���`r[�P�%GK.�:	s�����c��O�!�X8�{��n��J�""Tw�������S~��2���gta��ԋ9�1�%��hMd��7YZ=1bn��|���юY0Ģ�@����P#�ҹ�ny�nI�I�F��(� �?���uW�H�S?ɼ�B�v����Xkކj���?�8`	���z�zu���<�zc2��4+8(��X\�Q����]��,r��`���x7n8l�`wo4S�IYv96�G@b�n����CXvrmiP�+F|������{=��,�o�W�D���|��W���L�P�7MYɯ��⚱S��A]F}oE�H;ww�I<��F�3\���|�nr�&1\���t�dKak�k�4;K�^�� ʉ9z}�mJa��2ܥR���Cb5��A���M3��K$�\'��'ڈ���0gn�xM�k�a�`/w�����Z(������PƄ�.�R���;&޳*�z�3�"�x�X9�	PB�UA�g��&���k�b�8����ᠭ2곁B7���$�>���`�q�B>R��ex�����'&���G^�גsm��/R�+`cO�9Kr��WV>�"���Tn�Gd!0��ģ�����a���yA�����^�ŷ8��mD�rzt���SН�`��Q�o�*)5���v�g۸�R������j5+K�1@���5��Qn�h�J�ߝ��O��@0��/o�,_�[/����Dh�̮�����Tu
|�2�V�js>~�&~,C��"����/M��
$��τ�x����b��-=i�Q�~~Ķ���m&��ة�۹J6��a3j#>����;ӌR��ծhq���$P�XE��;�tv�Q:b�;L�}�ۦ�ڡ <�ʬ��!�i@��w��\A�A��H-Oy:��� ����"c�D�aR�r�t�͝�n+V�x<"7Z�u���hW߽��YlK`Ħ=�O�F��HE޻3�ʹt�m�"����M��/t��~�L�[�s�$��@�+K)�5�:��2!�&����5�r��8����k�_���qM�����d���)������A��$�
�Y`}��Vd#e����
�aL�k�\G\b-�;�9�v��V��`�qat�ΆU���Bu��4�l|(3�>�vMة��݄k�/4�2�����u���yz�x�bpY�̪t5�n�ؑ����l���Qf����)��Г�����z�C�(�,?�0�l����f+��a�*Atl�"^�w���X�ĵsS����0�P�bKAcpq��_�f�L�%�֞�E�Ӏd�v�3em�aժ��b�� ��g~�io�<8�!Gs[X�A�׺[l��D�y���]}�T����GR��:ѧ�,�c�e�9LJ�_�eH�q�=0>[�b�����l���c�{0�,wi�`K/.���+ �e�S������d㌌���]Ril���� ;���RF`:*�En�ן�{����|���{�bE/����x���r/P�C
�;9���f̃���gنH���me�j��*l�����i�w!<��k	�)RD}��N6��~e1?<�U�Udq;�p'��7�䗳EVC�p� �E�Ʋ`6��B:%�X�_p(����v�ev6L����(�Έ�p���UEG!�UD�O����䧌҃�<f�W7m��ۈ߯p׻�%f��f�~��{<O!� 0��fd6��tDRWﶤhd.V��)�~��]i�2X��ܩkW��>w�`��	Xa�|�����V�'ܲM���H�j1(�v�`�,���f|
~�nyUV7q�`�4,�����Yɕ�$!�>�|���\��qW�:��_]�	�%�͡b<�/���^�n�,W{bo��j��>��S%'⮥]݂��j!�k�B�W=��&9� �@��ƻ����һ�$Ip�R2<+��n��<r�AZ�����V��+��)D�U6�����l����%v��V�`L��F3o�DK�#��8�36[�5���|�ݙ��Q\��@\��B���t�К�[�KýK�Q�
Ӝ�b}�J�����	�Z[��FZ��f'�>˂Q�ݟz�,��$g;�YV�wA`ĘiUG�c�M �e�Y`7��[LP��5d{��yxBR#��6�M$m7�~lϫ��mfk�Clb#��D}K ,"���M�)~�k!�������P��q� ��|�#9Z�d�.��Y�6��trA*�m�U�CE7G����S��,L�IE?΢�ӳ����B8!�4��~Wof���eDJ��WS�:���3bi��b��(�g_�u���(�#-�����/dG���c"� 4+�$�Z���Wyk�{�Y#�ߖ�1&S�����~�*��lJY6��`�{K	�����5�<�X�]|��s1<��e4�d,<Z��>��Lx̓����U2H�X�H�� ���'���������#$��P�1(���"�L�v�p$qV�_&�����Fz=-�cY0��eUdD�#S(54F�#��X���4ܞ�H�ds�ZjD��D7Z!�
�L�@��+MN.�sE�igF�wU�0��Kax���~���.=�l��&~���j�����e���\��x���Kkkr���
67I�;�����+xTf�n��Fo��=
)3���=��Ej���Yٸʰj���Y3�-WP<VZP�lcE�)k�қ���,9g)��\��34�ũ�_.�:-\�����w������/���^����_������˵LF�R�贝c�gߦ��;G�:f?�� J?�B����'��@�-"���6_\ �h���h&ܙ=�<�eY��C��_&Fd�_t�%�X0�MQX��a�
����cM��m�p3�z�3�\�-z�QWk�}�<�@1��.��7���E[�H_����s�\�o�(b�Ңt��@��q��&ǹ� #3�<�
_�hQ߸�a���+�Z/����?�/[Z>�\�1�?
m�u�t�UI�u@,yϿ�{���z'Dj$2]������?��III1W�/�H���K_9�3��$`���-R���9�TD�ctZ�z[��1�J ���x#!Գ��U�bٝn�����e2a��:��,S�%6�/���.��g!���r�{�F�9��sQ��)�.��]^J���2���� �(�hވ��
lS�T$�IrD`Q��,пB�:���H���Z%*������~�8��G�给��=c��l7f���ۭ���SvwZ��y��k�'��.�s�o��\9�P��B��26U�+ZB�V6X�R��'�a��ex��wdid^3ñݪ}��]w����_����w�ޏ����y��{m��]���-�Y�]��9'���A���"��U�^n�Z�p��Ά�=|l��l�=�@�أ�5&&��7>g��ܓ���}��8+WC�X#��4���s?�\�f��)��M�kԹ�8q�f�Ŭ�Y���p)F�	t�?
覽��C�ӌ'e>��|�u���5�h�7ޛ��]$��F~�z�iqJ�F��=��?n�6���A`�dlos�evQ+	/C�S��?����.|���Cܯ��8��7|Y�F�=AS�澗}�6��k���_{��e�[z�F015�6��X-$¥X�������aR�:���lg4��WCIaM�<`t�XGsB�+�?��<��>���M�Uu�$YT&���ca��+����0d|m?���y�X���5j�y�Ҩ�@d�\�S\���U�C�,1�P���E��z\�5��&-}�"m���"�Q�J��jj��n�/���ښBHXI̽��&D�2^����]��#�[�h2V��]E�c�T�O0�'�c�<Y���s#�Ƣ�뾮m�F���^���c��~rk&�z��������;tf3�DnR�Ca����o�EGf����G�B�]mLTk�WAD���5�5^E�D�_��u#y�G����n�dS<�%d���s#j;���5��%��wĩ�m8�FeLވ{��y�����GGY���ԮѬ��f���p�g����!�u|N������S��ܶrx��R�ɴ��&��K��>����@Q!�;q:B���k4.�]u�qU�8��;d����� �UQQ�u$V₹8�~M&�MVvv������x�<��o�6�lKS	���NSl��A|t>�a*l��57 �`���L����Xb^�q�J�����[��>�KE���ӟ3I��bC8�b�d�*P-�>Z�f]T�C���b'�Eq�܀^�9L�A�>ʾ��8
���Ԃ1��4fnC�
�W��'��׿V��R����N�P���(� �¼թ���LYq�V
$]�������FÇ���ћ�d�\>���~ZI����j]�1�(�z���d;ߑr�3$��P���/1���!����������9^�x�ˌ��0Qڼ��_7�̀,Uz%�i��Bj)f�v�p����K�q=�w�G'�c+�]6+�'�kmA���^Ln���K:�fS�PZ��?�n�3�C-��c �����E�M�(��"��P�\���HS12����߷�oYd�Y�X�~�8*wW��#:��ꊿK���!sjﻷ�{ଆ26 �Q���8�`tޖ +�8����D[H�����&��e$����l�!���,��y�%c����v���0t����P��x�aG�u��V�\`�Rp�5�dD@xZ�S�_77w����E*�nf��<U_�g���������7X'ׅ�J�\��u� �����̔�J�U�,}__�"��+����YT�H'8��y�nsh럄hhξ����.������OJ�f��3.����̷�p�G=ת/�J+vQ8�������e������7��Cñ�i�&�]m��M�G�5�����>��:��<SU{��5�n}=�R���#rr���1w��� 3�S��?:��$��5N�>.+��]��0I���OI4� ��6:�+Rjhh�/x�?�����De�II	y����?��A���#ef_��U�縖_�k��Ĉ���3��W�T[���4�W�p����SI ����r�y=���H�E�G2:|��Z&��9���i��
L^RP��8�,C�9 `��?��:�����@���mt�/	b
-�Jb6��=|�ǶGٷ���>xQ�&�,ȑ�D��� 6��j�R���~܄�bՉl�1���n�K����z:�>j�c�\j���KZ�N�fxI�Pm����E)N��8��޺���F���P���k��}D��z}8؎_܆����3��h��5���PBAj � �R�S�ތ��3��K�-[L�����Y4�4�'�A��3]�b�qw�f��>DIZ�9?*^�ya���@�춖"(��MK����ԢwDEG]7m)�����L�~�Zس���X �B��>�2�s�γ_�=]��F��?�:����@����ZǕƔ�*�ެ.^����/��.9��'j�?{��ц\
;�ej��k鋾k���,$gG�b�ޭ��{��������E�����lb���d�TLx�������pTH�a���"�,��Z�(� E9 CEhl K��Ô�mw��Ao���3hG�g�98;�u�R�0�M�ˎiH�ɓ�D��K�5�����V��Ǎ6�����^ls���jM�	~*1��5��t�:��T�Ra@V�u���*�k�o���D��\�;��X�f��֜ɾ_��P��>u*Iŋ}����WU�X��J�)��;��{��H��楸���e�0$r��|�ܼ��8��G����?�L�� ��x�n=諞�ί>�yP�w�	v�\�ӟ�@���oo.�?����(.~z�/K��0w7����ڪ����h�yH���p+�(͘#w����Y0G4`�P	���[B�h~~9�
L,��$��E$; �xJ3�l���졆������)��sU����Sv�:��P�=��]�J`��J]<Y�*z����^�������}��l����*���a������pl�2x�3���r����\�ׄ�e�D�i
Q�t��-Ԟ�>�L�2U��[]]h ލ���.[�|p*��� �H�Nr�,���u�`�#M�	aMv�|�<��S
HS��`��!n�p��T��1x�x"O�<��F�;���m>_m���;���L:]���-Q��̊[�S-B5e�����K�l�������2��/������|�`�mSh7�.�q�P�x��&�X���P���n�q�ߴ�^H�!���=s��.�� k+k�Ì�}��:vd���M�s`À �]H�s�|�+��BJ�<�#���h.hC%�����\ӏ>G�ev������:^��f�6�FڿE�o@����=��>�fJb����F�I�8L��z�1 ��ǩ�`��4|�u[J(\� =�T�Ũ���b�+�k�Q��]�9Gcp�G�e�TmRV�"�M	��d����{�o���ǈ������q@���jj+�LpA5�@m�:!���'�3��(t��/�OC��/�/�:� J�*V�km��+I�����e4�/����?��l7��A��-`-�z�����L���ڌ���vk^��e͛.v�&5�`�-k����K�x�ĉ�W�ۺ
�����(��%H=�m�񸸅�&@�f�f�dl�L�!�`	MF#c�QA�� �+lu�L�Xkݟu$A�li��'�V�;���Q��B0��0[ՉQg��^�&D���,)���f��|�[�|�����y������F�����s�1U�bMgĠ�p�#6�����{C�*faN<����g�p7���,;�E�ƿy&� �8�Xp(�z�7ܓ��7�v䫕��*�ˆ�zX��a���yZ�HE�d�z8�㯿P�q�������C����A�2�r�ʯ�V�mA��� ��q��%8�q}K�snX`J`O�nb�F�4�׷��o�B�g�},���/&�Ē����j�k�s�"8�e�;AV��X9w�j�]+y�|:	ޤ�:P~,nhS���.]sv��Jwc����ï�IXjY.N�9�U��T��
͛𶑬ht�*M6|��ӈ���	�|y�V��:��<�5�3���N��)9i~�J�މ�KO�8�|�&ǩS�&=�O�(Ě�@�O1�O,�3����&��̮�E s��u�X��|3r?;����HA������|�Qu���VVƨ���2htL��������~��:(SG�n�a�W/����mL??
�S^���Z�k�J�F����Z��}\��s�p�p%��)�rú �Ȁ�;[�^g����#a�r�����:�N�)؁�������� �qa~�
د�o�M�Jq�z�t>\)Zz�h�es�O�&(/�'��ĒG�~8� ,�j(`$��G8�;����s[�U%|q]�s�܀���:���	��DM+��� 3�0�b�Su�kf��?�q�9��AӖ��g��%���x����B���u�@�x���Ϝ���R��9�O!��gW��?.� �˛<!pvjb��|K �,1y�#�Y>�ǵα$��@���,Ԃ�Q����쾴�e���>g�n�%0}�.���G���fW���`T���%0���<hICR+�#���|�}3%G5�x�1��Xu�2�t�p{�R�2��H����b�fwx����"/]�Eȷ���	���'��	�! �b/`���6�s�?�������9HH���`i�p�9N��vqw�䯽�E�*`���!�F��	l���_Aq��èY�Ѡ��oX�3nH��_�������z�ec��doG�es|sI����pE�K�=��'����IR$�
�C���\h	ȷ5mmi���D�"�ӿf���=�=8�\Bu������r��z��̌%s�4����g�����KQVl�U5�Q�8&��<9]��K� �W+ �|�u)8	8TKZv%�����^����c��o��ڸ��zO�U�h�ȦTISGk�.�h;��Y�< ��.@.� �p��d秷W8��ơ�#1+����qRek*�a�Ms�N2���n�<N��j]���u�ҢK�Һ;�%D��]����[�)C-ړ�#>t5�!橌�>☜V�v~��5���  @߿�o���������u�ӆ�0���*��R�L'�]ʋT�� ����I��ˋ<Y�@�t8&��3 r	���L,��!ǲ>�w0�t@��-</L)Q5�
w0�mq	����[̬�=d�@_�����M��fx2�Bk��Y�����7���a�;���|���<�����.�~,e� ����;��[nN�,Y��Of�'�U<i?�>�h�v������g�^�ް���H�'�����Z>�(F%�L�u�M'�`Rr�J~~�$ 3�!wD�OH��������_�F������b��@@N��� TG��)y��msn�ϸÀ_l����L ܓ�N@*��p> � ���>y����*�yw�1�������4�X-a�}aU����?�e`Q��|�ѣ����'#hV8  � �4�	ﯲ$�@{���cU:؍R�~�f0X��W*%�F������U�|�tHB简��+?%HP��6���Ngfg�(<iGai<�i�J3�sN���4�U�&+�An�0��Q)�s�a��;���>&B��f@$���*~���1���&�2_z�%^6�aR�u�+1(E�b� �Ţ������h7O.>ѐG���yy�B"g��Ǐ�@���>�����o�i�.r��Ł�e�<�x����j����V��}�xi��/E{5X��},u�`�Td�j~�J��:{��挌�R�$ŉ<7n\7ļ�VyI )�"��m����-��~�t��c��m�!����q}6p�M���w� &��Gm����>	X���٭� �30Y���S��OwD���#�ϰm!��L91�v���7Ԑ���T�}��m�� ������y
�'�&���6�t��k���叩�ɂ V�D�4s�V�`Y>���9-���+�E�Vo49�
����a�y�=xp��{ �@lᙇT�X��s&��mJϦr�ҿ��@�ٹ�U�t5mn@ۋ}��@ƍ�����M�H�*l����e�s\Q��^c��o�^^������<@V��[8�C/�aH��ǘ��sz`�4>�sq�eNe�E!� ��,*�N
8Թ�l��.Ƚ�Ӎ" �F���"�.�2�3�+�엥�Ŕ��&;(8p��TZ*qK�4 M9�]M?4�F�g���
R~��(i%xRF�$Y7��������WjSC|����?�Z�;vqd:g�V``�����gtox��f�0xo��6���8�^	�=�,.������6bp8i��$�0����z�'3�����	�LX�Je���kȀ���]e �<#����}�N�333��-�1�T��sE;�#o�|�z0Xr��D1�`Vq^��[�������a.����8�ъ��}s���y�
�3<?��5n���-u,r�&gvX�msI���g̒��o���v���V����j}�o����جg����[�M*�?�/����0�{`��yiv��];B��9;�B��4 A���:�Ix��U�b\[5h�9 1���� Ã�	�����t���T2�퍣���*�o���±M�9´��&�g��� �?P�@����>��a��Y"�v�J���Nm ����y������@-M�D�+-��/;/"a�� �͘
tm� �_�K��r�+��K����s3���e検K��]čb���_ds��y�n�xvEaa�7M^���o���T���|��`��]3��%�P���?��+U~�!�������02,.-��m�YG<�3 �tV����J۰N1h���-��Y��Xָ���G߭��l�3!�VL�617A~�|�R����Z��w��L�.��I�	��8���d!�m��eH�ifw�^�*Ui͸B'+`��117P�k|BV�[?�ѣn;�:�K �����s�	�M�7q�'���tZ�������W�R[�s{���?\��	8�%�nS��vW��5~FfW8�"`b9B�\p�Hn^��͟Ѻ�l}p�v�4���^G�G��_�W�طo?��е��V��N�9�B��5���={�1������ ��rb+�fO,�>:R=����@�0X� ��p�[wۙ���^֝�w��&WDZ���O;�Gq7&����1�8�3��."�������W�ϊ�H�G�������ҽH{3�_3ိQw�܃*�7d�i�����3�<e�3���&:j���~�9:�O��9w� ���@o��9�^?B:�,�<	�/��Sr�G<�t��$d.ܞ�yꘉ@~
mD+��={� �1��=M>�á�$!ã�T5��CU��zeZ���3��������RT�DY�z�!��$�_������:��\?��LA�7w��cw��Თ��������_3 �5r���I<�r�B�!ؕ���Þ�=���)�Ca�j�Q VԊ���c�j���Vor�t����M0eڬ��������)�6ˠ��䭔�R��Ҧehb��蝏97����3-�g�ɫ�`�R���J���J���׺��ij��d!��1��0H��p�|�&��߬ɴ�m�g��7x)�ۜ$�|�D�f�Q����y3�3�{Gȗ2������2�i5˸aL�89WM�Ƃ$�Yp���NL����_�d�+T���w���W �	}��uJ ���5����<'CsΆo���M�,.//1X�s�a㈰�?5=a%�ܰ�c`.``�6�%I0�H�<�L�l;4�����l��@}�C�ј�����+�����bY���'�'M�C�/s셅%�$��M~�w^��G@��,�Ѯ6W:�2����(e}�|��?�ø q;��"��s���\��;;�)o��`�p���8�>k�UueَY�U�u�L��Hۘ�H���4�;����B��c���1u5ЎV��T��,	(�G@�bM�gfo�$�)Q` 0�����O�O>fV6f/V�q0��|�-}��W6�sh�n�0�m�$A� �ǡ!@y��.^!��R͇[7oaM-��pQ db�	���U�M<�ӧO��s��bl޴��였\�i�����T�<tAk��֭۹��z}ʹ}7_h�7�:i衢�5���� >rz!w��C8���"c��0]b�l���"~x=Y��Gy� ���$�2��a�)B�Vz��]ݴ�����~?�ɳ^l,-���0=���A}`i{�R��@�}�'ޡ����]'������E.)h���C1��oP
��!) 6�W���-���؋W��8��)�(3^�0ً5 ��µ<"�Ѫ��l���tw ��<$r����ߘ[o)bXz��}��87��M̦a��2vS?/#��[ ���b_�v���&�ݯ>0v��_�vPK倕�{i�f����F�T�gpu���|�7g@no�C��6晿G�2��{�i����ND�ؾ�����iF6��6��������L
��n�jxq��=*��§N�<t��(9�.U%�.-��s�+HǏ q������0q�4]�(���$��5�M�5e��#����$_�h+�{��:0�>��ٜ�E	�]�9��J�������������r�*���u��SϓSmV$Ŧ�"�ƧUn�� �$i���&�o�qrNQT�l>Q�]ۼ��T�����s�ުc����:k
��y������'|sE̓�.���\Y��Z�,�������l)�% 5�eM9�؊]�W�P�*p4դBX�1�R����m)����,G���(u�< ^��	XM��T�v����b��պ�S���K�\7o�dS�(�����$���X�^]]a��y���儁3�'���g���Y��������F$�Ċ����N�;/�B�%�LrU��^fܱ_<Ϙwiܲ���3Ą����4|���
vÇs����l��u��o�jh&�4oٺ��\l�7��gΝ��>���f`E)<$@�
`��.���9��*�zJ���r0�!@�t6��D#B{��>p� ɡ]�0w�ޡ'N�ytL���u�#'���.������|@�7|>4���n��7EL0�<؉\X�� O��S�ԉ^7��\��H���6A�W�LK�4�~ ↡�lK�2M�gq@ a��M�|N8wW3���=fw���W��W�$c�<Y͎��6�3?�����^4�#�����Ak���>@�z�)eo�x�[�o�MyH�RM��M���  }��Zs!�l�^���Yf	ߵ�֨�c�x>�FS[���J@���(X6ڏ�'��g�/��Q�VSV�l;�
�XGV�Q�ބ}���"U�ܯ%�2nb��+OId�X߮Q�5�z)C"�N8��%)�8D��,�5}��Ռy*�7rK�8��;6W��=����-+�m�Я �\�)_��"r����"�����h$|�R �P⓽m�92 uG��,`um��p�
�(����7{�p *��N�8�ipl�}����������ms���9-:'q����4�D�;�Η�^�����x��YS���LϲZ �FU���s�{;�%�t��L�`�|��c��LxP�v~7ݽT�(���|)������%�m�?�X�Jg/"��X0��:y�Z*YyG.q�������[GP�P��W;����7R�4����\o�p%I�e�c�t�;]Y�#c)K��*�SQZ��X��������w�f����IP�+¸f�m� �Զ!d��j!d��8{A���.�	�+ d��zc^ie9���T]Ye@�ekk�e�\Ԫdm��Pc����k+�TrB��� H��	gβ��8�[�
�
)SAR�m���`�q�_�V�Mgk�ʠ
�`<�c����A��1�8s���av�pu��2�l�кc;+ب��'D\,�@�6/Z�������o8�0�W`�nۺ���B�� �����y�!��i;So�`v���èP,�N��e�몫��>����K����{�FF�1f6��H$N�6��~ӛ7o2�����l���`���X� X�ŏ���.�ގP����~`�M�S�.`尢�! �Cp|l#���á�w�~pCE:h��lN;xc ��G��2�i4]1�x���[��Ģ�l�x���p#h���H���%yr�	��M�����ȁ\)��<^��)��n��������0�B� �3�(ց�y�-e�U.��,˿�uaϤ��#^v�eU��++��h�㍇p�2)`� �z�3˶�9�,�c�}).7�,v����v�)�6u�^���/��:\���F�+�qjT�������VAȘ�s7d�Ɏ�I�����D��e�n��nP�|%Z^)���v& ��y��7P=7�/Yy�����ߑ3V�=���n{��=\�(l6�sJ�X*3�l�����<L=hoX0�׻> óvݧ�����F�+��)%��I�ae�uN8��%7:�p^e��%6��a��V$z����N�� ��*]����A��u� �s[G���i^�n7o�6����"楧�;�~�� �N���4����7�1jj����dP�ϱM�o7d{]K��fQ����OTEi�;p�������L�qT �\�i�4f��LSO���68�M�x�,�[�.�*��H��ܢ�2Q����s`�C
y�jl16����b��lf���cP�8�^?��X���},/-���;~�R����.��x��p�T��0!�g*�;53Ś�9��@���v��Օ�`N�B� C��Y�3Q��,L=&Uv%���2�2���T��$��s����;X��.�d�8�z�
���:��	@�N#��ӓS<���8ax.�S��3`&�srj¥���ffP1q����qJ�8����t�@��a��p��pG�������x�(��5>g.�l ��_�<��L ����%�YD'A�zd�{vS����o���^���p 2��R�m�~�]5NM¿�Y4�g�l��I.=a����X�6�R��"��R�+��Я��q́�[��b���n��/����5�|����5����VW�`�z����e ���č5�m�>0�����Q��;܀�Fd@u��������
^x��Yg�n@8��,� ?�]p��L+ѐ=S�� �ݢ�O�A@y���Ct׾]ʎ��2���c'�ft(��a��ɬ(f�u�cYȲG�����)`��`���-H}����ɀ������q�4�s��m�3���t6��m��{��ۦQ8L��g߄m�쒦�%��M`�3��-*=��ʏ�/H�������I�+���(;��o17��S8)ھ���p��ZA�^;�?�X��c�/���������~�`�̯bEt�|o@��y��/��=�ڸ�@~��yƳM��w�=���-)�X����:�ύ=��f�k3�#	X���Y��uF�{��T.����-Y�*�
��<�����+͐؊`i #Ӿ�sB�^HM���_�Mδ�Mj�4�f���z=��s��>��v^��)� ����� tU �+|.��%aBa����K�N��؍�\�p� _Xvax�
5~� V?��īt6��C����k�n�`�Tr8B�yB�(�M,�&�}�.2 �MD��)��H�4^fq�={wӶ�[�ُqF6�~�J:�<�2�n!δW��n��M뷕g: ~��:����
��b�G�)=]Ơ�ᆟ{/9���!�7�X�e	��*��7���4zuUD�auQ"X�tXY U�4TP�H`F�<�`���iN-]d����HC�l.���*T��`�,]_q�1X�0=�K���"9�pD�%h&�Dzvr&��(����t�,Yܭ��Ç��ŤR	����,?��VN�X�E��;v�$���1��&|�f� �r�-�w�$��n�Z-�<����>d"�d��ʌj��w,ٔ$+_(X�ʬJ}��Z�VR �h�e+a1T�.�f48/��4lRpͿ�7�8��J"����.1��L�bM��K�#�%��A�C�T�Z&�sQ��U����z��0�~�׏��v$w��=3�K)t� #�$��~�R��qLP�z���^x|wLB+�
������3s��#us�?t�5S��>&�离������!L]����9��<�FȞΓ��V �ٞ�ﱤͱ�����j��O�6`7p�X"T�����l`����+�@�ha�i�#;>�G�C^�]ّd����>�˛�@�T*h	u�%y����s���M����5^A٭V�H��� �ū�7	��:��+Y������b����Y33�,��U���gD�e���$u}Ѻ�ǐ�Թ�V��X�|	���@����,�l�0���?��e��F���kr폂�+m�����S6�@�`��=
��*�D���Q9���L�N�΀_��,�kp0_�1���gYPd@X��	��6�0�T3�4k���<=W�u`�+��q�E0<�ޢ�/���P��@uU]��+�ޔ��veT���q�(�e`v��� �	S���(d�B �d���xځ��m۶�q@P��@9Tj�}7�.8^�H�=�:���Z�l��2&VBd��]�t�:�c\
�ϐ��3d����u9z�ĹsQ��N�����:(~�E���@�{�����d�ƫ\ccm�J�H�߻������..2�h=L�1m/�����KJ|+�n�QeK���]� ��Q��r���54�ۃ��$���zt�1�7&�7G <'������
�}d�@�.� ����K����4�鸬dwN�oe��P.n��W8'� #
Εo$��ª��>�Z=d�SI�����+ӫ����:>5��d`�<��D�գ�uKP����a����Yڎ��X�]e��f�hJ���#����Ӝb�Ԓ�R�|�.��3������f"�`���<`�,c�qa�@;'v�1+8�̑���ɱi���U�)�Ѓe�$�i'��0�¢�W���c����Gp�[n�[50&��i��^�ԵO��-s;�x�m&�P?3�µ)��<�����2��q��c����I"� u��d���gN%<��o�3�$�o&���X=4H�f(1Ry��B��q!��"Rw=���n�ڭi�L;�Z�0i�}#a���I#��?~�%-} �$�Mʹi�����u�jF��Ed��d�c���Q���ʁg(	G���X5�l�%GH���0�Z�m���S���pT4%h��Q��쵦�4�u�p��\Z��`X'���k��Ղs4�EOh�]�4`7M�#Ji����@�h@���P��� ^�
Nc
`��ͫb���Z���H������^]W"�p�x�V�P	ncYΥ!����tDN�W��J��ΰQf0�ΏM�'Ld�j�A$!� ��^��	���R��_ل3W�l<Y!�����ӷ�<��4��+� �HŊ~���SS|� � �X����:����	�~N���b�8�a�8y��y!�	�"�o�VNӂ�;��x��B��W,[���w�*J�S�	U�����y��p$}P���T&f�(t��φ{z& ��DyAB�mÉ/�e$^\�4H��f��u�4eR/.I�eLt��1o[��X�?7/9d٣�����nJ�k��}ew�+������,��Z�����R
��Z�藗��f#`R��MQ�)��y�m����M2{�k老36�j��L�����ه��t��BP�@+����ү�bg��9,��%��T�������f�#�	��R�^$���t�A?h>Q��a����b�����������7?�%�p�����؊�����v�*�ӭ����c+;%��D� �EҺlY	B�?jg��q�\�6K7?���Y�f�~��K���2��.���EJ���f��~<;��Dd�S�qJ��Ʒ/٠W��ɺ�'�ڷ~��w������@,9�G��z΃�ȝ�sg2��&�es��s�7�hM^mw9�������B.`S�n��d�F��Ыp�#H#d�HL� H���F��FК�f�_Az�cg\jy?���V�ϩϐ�ހ'!O��=� Y����u�J�f�E��˕�U%��{j*�$��	}>)��פ���֑� 5q6ju+)4�j4��ܳ�"0^�?^j�<��E���b�&{|���Sed���+6�@��D;����k�wf�+?��4�l�2�h�2!�� ``86:&+�\A�8H�*�1h3V�E$�S� �.�t��`"@6Z�y\�9��h�qE�`� �c{��^=����\͵�i���&��Z��7���`���5��o�K��$͂ϓ�}���X��J\�:$�����;�dz���s�IA0��n���S��M����%�VV�5n=���āw�J�y�YYL �!C山Q�m�A\K*�Ol< ��o��! /D�0�xcmOt];`��?z�����>�=g$@;��
�K���h3��Ă���Z`�dm�"��}i��O[�̴��|� �~к�S@�~��t;�� Q9૷r��o��v�z.2!�����Z����hv��){L����[�8�0�r=s� ����M��� �����MF˕�>��=l�ƭ��v[e7��y�9�aK�0e��T� �A)�ZE	?��pj��N}[#�,� �9�O�U��Ϟ����B����������\ �}n��&�;�#�)��rضX7�'�{�}��ФP�.;P�z'Ձ���6J5gs�L����тi7�V���G��Sh�T���6�mw�i���6V� �<5�PGP.w��s��  ������ט?n֒�m��S���fbu����-~�"IwiqM��P�L����3DX�`;<됂�d�|�qG�2���@c�I�>*����ȂJ��5Ţ��`g� -��`�=WMK��%�c{��d�-��3+�$u~�sX�h�h.m�1�5҈(��L6�)��"�I&�Dj
��~CU�ozj���h�J�����=�rG�n�\��h5��K����,�,RȜ4;;Ǹ'�����~���K����b����M�s�����L�}������H��� r]aE��\pn�U қ7qjV��cyL�dcd4�y�ll���A�� hGvB�A���iˤ�ͬ\����n���1�B���n��mZ N�
N�~���@j�Çq|�]�c�)�07m6���V"�]X�3��YI��E"�����Y]�7ծlټ���N��� V�$���%�0��Ks4.�
j|1Z�Qu�t% �|>�m�n��ox�����K%w֐�h�P�Α,kagC�<��޳������8��m��2�~�.��Tf��P�F�ئ�j�'-�������7:��T�_Y�KZ�W� �f5[��vO�������f�����9��$M�EZ�2qXE9?/�7��F����@���Y;43�Z�!���F
P��P�H�y���e���:d��u�u�S���{���n���t�(emߓ���w�8��ip��b��������:�x���Ď����������y�!�^��m�a��qHW�6b��>({n`6� V�7x�4;���j�0�>�?{�k����G=�����'[�J��z�Q]�9N���Ӳ������t���E��J%���޴K����ȥ6
;H�I\@pgK�H��Zzz�~��|�ק�hΌz����%����\ �ľW�P[f�2~���{d%��{g�;�U�BUfd����5�k�q���ZBy�_
দ�H�׃Ui\��Ό-(9S����	�Y4i�z�w�������!k� �_�ڈ\��Q1#t}H���8����>-`&r]C����hbG9�в��{�c��k2��!`�����q@*��$��>����< =v�e�B"� �ϟ9C������EZ՟��;��N�Uس�Q��s ���J�0����(U,lۥ�__}�U��[o�Ç��T�pL�oG��7DG�_���^�0C��� ��.k���κ"����h�b�f�4���f��=�$w�R"�c�#����`�c�I��س���̨�R������1
������J�=�|ǣNc�1���SO>��H*Z b�z�Pɇ�.��2����?ގp�>��"ՀI�Ϡ 5E�c/m� 6Z��$�L�dS�~�#�|��7�.�M,l�Z�M��F�xЮI�M|u8g�
��[ƯKO�:O I�7��T��HA������YP��.�9i��Ӗ�������.-�(s�ʚ�uI��I2�\�`N�� 7�l��Ǡ��L�ע����a��,=}<��G� i�"�Iu�/6=����1$ 9ܻ!�I w�HΕ��*b�Tu�����b�4�Ȁ���I�O���pG���G��#!�b�L�?���Q/d�Hk!��v3q��&�?ي~�}����m)��w�|(8����	G��i{����QN�9+z�P�YJ]�T�5�QXͫ���7]�H�AVL"hR|ըҊ��%v�u ���lM�4�%\3���u�oIgM�+�N4�+-R��ue�o`�d���z Gtڃ�t�_��GI�
Ԭ����v
 �ߗq�$z���5�8I���V;�d�#�΅��Z��k��t���@.��x]K���	�I��	��`��?��㘽�����������IC3'8!P�=���z���Ə�&�.x��*c>�_���x5��o~���o��;I�.lc0
�������0T�Y���B��rc_��w4xd��&$ �q3�U���uO�{Fit��A�ײ�����8ڻ6o=yF
�mm�u��Ele��͵�5hk���&3��Ҥ�1��5;D�>;ya2 ��1��{8Q6D&@	�����0�-`B�:�']L�R67hE��0����O0��4�����7P�Q"�C���	������y��iGNI=w��h:�@*}�汏E¶:�[���)���MçM����㕅��_��, �j��M�c��.K:��s�E�:�#sKa�<�v���K�my.0�McEb�1�y�F���G�;�w��[ë�ka� �d,z� ��g�G��I]x� �e,8g6�Τ��Yer yN��� e�f�	Z �#k���TS	'�1��N��*����m��dp�Z��Y��.8	ح#H��(g1�˥�wl�g��M^)��t[���N��G���˪ͱ�m��)݆w��.��v9:��I�Q�:�ӣ�@1o?��@���i:z �g���6��al�<g(�eY�~��q�}pQ�!J]g�#�tT*=_�$��AS���1r��� ݐf�du-ł��M3t.�aJ���\1`l�P�_j',iz0b���'��y!�py��Q�f h5��ԆJ=��{@
�&]>�t��i�2ٜ�Q�g(]�@1A]��_ X3�h�99����E:���MFP$$e��h} ��4+XZ$��J2l���C�'���dG�%OT���.��3Ϟf�ٵ�׈{nܸ�Ȯ}&���>�,� ��@Q �8����^&F�6��=����;���{���ڸLd	V��'�9X[
]a�n���>��*W�j :.��
q�t)�3f�-f�s�n�y#��cP8 `�x��l#�B#.D�s�W��p-���͂����:�2���v����G�]>@��=�i�` ��/��x@J�����@�~aa�m_���f����c01� u_�𥛝C��Y��,�VV䌠��?��4.�@hw�t�$mV����
-�ܱý��k�S��1`ES�O?��}���� U��o�+W/���~�?�>#�x�ݻwf���#��ڍ�����{�v���&���+���֦f nme'3���F�C4v���'&o�[�e��h�c����9�[�&Τ��Q�	ط�9���g^���_�R�7��p�
xҳ���F�f��qD�Yի:��"�L*N�$ �:���\TI���5)3�ts�n�h$j��������51�H\���"�� �f|�s��K1�����$��)�Ϊ�\@�6�h��ht�q��)��1��>��߄��S���Ta`�6* 6i\�i�r�I�guc���^~H~�����6��n���2��9�R��u���4D��*s2F�m-6u��9�k�|�L���LAt\XsVt'�M����a��.�KAIRx�ea>7Av�j9��U�Ke�{�X�D�z#�,s�-��������CQ�ÎFu�9O�脈]�����x��)��sk`����I �㛑�)kUi6c�C�G%[�?��4=�Z(f�q&٠�^�a#5����-ж֮�Z���h���kqi�èmZ[�����E,��Q�UOӅ�9;�_����=l���X{k+�8��1@��}�R�	g�u&���8�P�.�iak�zS��è�\���s�w��^y}�5��"�����N����
�e��/ؿ^����`$�=��h3@�Pm`V����07�ynx�cc�,�i�D���NN�y�b�bt��u%� ����m�]�� �xޙ6���v7.���f��� ��|��������N���0����<8�(X3�t�Df�2�(���n޺Ɉ�i�/��*����
#�G�A4�:�A�\��, ��{�5`n���ص��ڳ�-��gQ]��3>����#4�S����D�*%�����F�(�����e�fU?Bݗ_|�=�/�{l��&X�"���YPH;��3����h�:��T�^o���g9~dI|y�"��0IDuA&��܌�O��_~��9V90*���h�����C���4���*C�����d��/��1QM�ܘ��G�o�ar��B1���GI	mI�I��.���ԩ�(򸈱7�F$��5���2#� `��1.&����q6ULx�4��䨇k���ـ���Hh�v4?��W���=��٣�n�q	���I���ͻ��WWRUM1y���ϤR�a=�s5�v0��D�]�"���f��E��CdͰ4��l���6*�ޑ,�uTӈ�kB�K��g�3*��J�'vBʃ>vL��5���)�M����D���_+X� �V�ћ�;�����c�z�k�b��f���$V]�6+��啢�t���1Ɔc݁9��L�V��*VR;�c��e��ڙ�e��NGn�P.r\]�Qv)�#|p��%w��m8r��1i��FA��e��΅Tu�����M:=N�t�.m������<����Sl�o�%�I����Ȩ�P�ET� 0���V?����G]C�����lZ�K)H ���\_[w�G�hga�g��'̲q=M�ʶD4TX�/��T���s���i��ٳ����S
0{��S�H���
��/PS��ӗ�OE2�� )ȧ�IZc�.U/*\{VV������DaA�l����,S�"��|ڕ�?!�M_�+���	$HIC�R�)q�D������e��h�d��̜q73=w"L���8�75�e8����$����i�G[ec�a��>`c�X�4��曍�m �T ����0_�Gǔ��7������B��s�X ����/L����-[	��e`���>�W�i��}�U����"ʪ��z�� �ӟ8���>�ܳ�/�X`�X��c/���������T�)���08��3�W�y1�P�L%��Y!,�m=�\��
P�K���=].
�S�s��c<"����Fvǿ*����l��Ȫ�.X ��S�S��{��g轁'�+�l���0��D� ^��4����!˂ă�D���S9/x��f%"��>��Y����A#�	��8���s�`�p��'O2������ �i�yP����H4R
׮^u�KK��t�U���ڢt6F&�l��I�Gqz�7�$��?�0� ��v�'=���4����:���縱�������>����Q�Ʋ�F��:!�4��z�)v��E��Ruhi�V�6��3N�Des��Q�y�'������I�+�I3�B����"�|'�C�)�"�F�2�*�!|�C��Z$+�tД��i�=E,]���Q��D���vǰ!�^�+��K�XB���J{ٯ��Q]x���BI���5��
$
�E�@�a�T��|�Tl[ӜQ��n�]�d��x�R���U�\J��9�+���Șҗ\�.?(����t��ڳ�F&�hG�+
� g�Wk� N �ö���`����Mh8�Ts�,�>vu��6ǜEO�����m��^���?p�8G ����7�u Q�X����6��kD���ǘ�6P�ߺ��[�Xc�,�E�[i�m�G�����s�v�
�sp^(��v�O>�$�� �d�cm��V<8�������/��_�-]k8!�f���R�4#`���-rK�Ǩ�����w�sj)D,�YGL���a�ɜo�D�;,�l�9��YA���n��S9(���v��Uh(�[c��S}�
.��58����L� K���A3j�ٹB[@g����&h#�&8�pn�|L�����ish0;�+x�ԤD'�����ܹsR ��RǏ�d��A�o���L����_|�n޸%*�V�h1�S�$c,��+/���z�c��s�	��1pn .��߹w�}�k	T͛�o������3�ց�����i�?�i�y6xR��H����u���'N���w�y���^�Z�m�t��=�Údd�ߝ���!b�F���y�_��� mYz,��w�@��/}s�`����_8�#?��O)/v��u����)|����P����l�J-9��;wiH xm<~�q���/�W^~E r�B�������` ����/8A�ǆ���_��]8��
�G��}{�1���E�dD�A]@t�/D50��Z�;���B��.�.�M����\GL�O:6g	�1U�f�-W�D\-}mg�H;��Ռ߸���)w�� l�k���.,|���x��]{�� @�� �A�WR�E��`Ĭ1����w�s�7t�ا��r�ч�]������gd�S8wx�)<{�s�x����(��]+�f�U���;w.��� o���V�j	7Q�p�06�ʵ�9�1��	�8V� X�~ܦwrC4ci�0�޸.���e��]��i��O{@N�D�T������b <x����o��g���qO 6Hɉs=C@�4&�4�i'���H1��Iz���`Z:%�o�,�L R��w���g�����&;]-���
���!�#���e��υ΁rC��W�$�7���q�?}�X!�tF3Ŏ,ٜ4��dS[]]O�٣�"6? \˩���}��1��;�!�{@e=����}f��1>�S\Y{���1�a�� �_�h�;6���hߋ����B�� ɇro��=7)'n�3�`����h^A/6ys)�2���u{��?��A�������~���<t��Yq�`�*CD>><ym_���t���X!`#��]��b>ݻ�H^�H�P��\�oM]Q�J4�������4JѨ��D����̴ԛJ[�V��Æyg���7�M��b��l
��&EP<|'�8S�5�sc-C-׏� c���t"���:�2V��O�`�Z����@�'M�,����p�
�  (��?�O�����s��~(�;���_�ڽ����O�q��ܿ��8��~m`���u��^u'O�2��u7�3��`������L�p�ox?�8���e�p�a�:��n�lS_0�+��j�kYw�����,@�]���u ,����[���1�q�!�u�)i���ݴ
ے��%��G����7��D"L?7']<lҢE��3���`�򗿢�ęg� �c,$pI̋i�,��Bs���}����A�W�'��؇p�}뻡�&#�r��y�ԈMVL�[�#���� ��*5B ��1�8L�U�	����V��M��c�?�pطI�7Pb�k6���PK!�;��Ҕ�ZT�"�
���!"shrr��7�Ƹ��ϼ�?�R�%���T{�� ;���KrN{~#Rʴ��/M��"���>7V&k����C�\��2�i�JR��0��ס� <u�"pu)2�z�4]��
@>64D�0N H�͡C`��(��9�n�.z�fԲW���?�F��x!���N6�
�߽{����_s����+���F�JۊL�vA�沾)&�`Ki� �G��Ս��t��=��`�Ql�g �=ش�E	�����H�e}]����T��вz�o�p�%+]�"/��6���n}}���kg�;3)H���u�1���uټ��Ң�U\����!u!3jLp-��UO��
:��vEkz�g���,�O?�<貱
7���Ν;� ����Z���#c�Ӑy�0�d���kf���9>��#hC����`]��p7T
�ǹg���9-�쀵�֎�~�``]�@���)�$ѬM�"��������*�f�'�צ���"6&�[! �К���|��c��z�ܻ�Z�+�u�b`5F0�*)j�V�Gi���v�C�r�{,H�`��(��&6*P ���0�-����k�="�Z�u�4�k4�ut����(�Q���X:��ma�5d�FL��6�e�:�a}�����g�!N���
s��ַ��{�q��3�$�W�M褦`x
��3g�x���6T$�2~��kҧ�C�d�X[y|��H���
�#�k�H�\���p\`K���w-{�:������p�	�~��o��޹u;Ћ�V�!�h�o,rk����*y����n!�r
-Лd�Z'�x�}W["}�� 
���7�W^~�a����r��6o��E�7^ Hӂ�����|�ؠn{ ��q�{$R~�)n�R���&8͵D�pMϜ>͈,6�����x��LK�0C�����!���<C���t:���@  Y�c;�1��f���<��7#��@Z?�&�����s�ڡ<V=wj��(�?6�B�i�]��_v��+�s���!h�����6��s��D?FĔ8N�<���02��I���"1�����\pw��bԬ��w�FH�GT���Aj��p�9����F|}X�����?!�Fҧ\�ң�N�����Gn��)�c�+F�g*
�W�����lot�=��E '4X~��^9ر}g���c��
��٠}��恅��^#�b�ƚ�m
��t4���G䠫�G����UnupI	nۆu�=nfn��,F��؈Z˲;�K�yׅ+δF��)�|�(�����B*{׮=���`�A�݄�M�%����H�	�HQ`AR�
�Cʉm����������#���zl�c���
����irv��Oy�v��r�0��&�����w�nx6���4��֒��Y�v$$��L_���ٕ����R�4��^�㞀���]̤����L@M8y�{|�~?���3��X3��a�1�l�e��`$�a�T߳���,�����Ç��W�\��͠�c��:`�ݳ��}��S��ѣ�RE �!=G
��6�� �&,�2`ì���'< ���������ƹёj\ �XD���R��BŬ1��>j�lױ�Z��k|z�/���	���:|2�X�T���*8�E- A��j�+�yԍW�'ڴ�ֵA�u+eqpS��>T���#T�\��2�Pw��ݞ3�Foj�:�vٟ�F`^åҺ"���u�\K�5����]eD[t����0~���^{
�WW�#�;�9��.u~��=x�U��cU��ܩ�5��L��b��#�w����'Є����y0���g��`O`7Y ������+�>�8�4Q�Ö-�o~N��۔ڀ/��/>��}��G�w ݔ��s��m�̤y�Y�(s-n�4�8wb'�-�춲Sv�I�|��C�&R8ů~�+FM�y�I��`��������!W~#�ꫯY`��O�x��>\6��b5��P�(Q�;���С�_r���i�12 .6Z. �7�,� �>������1ϋ�
"T���dU����5&����o�a��0��w�P����0�f�7�q���Û�I�׌?�0GR]�̕r�d�H]��L�"� ,� �xrR���\��ȟ[�8٨�_�JP?���$��H��xX�D��,AM8z����K���3D�P�r�{�0?u�)��7@���.z����߇���[t����M�^:XV4�7}�k���ٗ^�}�� snq����7��g��WH��τ���{��e\/>��}�T_�q�]�r�}��g�g�￺{w���f�x����DU�V���������������h/���(|���z��Z�x!Z���cGV#�y?������hc݀�D.WV��{��=���K�B@�d�^o$w-�1��Ů�;��v�ڑ�������|�Z�.��?��X�Rx�S�p�>��{�3��<��c����໌����pm\d�|� �����<�X��\D�!�p�b�9s��S�C� �~���5ߐg�s��s��a����ܽ�x�����[L���ꕫ\S��"��ak'ӹ��dy����*E��i܅6�G����A���?{kٛ�Qِf��X���s�7�ν�����K�T�T|0��ʀ�T��Ù��jBf����rBg�?z����������_>q�˴� G�����K/�7��{酳t�8KQu)�<�&�tme��!3�U���ڹ��={�Y���_Q��E���C���A(w���Y����L?K��rf��QU�'78I��_�H �W�����4q�m�s��{�0�K�!��6%��:,ڔ��4���$���R0V9�	�L ��#cGp>1#�>)�rV�@�*Pry?���ꡣ�J����#U�!0*dľm�lZ�wH��6lƃ4I̬�ko�	 F���:�6{òWJ��>�Vt=�P���7:�" v��Ѳ^0�v��]Kp��վ�%�թ �p!b��u������O��n�V���l���v������\��O��{��W��'����ӆ/8O�+�%AF��Q�l�`���Xs�k�ɵ�_�������>=�l(���{ꄘ q����! f�z2���cڿx�=�(���!���3�Y$�P�k�c5o<J�18�8>��s�i�g�=�7�=|��^x����ߧç��Wz��9��T4�T���ƱLE���B<��K/�$ѩ�>S`KK�BBd@��g���us�DҨb~�63Z�O���Eu (x� ��{I5u)�'9z�>�J{�B��c�@TE���/�c PҖ��3�V�i���;�Dd�5��pS1�%&G�ӟ[@�5�϶�2�}iɴ�����mஅCV����(��l�_�$���0F���cMI��E�K�=D����k�B�"��:ĳfH*C��c���2�/�
`���q�P���K��B�)��>�kn��ZfH���^�k�֤�| ��W�=q�۵s� !���|z��Bzu�䐤�l��v���2���:�{w��(8k�2c��ǵ��L��b��i)W�Vl"X;�_�Q�FRѣA���Y�Ϊ�v��� ��c;�.�;h�0n�� B�6��^Y�_�A���~�*�����kmc������,��:�lʞ�JP1;�44� �؈J�Ɩ���d��y��)-9�F���;��"�	J�C�ݒ��9ԡ*Gѩ	���}��D5�A~�)}���Ţژ�5?<#c+�Ӻ�9ͲƤP�"*i�'�l>s��
�Ҳ_xƧ�z�}���`�5w��S~^l�I��fc��T��c��~F���k`$M��,�y�f�o���3>gc`Ξ=����;�`�0Z�Ev�^X'�$� 6�	�,�jc����<�ԓ~�x�����ߧ;%�/2��[ ,T8	�%�+O��&�L�FIW�C�+�2�!-3�"*ҍ2�mR|^��`Ŭ�Ɲ�^���	](�:���Y{Z��Աx5M�%F���̢����^��o?c�'�PB�wk�U�9
�^�Bc(���\�-�6���ދ}�E�[�ʑ!H���l�8�9C���~�yԠ0{�O=���N�:Y'�Dp���v����Q G���s���?�������`roupv��p�����:(*
�f�F�8h�ߓ�J��̑%�N�`D����_�*���3�o��4[�n�Φ8!�$mQ�)���5�umIz,F�2N̮zNƃ��6S��i�J� UG ٟQ�ڣ92�O��E|1�?$2�a�qa4μ��{��	�Q(R� ��s�y��������"�&м��9�Ll)eD��A#m�TC�׏i���:ō�׶�$dw��<T/`zJi�ԃ^/<:��F���~�;��?�1T��2��Ӣ��6GΒ�c|~��'��6�ݱ3��+vx�>3���?���s�ܱs�Y�ɹ8�X��Ɉ�h���<�~��Y�(�9fu�[�����	��E|�B<'iE-�F~��n���F���@�їND�Ei؄ތ���n���9n������yr���k.r-eA�����ļYqoԵ&QSI��8y��2F2�rP4`��3�1�'D�p_p�z � T��� �s�����uD���g1*���K�ғs�,t$����c�y��f�D�ʠ��-.�'��t����+�s��"|��85��B"`���S�`ӓ�e7� �t����f��t�.����4��Pr�C�������5#�S��	mr49�C�&X$<`�mO#/�(���x��\��(�V��dQ9up����-r,�vԸQ�;4j�� ��ڂ���~�m��o��ǧ�#�@>;�?�U� ؔÞd��;�4`��T�q���Q�SD�|⤛_�w#o��q��gt�^���o��<�E����]C{����Q�z�Sac������r�t{���ŋ_I��:�=U����L�S8��~��b;��Ü�v���E��"�%��L>�K�6�{�h��v�P�m5*l[���cƛ%��3u\�"!�nW�s+NG,����D�&��I�׉{.�rݧ�^8����}��#�9P��[� ��VJ��b��Y��eO4{Aɺ��&兦�FYp0
:��Q��|-���Nh��ƨY,>f�^�[7o�?��O<��~���,�������������sZ����ҥo<���۴���>;��P�YMʓ��0����� 7���x'�[�x��N	�0���(Nп��<@ acm�͸.^��>���g�n�m����(>\�+"����i�wTG���v���I����}���.z���]���  \��Ո�bЖ�W�W��^6.�fX�{��'����6R���2��[U⾽�ݎ��AA�kw��'����g?���$a�XY}��`�'z�H=/�w?��ܑÇ��|��E t�%��D�qD����(�� ������u�f����P	L>��T�:�<�c89E��1�^��>�0$�jS�P���<���s[4��H�na�ȓM9eR�[��'[v��t����p�!��ڮ!�lð��O�� �\�KT��s�Z�F�J� �--=r-zן������w
�Gt;4&B�/��P����wθ������	i}������B��~n��������7o�� @���ٹm�����# �G�6�1J�E�7w�[]�[�P^�t���mox����=z�D�I���j����` �*i�;���������]w��U�����
�G_z4q���������q���#��6��,��s��Uɟ��<�*�|��ȆE��7�ErNo`Ǣ<p�p�Y�TH�cs�_,I�ba�9M)�c��ʵ%�#v��׋M��jx�5��A���C�,�r!�K�z��
Dq#
�0�#�p��V4���c�Ն�J5y���\���2~;��GH�������A��5�ғg�{���#���3�πؤ�uJ��˪u�ÜL�ob�yV�H�!B�c�;��w2�h8�g�<φC�;@+ H�6𒲖���	��}�v��L> ����'?a�������� ��gU�Ӣ|b�������+ ـ}~>0E��F�4m0�$t��1�v��Ad�	�:�pݿl(�M�����z�<��w��J�޹m3,�z`�}�][+i+M�XG�sܯa�p��@�=s%הMU��+\�"�P�֧�!G��x X� D�KE8���-EJ���K�t�;fi�ގ++�1fT.Z�p�0΋�K��Hg��{�_�8ΰ�[mQjК��^G�x�����/~�������1��E�6T�ɜN:������d�0fX_80�f�޴���<�|��/~�~���s�A6��:ɴ��Ѓ��j��"DG�������@6k-���/]��)��k�,�:~`�QD��zmv�f�4!��*B��J�����3Tu�+�
�q�Z����T#0� ���Ϲ��>�a�J�u�,E/���$�����p�-���s��������3���_]t���o���4+|��t8�s�=:�A�c�O���"7�B�PS�C�^�Gc� �?����0	O�8�+�*�?���P�iD3������<���!�U�����Kۥ`�)؍��C���tnjB&� l�,ꨛ	�q&I�ʉ�h$N�V9�����&%�1�s�s����3�p�y]����o(��,"p#it�v��%�����E�i�,-��� ݹ ,`�E*��\3]ܘ�]��>e��X@�@�Ş���@:�zsS��پ0O�8� 9������x=�ϫiPdDL�~���"E���="U����\5x��D� �`��'޳g��{�V7V��e���d-�PI�
�?l�X� -�N�Ǫ̀��YD�77<o|�*B��� ��Z*�L�i�����S*��t[#ݵ
���I��C�2��\"��1��)�7�)M�����[��y8��d�[�M�B@	�.�]~������(Q���o�$�2��r"vo<���u���d�N��W������|Sp��_y ���`dלy�V%_�0�g.u�E�96������jQX݈�"r��A�i��=�GA��] �8�s���V�#7��P�_UE���^�&D���x�w����mbb� �?�AÎ��~f�y'c��JD�5dƪ��� ��N"�g�.1���`K���)N�?5
{���3��H�Eu|2#p��:f��Ӆ�$�P'���l��8�lYsƄ"%�2R^s͘�6�<��5�j���K��:��W�t�Z�������@����p�dXZ�{Z#�I���dϢ����&�.|��smmCZ��L�Ӑϭ����X��פ=�ݻ`�upW�Y<W^���^+�Oy�ѐNR�xM(i��J�K�Ơ��O�����^=+ީaAq!riUSy�-��]�p�y�dmz袂��`�1��l�x;gQ�IA��#+6�S���G��nH_�0ՉJr-�OO?�Z�_l�\�pY&υg��/n�a@M�>�E��.�<S��>�V����d��0G��� ǣ���Ҳ�Ȯ�/����Xp�c�������y�ѓn��2^��(Qex��#�����.������~@�y�������~LRD���*dC�@�y�(��txkm�i`7@��s�,X
g� d�KS�xZ���sA�Xy�����i	�4Q	��I�]������w�	�8	=e�M:�� ��,*���.�hU����g�l&(ބ�'�$-.`'����^7	r�˙,ui�������:=:O�6�yMQ�w��\/�C1O�Z�y��A��`v�����H�L�i;���6BC��(HИ�Ɨ�7W'jڄ�>(.8˱Х}�Ӳ�h�+`�֧�-��;n���3���2#S����E$�4�;s�K�n�[i��l��-�jivJu{AՂ�_:Ơ����� ·M�ў����;��@��e�󛟗j�Z� I�w6�  ���ȧ+����{��i�[�ɒv�rZ|�~�@:r؃��Q���R[�Ln#D}�ꅴ{�7;Z e�d�t,6[�Ngl�l���'ٝ��<�5�+�hpPv���q��La��Yl��M�VWHA�X��+��C8�l�R�����ypRl���^+������t�)�~c^�s��&f4�V���#�:�B���ye![Ҭ$arԔ��}�v�bݒ`���nW֞[9ڦ�3b�"b7d3��
����2޶���isH�*�[�v�!M^A26��hl$]i�V��+�YY�l�)��M錈�i4�"t�R�t�<�*� a�e����k�.3ZBy1�H2�vY�kO3~��iVF
Ǻ!�1�̑�X��K�N(��O�l�#M�����sM�cB�T����t�x���&ZUF�D���#�n�/��ʽ:�S���[�L�v����pSF(���ۗܲ�59���N��@@^K[�B���v�C�͗"^�2�͹Ȁ���ؽTI�Y.��<�v�J�ڒCf�DH]u� ���p#��i����\�]��t�>x ���q������̲��*���4"�x�EE��x��P=Zf��l��0
��ǟ|L�!��a�Px#""����@�� ֎����O�n=��_�8P^����� ]��lRd�m�"�P� ��Qs��ѐި�ѵ�T�bZX$?�fi+U�U���"�6G�Y������+
K�db�E馡LKZ�k-h#�>�(O�	�6��ߴ :��l��5�Z�s������ߺEP,Z ��g����� ����ֲ������n�N��^�ys�?��A�K�s!�4b���&! #l���-����'?�)�/��n��;�w~zf�t<  tr�#�B-�ń+�{��N=��{���Ce��6�'k[
>�4���i��פج=�nʂk Ŕp JJ�cº�"��_�����p��>O�)�\P�	.��>gU�,(���!�g������!Z�Dʏ���*<�A�6� ��M�%sp�<jc��;R��C�to� �"W�Sh�Pz��Nna���߽w7A�s�>KۂyQ��^@���A> /��ho���n��`�-re�l����a�6CT4��aJY�F�:F���a��B��MS�K�UK�*$2!^1�T � �0
�Of%��\�b���6�
����{���V�^��so�>�:��<�[I�E交K�9������k�C{�����2�7M)���ƚ��N���B4qc����^]��,Rʅ�=����@s�S!���=�˸2fx��K����<��t.v�+����vYG�J;�G5��>{@�7�<b�i����"#�������eAK��N���W�m}��B[[��Ŧ8��L�\�\�L;���f/��Qs�2�Ƈ�s�$�*Z��cgRO�Z-��=E�p�,o����;��	��L�ݿ9�����N�龴��9�ؔ����B]j������ϔ��� �Z�A�Ԧ���V��OGG�w���`�hji�C�����lY�'�q���v4[V�s-�Qu�3�1'^�[��^�r��(�Z�!Ŋ��'?�O���` �JxH4��j�"ת�ر��bz�=�ٳ���~f��֐ʠ��jV�tI��:6�SJ���-z+Ǽ׌TuG7�ڊ/8Y
�f�0��5�L�$�@ C�@�d�Ƶ P#
���a�!a�������	��&�<L��:T٤p���<Oy���,~J@����s?�R��ãwh�P��+}nu
 4��z�M�f��1�~[�W�st�s���,~�I�(79Fv�06�z�O���k�V��k!��L�=Z�k]|L�\M\�uJ
雔���:	Y��9�K��#Ш��C��zo�o��_�;���.Я|�@�{��\(R���ddR��ck�i���8e�Λx��9��qF7��{��ey��T�s�ԅ�����j�h���N��2�<Y�iv6��B�5�s����lzn������#`����k�k��g�9�����yp����-䛳�:S���qee5H��:�y�۰��܅z�ϴ|�X�W�&�񐑱�hS��d�F�OO6:��i���I9累b�x�Ql���z���~���e�1�M_#3v]����Q� z�������^�3D��~n�N�=�To����a#\s�Ѫۆ,\G�-�N��u�[z�V%�u�35�匀}խ�.�k�柟�K�p��߾�y'��O��GL���ݻ�[o��y�+���Wn�j�Xu4zב�4?��P{�X�B��b���m8��4)[lw��Z�H��(_���e�p$��y#)�*(X����B��cbZ�x�e9M�ASh<�l�E\-�k{���uh�21�
�6F�>]*L>�Ժe_�C�H?[hzI&h�!�q�9o�q!�bL%�Yk���'��J�#CV]s����Ci�l�&��x�с\6�¥J��"0o�I���}�+�_e�,��O��B=���0�D�%�m�n�j�B��P���γ��5U���+�3�o_��x�O<!m��7qal������P;�`(z0qnQ�#)UXڼrX�(�������] [lB�6����PS,�ܸ~��DG�MK��=���'��M�J�kyn|�^�����������g��h���Cnd���Ly��8	LM����&�a
y��ٗ4kߐ+Z��W�&�+��nEY�F)*�7����LyVm��`5�[	OZӦG��4.<'� �?$ib�Y
�"���S#�T�!X�=����J���9M�Β�pC޵:;&�͈i�m�A�&a�'��Y}Ul�z#$��F���J�TbL�A�o* ���3R���D7a<js��5�a�������粠�Ɣn!FseuE�t!
3��> KS����v�:��!�g�/Z��1��r��)��D��
|y�{G\��v���&����49�#
GwV�^-�`6v_lo�*��T�(:!�7)�����[mQ�$�C��ҽ�i�96�cǎJ�+o�-:���vv4�ɦW$z�2*��T�P��*l��}��^�ejB
��n�����u��U��:�<B�h���`�����Z�Ɍ0 ��I�Ut��<��[d��j�`��
 *s�5�dj�vVacM|�f��4��ew��U��`��ר�֒�X�۽��ٲ=�P5�� �	��`�!`�Jױ�a��R
�����|LM8�˪�ِ�;n�������C&�^D�� ���*�eK�9��x��*ϹA Q�Z#���z�K�k9H&��Ӗ�> HC�U�
���d<A��i	�M���F�n��:Mp�!��:�G�wM&�3�~ȆY�K
KJ������Qp�T����@L�X����@�����S�
�"�m�+��@{[`?��*�/�k���A������L}�XY6%�	2
S I��T?��QՈkN�QCfBje��{*��X�p�������|Ώ����e��V��i@��%��O��ۉ2�W���D�����n�H!	 8V(��6-<+�2z�&4�>a�5
��,�-�Q�8��Uvn@"��k��@;&�
�A��9"e����_&0����yi��Mv�!� ��{�\��*��!�RG+��<�B��@〢�|�Ν;Ǣl��|&"@x���#-���訔���:ymz�Ky���Y�?g�)��5ɢJ7)�����1�g��:6u�mh� �`<6��`ˠ4���"��&�X_pl��GAx�w�*Lkkh|�}�즛 ��20�55Q��Ao�B
H4�kf���"��PЛ�t��tT�Z�Jz�]x�(�t�Xf����| A_�����m
C���n�"�h���� �L֚Hp	G�ED�ɕ6����o9RPD5��u�/l���7���*T4��Hy���u��TN���Z]���f�55b�F̘�_ƻ	�&Ъ�	�a�zl�����׉ٙ-����
 c$<iH`���&r���ڊ����t a�0�q�th'S� �6�%h�ٓ�e��2��	�;���k:nc��k�I���'�X�n:�5��P�d���D���(@v�e�s�c�����Z_[a�?TB:���<uB9z�l:��3`8ҨnZ����pQ��*�7o��f�\]�
+W������A�-vl�p�� �(Ȫ �bޭS�d3l�\X��kk�: �Iu���cP1���6M@=X�r��d��e\Ȯ�8L��ݻ��D��5�̮��D��E`��&�����.e�e���q!�;G�~��K�C䷖3,'�Rנ	?���XS���Z�n���<@4��4�� �6�� *��.�������G�2D�����<c�Z6�&X�N�oU簢T�mް����q5Lod���Ӿ�I@ѝQRm��vS
��$;i\�4rj��4ymR�Z�@Zi������p������U *-<�,d�E�T�د8�x�R�� 8K�?�$�^�J�
�¤��*o��c�hs���8�F*G4�:D[��#/�����]-�ER��[32�*�.��/z4,�ڂ�5� ;V~��<ଁ3�B���&�����F�����K�ә���� 'uH���պH��^z��]H5�Z��f� WU-_V�g�������-��Ўp}��l�a��8x��C:��RKQ5-Ó�d,�qc��� �&���vO��I�)<s��d�H�|�#�� 2N)�����"r�P���Ї�[t�	�a��h"�� ��n��W�nƘ��Y`-��V����*l�P�����z��gl} ܃�ƍ[���v'�#��y���Glr���)%x�~3G���6��D:{!��y�⓲\�gXу)Fl��T��K�`�	Etojf�;���C5:6.F�=0�t���uJ�� �� �$޻w7F�,���P�]�.�A�t(U���6{�/ݗV��XO��"t^���j�|�D�,5�"��!��� s�5�5�  �&�`���k
��^^�"=�\E��8�l_ܓ41Z�f�2Rͺ*�P�(��\#h��:ܔ�M�(���������2 E�iD4���7W�Wt>���Քn��}���wo���9�wt�[u+h�B�,�O�2�P+P6n�2�}��Bq�q����Ⱥ5�:�=�;����	�|~n���4����i��.����hl��� ��uB{}cՙ���i���e�"����y'jum������/�U St�<��YfB�A<6_��@�T�����Չs.����I/.�C�q�!DgD�b��Z���j&�R,7P��nj��Z����aA8�7?V�nr�G�&+5@����Hf����B��87��`;�<���XT�k���E�_tמ��WP��$�e`t"
g�I�HA?��zl"���v1׮\�������~�j������#����mH���BUj~���A��{�=)T�&�Y�� �؇D�e�E���!d4ؼv�������I�i�A �z��I���-v��B$0e2�RS SҚ�^��&��0 Skj��F1{�H1-[GPc�2xTշND�ަ-{�x'5'Ey�R�W+m��?��wmR�S*��:�Rx9�~�>�<y�]��ʥ�J����N[U�_���h��|^B���\��5�VH�Z�-ei��i���_L��%�U�&?�<�tF��V��Z'��Mg/n�a&L�㱷�^	5=�X���SM��>R������"̓ٙ��CaJ�
�6Y��s��H@G����D*�xQ~,�Ð���ϑsZFm�D�}A��f+���ܒ��Q]oi��w���Y��=����bCN��" �ХFKc�L�}��]I����s}���Y����������+oox��Dv%򕩠z"#UmM���K/!�F����³��݀E6؜q
��u�;�iH]e���e�ܾ}�ݹs���_+��.���I;
Q<_De$J&
+���"TP
����s��hk���&Ю�f'9.kF5�������  p��æC�4�)�{���L|@��@�� -c���"�D�Q�X�>�<����
�۝!���W([8R #��r�+-�a�,�}g�O3��F%	�JxX����"#��N"�r��C����s��(6���6}\��}kFvBs	�6�2}ar�[x5�<���̑ٍ�Y�;u*�e�r��hÅ�V-H��!�����;F�fJ.y��3�j/Qitx^��o�`��ZY�W�a^ҙ�p�;t�0�����Wj�^���><(yFG)�ҝ~�v�`B�����s��\J��0��#M9��ػI�����j�΅Z�Z�q6�>�-n?3�u����EVbu(�0�	M��(gt�NQ��;|��3͂��@v���CaT
p�t�!�D���甕pj���Â����z�@�Ϋv�-��%[Vc�co�
�V����,��\s�~�Op�R(���S�̟{wyp*�ܾ����c��I"mM��`�AY`��^p/�|��ݳK�Y���E��v�: &ug�G
��iGu_|q�;��ʕ+̙Fp��6�w�
��66nkj��L�A�v��1F��t�0�7�K��A������`/�<MBB�-���v�u�Rk�mg�XԔzg�x$�5!�m����o�/,�~޹c�{��3������1T�5yq*bS%S�o� h�+���f���Z6ZU_Ć�ۜ�O�YK��ӹ�&`�(p�1l����c47I�*�
��bT6F�E/��mG沱E�����M59�}��\K�2���D!�	��P�Pi�j<��*|�����E�kX�#��U�����Uww� @�[^]���pҳZؒu&��J~�k�>xSH'�w
�n�����S��K:�	��7J�wλ�7hH�3�0���۷�0l��/3��Y���qm�5�I���[젃>��|srq 2^�r0��+�M��H�^b4��Cs��=�@O�:pk�F�cj��b���.^`��T(vl�r �a������*���	)=��!۾}�ZA#�(�5�4��Dzۆ{p1T]M�q1n!s*�������y])��F��:�4g�ѣ�uF�H������&a�}` �s��Hf(�&"�Pn֫���2V��:��^s�����:�@Y��ƺQ���1���q1ۑ.�[�-��9�,�o,�;.�+H�T����L�8)}i�P7�����5ʕQ����"���N���Oޓl�,�"���g��;@|���wH�yk��-5ڏNd���t��tr<��� Z����~�!��'Q�"Cds�B��R@J:��E��͂���w��Q�� q&{lE%{��d���:�f8QǏ��9�+�I����̏x�m���I R�j�y����-|ˎt��#�bhSxJ�+��J֠֨o%-l�؂�9-Բ�sӌB���H���s����~�z�4����QYǹ��
��}�B��z�B�`�K]ZHg�~���{ܽ��K�W_w�D�*��dǳ�F���6\�&�C���U�.2�qK;SJQu�^,��4.* h�g\Ǯ�;ݓO<�N�8����m3I��X�˵%ݜ�5uރ����ݯ�#G��=���:�ƂϨ���p�E{������X�7���R�JUR�����F��E�� 茽��M2<��+K��\`�w�����s�߭)�'�q!%���V�����o-��t2|��$ܟT:�+Ka��bDص���\j�'��6O���Nk�e[��e����p�BG3~OMRTr�����c��7<��i][� ��"�-�s���Q ��͛�b�o�a�wA�sM��;v.0�xǿ�����}�a���a�3� d��u� ��1h�s߼��� tz��@TQ:JZ�ʕ�n�!)�ቓn���l<(z�<ػ��_�)?J@�\��TQln�\�.'6�[�P?��9����1@�߶m��C���­�Юxe�@�������m�o��������kW9�"g#\?؟o�����e��������]>3D5\3y��p�m�L�� '���$���V��)~�>�=����8N���ʠvԁ��Ι�]M��T�MIpn�b�\ ��p�|�fN�/��ݠc%`
Ŕ�� �t�ø)%_��s��� ���v��Z�,��a �hk6�$+�p�f��8�h�+cTZ߇�Dw�۷k'���Q�H�s� '�;��mE��C���g�S���T���v�Pz}��V��ΈIH�c�C.���6���Z���ਃw��a�[ ��M?O����]][�@�kϋ���ttH�ŏ{����;+�hΣ��Xw����E��&�n���|����{s)sۂ9��{�)�8Gl.��v���h��a,,�%��� 	�b��[v�����gs�
O�}ŀ1�=�;w�����ʕ��)=XЌW�	�8�@�[؂N!��D���rX��eJ���m��HA�b3�v��scW�:��B�Z�^ �!{PO 0�&~�2��ϓO�b ��!'.��\�[�'Ex�'�s���s'�w�?��;��9��V��a�N(��o96���`j��&Öʒm1�Kﾐ*CcXHXu�@'Wp�7 ޖ���4R3)�	�p��%�q��\y�&.ώ]=��3�g�)���[��,zD��Hg�Զφ�����ΝcD�i���MpR�5�;3���y��XfM��6�-�>r��)����4L<��v0���I�8�5$��Q� ���dJ+<v���k����w��?;=O"G�J!<��#���Ƥ�������id�Ѭ����~�����/��p���[��Э�T��%�@޾q�}u��[���SG�[4�kD`����������*[C��Վ_k�|}���s����2�������Lo�@d �`z��M �cb�O�Q����%c$ʹQq�a ��Y� ���<�Є钬�d��1IZ��ݳ҂���C�s�g�����w: �l���9�H,���y�@�C���OS�8@5���/]f��eQ����z���h0~�3BM��:y�%R�����f}��B�^��M��&�)�:�ܹ����ۃ�#Iy����g��ů.8�:׸λ;�����a����B%���A�Ӛ�T4e+cck��D+SW`fY��[G���]���B�,~;�No)��W�p�g���uX���?kS�i�~F5qO��?r�uLխ��j&w�voG�S3���9{[����?x������9�����]DAUBw�?��C���_���y��E��̐x��wg,��}C=	��<X�N�b��g�y���h���}�b��������p�ʥ �L����� ��P�����h���s���(�d�@�jT ����L������Ժ[�M��:3l�+R��U\]ka{��gϺn9�P�7+��Y!�8�"f8�J����@je!�w0��������~�TB�+�#�B��;���5E����	�_�'�ߚ'���vH�f��w�ϵ�O�?�mЬ{����d�����v��򭭋$9��������*��mam���Y�X �c��_G[�p�����:���.X~��n�����>0`�Q�4�>���"� [
���:E�B5��[Ѥ��m$B��F�; �00���E�iD�Η�5DK����={v�g�}�:t�Q+l���4�Zт���Z2E��N��p=�y�i�3�1)W.��j����Fv��IZ)n���- �M�_�3�P7�f	Oʨ.�ί�=����B��1:�'%`�D��T6�@"��/k��EN����i �l�H��6 Cz��74X�w�:*�#?�v�Ӱ�0��3+oF�pv�
 �"4i�{@�T%�ByC� �$�֑f�� !��먽���I!��"�D\�$o�qNAۺ���6>�R�+ yk��[��5�7e�z��Gx6 ��B#����ڀ"]��撂`����g�R4=?H���]��Đ����A��\]�7X�ړ>�!�������� 
� &5M��p׮_wW������;q��@ԃ�׮3�Bq}<��Tç�s�Ɛ�� `�w<O<C�9Ƚ�T��q(���/���Ɓ�����`��$v�I��LuuS��qG$�Ңø��5ek�H��U�[:Ť�����g;%0@3Ha��3���׃�^;�!"��).��2�u��$G�ɵ̚�!��]ꈂc�nj])0D38_��(��t�fݸ�71S{ �]�\�>l^�E��k0	]	<s��?��'�y�O)��t�N+껤�tiG1ϐ��l�_�OK��7���;���W�1ݼq�N'�ߎۨ@�f3�0X�?���:�
yFn��+ Ӏ���vq3�R���}��ϹSO<���@���`5U<��6��N
�l�j�z�ڱ�a�]�s�nࡷ�C#Śp@O�<᎟8&:��ZQBP��ҹNZ������n��� A�>?X^a������[�e�8�����֚:�1:���ѤC1A��r�x�P�`���:c�ԬE)#:W]c�bF�4���#�&vUs��n��?��W�%[B��0�h�(9�NKk%��sG�!� {i��&u�c�A&d�Z�ϲ�� \c=���qѶ{JD�����+ۀip����0�.H�d�:Y��-���q��qv���7�UF��J�N"M��2%�<]���6g��R��v�H��-j`畊�����iE�R�kU��^/p�'�,E�/��]��:�ۓ2j܉��Y�nMT|�����c��#�pM"H��xM���r � |�ɧ]��b����<Sh.""������C&�0Dt; ����Y������Υ���j�v�����̰��@�P�Y���gD) 8�Zx�b�%F�a%��	��/���1��i̻��ﭣ����>\��:B�rW��\�F��v���m66�3}Ɲa�� ��n��(��A�J�Kyp:P������*1t�yr�!�b�w|�u1Y\(ȓ�(yٺ!Sw��7�R�J�9�n�N�|�.
��PMSK��������wn1�̮fN���C�N�+Bc��b!����d!s�Ϙ�C�R��YȘ�F�g���9E{u�E����� wV�g���OkV�a�F�l�d!��P���B�l������f&��V[V������{��Ё��xe!�0����V�%-ھ^�øw�6h�����u���\�L��B;�N&���.f�jf8iC��m"/�h��)�iR���ӯ��(|u:�S�[*��a_p� 1Q���c�܉c���>�Ì&b>YĹ�σ
��lSG�
QjrGu�N�l���!�l���罣.�yHGL�/�k�(�͜�z�M�����(��F����&��XI�P��-'-j����ܻ�����w��6˷�z�e����^���=��N��-�]��D�%B���"��K��kAV������˿�����?�"N��=�Y,m��HU�Cd�9��f-,��5����pˀ��k~�_΃���։C��tF#ܠȊ���v��t�#-�.e^7/�Y.^���ŧ�ǅ�l�#�'��Hr�w�o[�1�͡U�T�Jy�TO��5Z��yfƱ��@�ɧ��^B��0HJ��\""���&�M.�_�4��'�����Mxh�ZB!�:y42�%pj�ZeG��Vu��O����g�މ�43�g����VUm�]���\O,, ;!��hW{�ߪ��iCX����f
ƪ��X(8����`z@MC۰�I�u� ��E|ZR�����q^�1�K�`�R!D��k�Ql3~�g�%��S5V�6�����VV͏m�{O;�d�q��B����"ua<�禔o�HG$b\�|�\ʾ��S�""|u�%�TێD����!Q����dkX~ẚ:VcK��8N�]�:C͆�G�`�i�L�B�M��D����N�j�:G٩ UJ��r�#&��ϴ-0��s�<D�DS��m"K�$'�k���+mh�A����"�{�f�me�v�*�E���Ai����zhހ{�����K������ ��hwZ�g�����%��Y�K"z޴*�����V6U�8g�w�(��۽Ŧ�`���!mYEG��%B4X�Ph�,S�}EZ��陦�O�6
`s�@�bMx(P�iw��G�DW���Vڏ�#�����yIU���,F��ϋ5pC�Z�B��1:Z�
~�qZgj�R|Z��F�a��]��T�b��I�\H)�B��	:��
-�isқL���Q��6��iY��\�MHW/kRx����{�H+��F�	�JjRK6,H�$6� @�b�h!Ai����! ���B��·��E���GO?�E��K�⍠t��w��3�6�8v�������֙3�3ky��S`��N��`^'G��GYf��Fe����#��2xP�]����]�Dd� 2�n8R���)����5*G<��s�?��ܳ�p����m���}���H'�8OQhf��3g��B���_���i%�a}�����{۝y�{l�~7�f�`N;`�t0���}���?���0�:�Ƚx�j ���sҕPO���Q<f��"����I�����6�:��DAo~��Jw��pZu��57Q�Y�VWe�� ��]�Đ�}�~h���I��܉v%�����b�	аB�U��vm�2M�|�J>W��H�kQR���H$���Zŷ�1o��B��H���)EGr|�d��uև��6H�a������<i程%�c�$�2Y��S�fcbm��H�^�t�v��*�$mD��I���=z�-j�ܹ�Q��F5��ƺ��ۿ�Ք�r��Ɔ�M��%U07;C�ա���6ؕ��H;�5�ܡ
�믾v_]�����k�m�㚦e�}���cG���d�aإ
)Α��4�/��Ŏq1Z&��FÊ����K��>��Y���I�ݲ㉅��&�L
�MQo�(�B7�}�|Ĉ���I�T��tl��o�}�#�2N �z���5^�����"Ԇ��/|9[�MM�NP��X�N��ee��{�fK�`V�=V��X���3��I,6�� ����!�n�.����)���mcaw�4�I�ӖbIgM*/�tn�:���N��a�.��aGVi�W3H��z���Q{#<��Ə����ߐ�����;�ܸ	���N��c��iM�'��L�%�G���� �=��Q��%�+�	 $�}*����;>�_P��+����1ַ��sF�:�Ʌ�da]%ΒEfp-#?GF�,�c���YY�Om�ږR�غ��Qaz�4UA,^l�"75�&ˑ�wjA����6�,��RPS�V�	���+ �8�p3M��y?� ��pp/K��=$�ƶOb6�s���
�j�[
�m�Z�%o���	�5�)��2h�[���vߓ ��-�.��)���M+���M�������c�xbp|�~�i*? t�^�>�tЄ=u�)�?p���݉�q'�#�����&��I��,b[;�2ؚZ�v�٬SO=��~�m��+/��ۯA���-Z����#[7
x� ��J�
�bO�>��������ˠ��������;{�,y�Ȥ��~�2�7�2w3M_J�	0��ʦ
k!c`$��9t�{�׸���j��:*Ȑ�F��W�.�{�{���B#��4Y����N�J;�W {�;��%k�*�/_kS%f�@o ��#Q�&���~b���^� �4���|��Z� �N:;�\%���h��Դ�Ö:����a��ѻh������g0��NGӬ~��d�Fd� �O�ݻv��T�t�����F��߹P(�X+:��K#�x(������_%��CW!���������c���:+th[M�dk��,�w�ZDJy����Ǐ���?��gz����~@�W|�/�@SMj�،d�F��Q�p�������P:ƌE�o�}�����������q�3RQE.-8��!8d�n���Ey�|]%��п�@�t���Z�]�eXΩ.a�S���~�<K^�d1�im���԰�g��/iz��+M�����/�1�kT-O�&9z�nE@o��;�T3����d�UA�a=,@cL�Q���O6
��PK��h��2����c�3MF�FX���)�I�H�K'�:��t&=����3�.o��S�	(��2��X86��Zzډk�6��b;D��5��8��da�����q�1���2���m�6E�Q�u��p��������ˍk���	��"}:;3��i��oQ��N����Ʊ��Y��`��4��Qt�`���D�P�?���7�	�ƴp	��5,ٺ�[��=���f]iՋ��n�"o%|eib �tE�l�
�d��Ʀ���E��_ZB @q�|Y�r�F�9�Mۮ4v�	��>a��?���Ɏ�:ͬ��
4�}W��D�IY��g����'����L�[[%Q�}A�؈���]�����s2��@���	��vUV.�|g�����3]	sJ1�-몹	���n����\3�3E\��4��?���PhTp��I���_fȌ��]�?wޝ:}J)F;���{�Gf�;�wFzƖ�[5<f`�K���c���U9E�Ug'���/���G�/��Mw���+��%�^��ig��lm
Rk�W<EV`��"��7>��C��{?�@���_��A��p,)K�@%h�u��f�A=������־%S=��`_"}�9D�
�n����Ӑ�Z����=pG>S��/�����uE��# �(#���!�e<�6Iѫ� �,�rh7]�����P�~����C�t��AinwS+�['�Ѳ�V6�2���������7�7�I��-$��C�@���$�5�f?�U����݈�28z�8�RR��PU
�RHɒ�u)-�4�
z���L�������ܯU��7n�r"�8�`� �rjwMOM�G�C�Fi��:u���g?��/�ٳ��Y��Ж��.���4\D;:���ЫA�ŋ��E ͎2q#��iI+��7�yP����p?��v�>��RA�$�c���Ozt�������� c�����K .�w?����i��[\�%<��0*<��I�S�C���T%f�/(om+/\\z�K��� }
LCM)�Q�����H�X^�m�:�NV�݉V Ò���E��3��;�f���*��U�y`!=�	�`vS��|w��㛾L�X�8 )S�(x������q��m�0U&�N�	C���1Ռ�L�� ��%^���������\���Jߛ/�Y���|Y���k��Y�z**bx�>�g,�#�FkT Hg�gi!Li��bj�6��>���X����|��%}�R�I*�T����`̣���0 1��_�IEG��PQu����N�%��,���@ߩ�,�g��~꘵
j@��Q/fOӀ�L��2��i\�sf^�ќ(!���U^B&"J����/�EP>u����ZG�̂ M$b���"ӏ�h����+Q�:y����NH���x�C��Q��Lz50|��G���Y��(&����� $�I4���`䱖����i9󐭖��udq]�[�]po죿����x����?���+�c�c�{�[M�+5pJgC�=Vr�.DO~��LQ8�7����*��=��O��ww�-��K�'ۦO�g��8��F�1�L�O�.�$��V��8�~��+L3;x�`�^��%@��R!:3�B���J�����E�
�Kܖ er��'�"^��"����P���7ָi4�P����=�(Lİt�I[p)l���7�a�:�SH٨c-����!��.%�;{���x����5����ݼP���MeI[q"��6ܭ_G0�5C���PԲ�'���,p�E�Z��5(<���Ð��)�.Ý�"X� �:$����q�ܤ�y����Q�XF�����A�Rxώk	�<A6O�%�p``5���W_��{��煰^��-����$�3�&���Y��ڡ�����t�	]�6K���5���������ME< p��g��˗�b갭�%eBBh�¡'tE󺨧�Q��\��/�{B���]gG����
��C���G2�7�Y(�O�VܫL-�>�i����5���H�JZ��[z���6(Lb��#<V�(ӏMUz�]�Y����4�<���D=��W�{*���<.yH��݊�ʧ����jJx���S�!�鴪�qYq��bW�y�h��b?e�^�[Ȇ�팉�l����Z�K#��F�j�L_�?V�M�%�t[��ꣶ7����hc/��-6�9^�t`A��®(c#1O=ޅ���1���M6� 7�XH<1���6X��O4B�G��r�x�%R�۴���������᱖���s�?��;G\�� [s�,=^!�Kc�I�"�Np�6��C���~0�K(���.%����ϼus�KT��Y�����qH��FL��
](�r����ӈ�:\�W��+�sM�g�'���63Q}%#�..۷LM���l~�w�� ��~\x(�@����鳧ݑ�G����}��_�B�����{�w05X�0�kZ�tϪ�,�30V+"3�e5*�0z=l��'#��DǷ�g��iZ�M�3$~MBHsc�d��1$�TPhvv5]�����g�#��u�hX��ne^ �9�j���ފ�yS�h��)�!M۷���{��t{>��ʳN#�I���s���\I3�'��b�λ���as;ʌ�h\H�-�ZN��t�S��`��ȝ� ]H#l���h��"v�	�f��njU�^q;�'�%b���G^^�e�r�o�iN��#h���Q{��!r���3���tw��h�V>}�9�����6vK�������)j�_+ѣR /��(�v�/=-D��P�,;��فc��-�x����d}��˒�m|�Ȱ*�I�.�?-�n��w�ozz��Ѝ	���~F��� �u�����^�M,�OT��:�=|����ACx>q�lI��-����l�5������EU��/�{�O�\%Gv4�5���w����棏>���7��"'L�X�h���D،'�D��09�u#VRU\�>jሗ�N�F�ϑÇ�E�@�y�ǁ�:�ƒ7�q���yǓBp٣T���B:D�r�B���>���U
�Z{�$<s�/(oi���+�٠Ċ%�J<�5OY������J�i W][���X �$/s�?G��x*�^]\"�-�++).�<W���ң����K>�i�l
��]��� �p���Wkq�M�
�ኢN�ee����O��ҵV�{�[A{?l��4J�f1o��W����(�zF��o3����y�y�&�	a0h�7hg��4R'!���90Ze�x�(&��1�2:G>SS�*u�U���&�K���,�� �4��R�D��˟����5�[�<w��D5G�8:����_17Q<�AAAO�>���i�m���>��W�H����̙��w]'ٝ�k#�=2�/�=����wN�|�itMF�l��=�%����*�~ޥ�;V*s��^�^U���h|7�h�i�Y�� ��"� �T4V�?���_�W^�w��ᮦ���d4��ǍC��qXK�Bh��l�/A �}+���|���0c-�n+8
�$��Z��q�����fc�͖��mH��f��X�M{a!�v> .0�Fԭw�ܥb�v�{��f��O�T��do��P�O��a,Ia�"##R�(��oL|
A1��{ߐ)m�qo:�7~��ٙ2�FJg���)�k����>g��pK*_C�)�7꣨��N�?8������A�`�~s��[ٷ���թ�h�H�?��d���ɹ�8ׇvǎ'��w��8l�wf�&A���'��:7,�{Zy_~/$#���r �7���~�<�?"�sd	ʆ��8����(`w>pw�I�'"�ډ��~�� 
��z��Qh�&xZ �Z�.t���to��ٻ��ϹK�/Ё��p�������J�r�l3�b�ɑ���
+|�婧ȓ��Q�I4̭�KծZ=�7B;��k_n2�|W;�z�ʲ���u�t�nS�������Ϲ����D�('�/����KY>�`݊`�x1�i �v�&�t��	ْtX�T�� �s�S/����҅�n�v�����ﻫ׾�ǀ�cj�P�k	��o[�c�{'��哒���k��Y��o:F�"Y���}\LP��C�L�4�d�Է�n��<{��O<��v���D�d��}w�c%��x P�����R��s�U���%O� ��S3��{A�����Ã	i-���9�2v�+�f1W��v8W�K:�ww%l�B��yʧ�{N�,N۠5��EW�OsW��2�^�dt�s�����\����'�A

����*K`���~U�H;[zbu>����3�ͥ����ɺ �Rs�t��`�Y�/��Ԃ��ؾ-U�sت{�2	^(t��J�����!RsJ��s�'L%�q�6�ښl��+��X��m4��Ir��y�:*���&��k�E97F���3���6i,��i��F�R��A�d �ԁ��:�]A�ʫ�F.�u�H�jt̀#������PQ>�FR�.]��^}�5���K�������w��;�0z��5
� p�n�)5����2�'<�������Z{-U*C�k't�9� �v��?y�����J]�H����v��ԿzNhӱ6IN��v(����M!y�|O���]F8LN
?u/����(�ݨGݤG4~o�ø�@K��_xe�3辻��̀Ŋ��)�je�Rԇ=�>9`$R:�R�:����d�� ����sG"�E����� ������|'xH���Q�n&Ǉ�8�`�Qv(�@� �O�j��["о}�ml��xTqG��M�3Z�߿�#��9�N�<� RiI^�`�����I� ��JC��+�ZQ8�p����t��v�Wאr��)9;aF���g-1Yݸ���IY�`k���(C������ݹO��7ǃ�B���R�B��!1���&C@��[�}��&70>�4����Cw'.�h �p�\\��!��!�@0�I��Պt#����%vz��$�'� ݳg�0��c���C@���t������iA�g�f3�e�0�aބV<r����k��S'Np�N�;Ô��V�� ��$��V�<D�2�1rj��:fE9 !Y�PZ�/�a������}�]���v�~��t/�w[���>Ӡ �fp�f>����G$f�O�s�׫Td�F����1��?���{( 7�P��|�w+�ג�2�n���1���޳�`������~n�럔���]S�������'��tfP ��PՒ�j
Jߢ V%�k��՛��"�*����<Ix����atS�]�3�h�Ov�O!���1aͤQ��^���z�������RV:�֚�ξ	�M�D&��P[+G���,)�P�6tw�� C]�E=G��i�� p�g�b��8(1��΀A���GI�X�rƵ�@����k�2��$�#��1��@���&ݏ���B �{Xj�ݱ��(-�s4E��=�������r�|�M�	���>6߼q�m��aG� y�eh��jB���8w$?�2е߳¹��8
ͤ/��z4ر�ȃ��q��y����y����}&����Tbp9���K��p惢3a����d��m� ]Ls�8;/9<n{`6�I��]�7(t�ww1�y!����gz&N���̭Q�&��`F��cvQ]��l�V������i�)���2@��P�E|,T(� &w�?r��2R�дg{ӥm��Yjaݗ�q/��_q#��s�z\c�&"ցsnm�2ia��[ �`*��ڜo�q.R>�M��d�����˨��)"��t��\g��� �'+PY��M�T~����
�`w�.D���=@@�`y��G��0�a��}7�|+Z�[�L)n�n���ھ��ƣj�������Zc�x�wn1�#G�Fkq��C�!lF~쁵�, c�w�Qh��M��ֳ��C�[<m�>���V�֚�JAQ�� �-8�m�`tf��W���%/N�,�����t�A�����b� �כ�C�he���bûni&B�մ�Ym�<��?!��?��3�i'� ``5~q�Z�.�)RzUE�ՕS�����h�j��G���U��}v�w.�&�EW���N���Mz�יR�ş������u�/����dq^�*�htI���D=�ͼ��=Ϟ9�3?�2�#ן5�O�+zRC�����!+�ʘ76�kZ1"�x�V,S�ZF$
��F���P�Q&9�b=xp��c)�c+ #0᛼�y=��-]�����9QN^�R(��Q���ȉ'b�Y������Z{��*�Z�Emn�Ϛ��a�D���b�L�iM�D�|�{��?O-%3@^G���ך;	��.D��,��+����}�����:��h�{�~�w^PO<�YG�$�p��X9r[�%��
�%�����+L c��<D �S�Że�cB]8�לp=�)����Tn�ڋ�'HvA[(,Ù���/D��g�r��5�hw���$!(u8%�V�g�[�ck��%E`��J��ii���ǈq奦��{�ҳ�ڵ��k4�{u6�ި��9�v�*�h7&�1��9��KJBA��^=���Ӎ��]��^��&���Up�Mr��lGP����F<o���t��R�j��ee�%q,�bήZnB�`��5����Û�Mi	� ?2T��@�S︇��d���*�k9��Q�ݎ�Ÿ��F�s��)�i �\�Q�Ah�i����
7�
t q〯�OW?��ՀX�B�n>|@����ă"����������)�	��pן:}����dk�7r_�	�C�<CN	�L>�H�%���8�:�͙�s<d��h��J�? �Za؆^1m1(������"�p���Y�V9QJ�nַic�� �U̵u����|���p���z�{0w�i?o�7��l	��?�3^�Ñ����!{w�X�]ۓ]mi����I�V��v��) ���h��G��+5���� �����	ެӱ��h��{�y*+j����H7͸_%o4+<�f�����^�ɪ���N�<�4�#���h�y�N����6`�����>ηZ���X�������0�yB�.B���[ӈ�8�zj�x�ҙ*䑂�`^ kUx^��[Ψ�)��نw�6�18�Wwꭇ�ݴ�l$➳W��Y�P7�9BGT�*���Uq��ȂNp�w��Zv@�/�����0o�}&�Zz�?�,��`@$���g;Z���Hε���\��ZX�S�c�������"��ݞ�{g/��n�o?��mi�Z�<�Xχ�ܿ������ 0W�F���
�D�u�%Yg@�C���i�ﻕ�h��6�6��ЄS�t�D��;+4P���}�ݏ�)�8��.
��\��gH�i��~0�)�Βs���t`m��"׮]s�G��h�]��?�=���z��{8�x!�ԓ_A��R�7?z�'xv%N�����@iԚ��n%���@xC+��m�j�V �w�:|��;{�9uw������U�$�9;�����g2���܅��7��`G� �g;艽�y�d.�wН� z��ʣ�#�2����J�-֎��3�Ȼ���hE��5L��}�Ղ�4�Pp�+�ބ�\ݷB/襠�B�:gZH���I4T�R�AA6ơH�j7��T,�����}�fY�ƺ���V�.-/h����h�з� ��7�%G
k�t�$1'��Ϸ#�tU��S��m���@�c*�sCh{�Z���������ΗU�d�j ��P�˚y�ڀ~޽��.��^k����wg���%,:���b���M���7�z����S�?נ�V�O~)�O�n�ː������5�c4��|#��-)�&�����qf9�i�9��P'rw��ƿ���x�7�7��C�fg�6q�x���	�T��Ξ)�7]������\pD���������@��*[�F�u��e�ɼ`��v���^�,�)�?�����}%�˸6K�(��'H�u��A
��ɌG��ڕ�$-ڔ5�{��L�'�t�"��믿v���`ԍ�l��%��@�h`��[��f:d���]��2�wܳ�g����?t��;;U2��}���s����)���v���c�Q�Y��AOXf8�u�C��P����g󼺥I�Y�&~�� o H~�ɧ̏E.8>�bM|�E�ХK��#�o&T�q�(�����A���Dx#�[@y;>�TDK@	'VP��й�e#��5p�Y�މ�4������Ѣp����4;�z � ���h��y��P��
���@�onm�����7X�[7�E��B�+�.��[w`�#RwyV�w�y�c�|^at�z<�Sč����6�S�p��`Vy��M���������ځU�X�x�����$�?v�]�.�����;�9 ���>&~�� �9cާ���I��  ��IDATvؐP=,$��@��	�Vt�Ν�� D�T�����8>L�m������ۆ,��-��i�s�6l,T��7����O��D��T�H�Fka��P�.H�t����7�y�=�iju<�� hƲ���N;��-DA�c�I�sU�pQ古uXj�Iq�~����tǷ�A(y1��ǘa��9}�EU#yi;+��֊�U�(���u���� ���l+�����x�Z�w���*�[<e=Ϳ62���u!M�â��&���QQ�#���4NH�a�+{y��W��z��5m�}��ٲf��J�n
K��U1���ا��Û{D$r�L����~�1��/(zx���gGYW�<3�BAV��-�D�nH{�R���b� @�`x�W�F�u��e-��u͒"����Jy -�6m��^�*+ڵz�ѳ�"AT #�c�G ���{�;i��`��m�r#�s;Ί��6����5���n�٫�>gN1C�r(btAA�|e��z�`8���D�\���,�>  ���(�Q�|��Yv�D^g��I��5���ҽ[7���e!�e����~��[�XS�������V��/9%�&s<OϏ��Y \�������+����g ���4� �]���ܐ���6'LhR{�d]�|��#��w����A�("�W�\ak�1#'�Ԣ]�D��-ƠQ����i{/�{9S��}�Ɩ��w+Ӗ�p��l1x7~��w�7U쳷�">䨯9~7��G���C:��Յ��|��F��E��0�ĵ(A[�R/�<�L�7��"�n��\���UP3T�5�\�fk��w>� �Qz��C6�ߓ�m�5���_����>���� G"���>6��c��X��:~��L��[{�g�8H
�*�]�9z��}O�=�C,&�c���;(¿�%���8\�]t��$��Nnr�H�d>j����#v�ţ�t4ϳ3G��L���p@,���#�!U�2Ǽ!���cօ�Սh�����Xv�ve�;w��⡍���O�?����^��8<�_^������n"8'y�&l�t�tԁ5��q���Dr:՗%��Ku%*Va�@�ؔ���y�%	������X��r��an(<����D�~76���������
	�޷�pYzT�y^J�Su4�;H�|J��� �?��c���5�`rr�6�ϸa<H��� �xEAf~��tH���)����[��k���_	�ۧ�\��.�'_X�|b�B��؜/t�̛a�����=��9�8ŸK�վV�}K����4�ڨ���T/���Á �BG��f0XL ��u+y��y�!�����zL� �%P6o�}ߔ�D ���>"x<���D�f�b^U�@Jh>��7�&��Z[PBaAi���*}`���P�<�Q@�ps��J�W�e5x/��pCq@����f��=`3.�P|`�%����u�'�ǯ�k�31Z�gB�xx0������á�w��ӣ'{
<��d{8�����[�����@��?�W��_��mD��°�w�^ZKb���{�E����M��R�B5�}e�'.9:d����_����D�H������ (Wx~��awWZǻ t>��S��U?��S��H�*`�c�n��{��� ��[3�Nՙ��(]��ȇ�h}����p"uM譄��2����>�~�*��n����햎u�(�Nѡ���O��	<��i?�cc��uv�4&�����Eq���a�{%�oD�#��WW��gUb�y�`�1�����^[nt3Q��CG�.��S�IzO��&Gvvvҿ���-�t����z�X|*ea�c�����7���q'O.���nj��5{`�ap�ъ��-��#��W_
�d�jTp����x��ԩNqY�M;WR�ZH'D�u#��1"��Hð"������َ��=E��f�E�*2]�`r��9
����q95 +IK9q�� ��s�s/I��Q]z�m�#��9�Z��km��#ړ�!�cg�	[���&�H"��l_Gܱ�x��絵���0��g��>)��I�RC����SR���`�(_�i�/�2��.z2�1��\��/��̳�/o�7�,C	c\! 2g�Cv�����/���}�uT$;�\A�!�*�AB�SFC^h=����Ҫ����i�Ƚt��{�bN��](,��k^$����]rā�J,>+��}s��>��7(��U9nD\{amh\�s5�g�	ٜ:y�������Ç��&mV��
#�㍁� M�9��>�-(h@ ���!!0&��6���:{C\y���ˠr'����J���V� @E'��S/�0�@/. A�dPQ@A�ua_��!�L��Uj�`�k�KnZ>��@�NaO�2!�;�+���K�]���G4�p�m���1E��U*eX�XS���]+4��������.\8O�҈~��_Fpw��ƻK��&�Dc|��#�0���!ʹJꑙ� �ٮŨ�co�����=�-�
���O�Ӌ�p :}�t�Ix�]J�� � _E�Cь"��<*�������w��^�@�������F���a����w�]��9�t��^�i��p���ϝ=���V����+T����h@��g����my���ч��Y��4�j�4^�cm���7�q0��)�@���E�ߘB�wO��Ѯ�9g0H5 B���k������c�4��������՗�^6`[ J�?d-�R�V�C{�w���F	hx=F�'�t̸�~���;9b�,��0�D�O���f��eN���� {{�����A��c�u�N�5�䑏ss�}�[ϻ���O��xF��{�{hF(d;:����;`�A.�=�(ΚF�~�w��i}��m�]k�m�dj �.̛5��}�r&�A�yW9k��ÑxY{*��q4�pF9�27Հ�P7v�w���F�a���D�b6)ˠK:B�y��	�	X`<�鑛�r	�N-��ǜ�v�W8c-hS�o�����<o�����������NNg�1Yhť`��.��bm1�ϟ�]���8^z���+#,��9�eS!�1��]����D��#���iU׌��<�vRV��s�8�}���4����H9�z3���d�	���N�{a���'l�遨:��S��ŵ�(C�::H] �Ap� ~�� ����؉��Fr��]w?Zz�I`B=\�8���f���E�|��#�W|]�.��
�mۦ���[��r)�[>��[�[Z��e$8�ҥ��ŋ���̃�m%�j��9,[Z��FA�X���`n�{�U;�-;���c����A�� L�j����~���Z9<m�^��O	���q_?�x��n`^r_�=W�:e%&�{8�Qg��x�E���kki'�LxW�*�<����W�J~y]������}��U<��Y�-(�0�\p�j9�e(��}�{t� �����>~�[����}�~�}Kb�f4���*|���z�����k캇=x4*ܗ^z�)?8�1�/�8)]o� G�x6wS��O(N
m/|���~ӈ! m����Bx��3�Ύ�?���w{�6�{��3���<?v���Gr��<���YU�R1���!��7f;J�u�ϟ���	���y�C<Cwݝh�&�y��ؒ �n�z�����^d�[�kx_���}*���*�1��H����ӑse�Ty�쓺�4���(�]����(qK���)��X�WV��5��@��Z��h��o��������y8�"�g��R`L��i����U4��&��v�)�l=�S�MD꼥�,xW�W$z����X���bs�� ��i��3�d��YN4o��cV�����8?k�9ѐ��nf�}���R ��iP�'�a�]R|���Tb/�ߏ�hG�3���@Cp���ɧ���׿�߿�6��Z,o5%��'�-�4�ǳN���/��J��R@���@��Q<׍�]�G)�4VO�퍔��l�_X(D�5:R�����;C�-.-p�10�ֵ�(O0�� ��ڲ�Es�>�r�v^F���l�v���u���?������v�$�����>��O���|�)ʤ��N�(���]���9���BDC:��)�I�\��j��4y��.�G���3��i�.P�c[Zu��_d������W*pX�f��팤j��K�үeT�.�|ή	F+����l�&��LEռr�����(����=s|/=�����]ӹ�H�vR��R����D�eE�VY��3�f�xP�a�U�d�vMV���a��,�ϨJo�8��;�.-�X[�Z�����!�
]�P���ޚ�?#����w Ӯ��3��[)��>)�>��[��|��B��13J4xR���ċ֜Pp♽ހ!ɉ-+��Roy,��cѽ�6`���'�d�d��A���|n�������²��j+�G]P� �?�я�VY�һ�;!mf���������w�~�)��o�����!f�1� �s�?O�n�M7 ���s�=y�J��ƺ���kZ�x������潻����A~�W���[�u�O��^�o?~̽��klu������9�J ��;3Ҧ$��<�-@���Q�@���� ��f��Btss���%>�^]��~z���֭;&b�W�O,����L�YZ~��0�E$�|�B��I�9��.�q���Ï>L���kM�J�̓�]��2��9�y� �m�/,-�?�`4xH7A�D�a8�h���E�!@w��=��>H���xw�a���q_ɗ[��s���U��3+tJ��%�,�-�
�Am�K#��=�;����:�	)�^��V��ܝ��ZQ[y�>wt�eu��T94���-�� ���!�'|G��4m��c�b�� ����@��U�|$�k�,��^�?�r�^���� ����>�����o���{뷿���-F9j=,�{V�2��������,y=�ѓJR���ַ^�̸��W�V�^7 T�(�ek�x_��-����B��fH��o{��s.=�f�7���{��E�{1��a- ��������.]�Ĉ��5���N?��Sn_�S�b��e�=7�de9^�r��#����k�%���Xqv����o�9��Rza3C�M��DtC����p�E���|x��=��R$��7��7w�;w��H��*�U���(x=릧�Ҋ�,E�Z!RA��"����Pgk�u�q�|`mJ�^R�E��1jR���4֏�ش� �!wD4��x�1�9�2!xnJ�DW�s��e� Ó�,��Q��W��YY��6��j���42FYLvш���m��ey�.�-�y��7�3�^ؔ���v`ū"�Ӷr�d�A������������F#�Y�;�����*=�f<t�&yϒ=rHevf�T�{c�z{�5ݭ"�g:����'����琭�C�-xK�,��EP�x�h2V�XNe6��7֪����˼u���ڎ��zfw��%ybE��5@�(����Y��1�!�,��՜�Z� ��0N��B� ��s܂Y�����{у]�YDXA�C��@Aw�s�v�w�>��
a: BS�2�N'�{��y��3�{��1����;y4�y��IC'<�~��FΨ�N7�o���}ڋ���=d�C�FC'��~Z���! ���`uu��H��wsii@E�|w��(ü� �'�n�x����t�H�̱�y�8-w�<Wx�zker��a!�S�>��K����U)*��e�>DW��q�[^Y������2rh�p3֣I����g�tR.'zڏ&��4Z�C�����s�$�	Ғ���,�"tb�|ǽr��i�v5D����o��ot!e�Y���E�4�B3%k��k����G4�g�% ~�����s�����	-۟��,/~�E�ʪS���\�x�N�dmW����:y������~�۷�f�4�m���(�0 ߨJG��H�Z@�@�1��Nbt�B��zܧ��x�G�B�朾`DC�B>�L��lQ"�9bƾ����_H-��q���E�՝8H[�$��һovDF(�$]��Paa.qf�F�,�Ź�No�[;�T���E�r�g��H+���_G�4���vv�v ���]�&�qT�(7K���A��jp���8��)y5��+��I�Hw�n޺�>��:L��5-F�G�6Қ��Ǫh$c�`����Ǚ�4�ポ����Q��WM��w�2��
�sRO��,?����c����tU�)'�� YdjIz`.��f6
�j�ZJ �����(�_���ą[ٷ����鸹�|9H�U�M��O�k�8L���	���.v�J��5���\��6me� �Ӵ�Ҏ�	dۂ�΀��2�mIŉ��8Z���|��T������J�bMZ`�|�lAV���i2���8ajH5�6F�KÐ5��R�Q���)�F�
2��Ԍ.�^	n��1N�dgp3W~�\9l���` }��m��[�^��8��0Z��#�5�
	�7 V%]3G��u2�%"�u�Q���^b�����=|�;u򤼑
g�uidJXlue�I��q�8�
�cMj�M[�/�� ��J���z���3ǢD6�\ B{Q��q��<�_G]�rC�-*I]��>i�(�&��;z�)<���OCP�ǋ5A0�,3<=`�ۘ�m{>��p�|M��� p-G (�/(�74��u1� { �s�z�O��fe_�����LcM}]X�.���@�Y��,����	C��7��i>�QJ� ?4�{nn�;O
4�*�
ˉ�t�Z����h�:�) g�3y��y���J��]��#_�<����{1L�
h���yIy��.6����/M�
*é9�gp�$-���o�;ơhw3�^x�1�7�cF�Fb���lJ��{���/>ǽPu��s�{�sM�y��+︷���J���6�9;z�sJ���ca�H�
�Y�;Ʌ�'�}��m~a�M���/3R��o˼i+�������O�==��[o1�L��k�Ҽ�v��o�7��h�9���j^�D�'�1��_��*�+0�24�05R���*4���0�~�Ę��>�մN����SPk�)A=�ޤ�#�pe�p�l)rE.��׎[]�a��
�`{C�Ȩe@�\�Uԉт���*� qCeH�tMf�����=�>c���;ƚ���\�U vشN{�\�9��1��b:��5}3��Z���o���
Ӥ%��s�9mi�Bg��]Qp����p�T>�zax�4�ڢN��Qg�w��v���922�0�v������R?y������s5�Mi����gx����S�uz�E7Hz�m%���ר�BP�Gs����s�b�"wB��,Y��;�����=�]����Z���2;��$%��Wfx!<:l��`�yl�ͧKx��2%�G�R�"�wP�4�C~ZЍ����.x ҼB߹�'�Ķ���8(Z<`��$RWm�GZ�fҤ%x��D�!rS�����{p�O4�J&%3���I��h�]�h6�D��ʧZ;�L�գc����bǨ�����5�&T�>��-���2�� �C,�ڗ@����u�ƻ�G��R�r��x	�5�x<l ���K��9M��z2��9_�}�ǉ�
v(<�3���j��L�'z������3��{5��}�#��G/[׍K�[ε��M��G�h�0OV0w�G7 \4����<�z��r��P<�� *�NcS�!J�4��zHd��AzѨ�v�o��5*$�U��~@��m����������<4��66%ȕp�������3�(�XUڮ5�Zp���n:���x�*JVx�����Ϻ�_}���_���^ =���&���J s��D���
.:�QK>A�*��[�p���*�`x� �W_uo���^��x�g��wP�MI���F򩓌�"��0`$����CF.�u�@^f�ԙP	 ��'��x�&�xr �V ��Q +D����=��4T�c�|�?���
��9�"Y�<q��ۿ�[F�`�c���� O<|��]K�1���z!^[����Q��Chi�F��|#�s_<��nO��:���E5=簡�F���#/��L�K��h�/J���nǨS��	��� ���J8�k�4��a!&��97Q�ܮzz��"��<���(�:F;�$�e�����Ekj\T�DΚ>�)p�C5P�_TG�EZR����=��4W�Q=���Q6�JQ��Թ�=��s��t^Mn�1`�"�_�(�i���&�Y`�'bc0������D����5K	y2(���+��J���w	��U3� �V闫��u9�u�7��rwq��6�5�M�@v\�!���
�����z��gan�u>��	n���Z.9�q�j~Kև2��J����쳷wg�����1OcR|�Gi_����\�ww��E3(@t�}JC%�G�u�/3gq�J ;�6��M��M�bCm[��TLw�4�~]C����KOQ�t���?'��6��2�������V'��(h>��3��}6](!���aG ����ŋ��%��c_�e@��%�Q�Hͫ�f��l��Ub/Gp �K�˛��y9��Ix�������(�P̉s^Y`�գ�0X��M�{Q`Kt�gE����Eh�e�x7%_���y�_E𱾎��]�!B�w'
]��q�{F}%��p�^���mB�ٯ~�+�U[Yf�6��ݼ�7Pi���A/4O[�[rO�-���j霪!�?�����WsU�_Z�'�D��#��N�ݲ��+lY�w��a�. X�����;�v����PZ<R/.�aZ�ZGH��u����& @�7N^�50���k����� �{�9��8��{��7�e��J�����[�Sg�B���ZF�w��9R���w�g���CX^��sk�8��60��zܧ�HqX���ܽw�E޸r��� �����ܯ_E�
����X9��������� �s��_ჯ>�s	ü�[�a��aL7D�pL]���9|حX�Ȍ��ƕ钦_�q��MY8���'F�9>lիV
�_�b�����!Ly{����K+M!�1PK�I5i4�'����e�Է����0�9;k-CR?_�t�̓T��C�?���Ȇ��!Kϲ�#���P�2~��|Z��E��K�׳^����W��#��F��$�o����I:�����q��(�]��B�����Y��K\�,/&<Z��K>R����N.�ӽmq�^���^aCG���o��νu7��1$T�1�=��p���A��Q�`��S�
�Q����˖�t�. �S|��\�+yWhB�����5*�;�ޫ���QW�BV,w�3N<����~�Y�����C����V1�s��?��i`�֜��w��WY�z�P`%(�k�Cj�_�T�j}�,YxU>��#*V�}�B\��C	#�O��_�L'9�`W���X�1Hn�������6��0���O�D9j��2O�+�.��_~��ZHgXТ/�؅�<ax�������y��SI#+]�2��{���o���1
�61^(�F�f-dJ�RH*L�4����a2H<��a_���/�3ľ�`!w]��f�y��q�k`U�M���y����q������Txȩt�r�P���������\�.���_�3���u�nCPH��njā��kvz��Xh�ͼ.�9��r/c�����u&���h̠s
���KO� �e"����λg�}���i{^ܿ�0qW��[����V���Ȃ1V���S(-7[�2#�F#�h�� �(�D�<�dl�x�A:j�l)֨D�ĥS�#�G�uO?��{���l������Qc�7R\�K�(MKv5W��G�|��7�C�K#�^f����W�
��h�{�;E��4�g��6���O�|��/�����y�i�0�sG�R�Xp�:��H����|�4X�s^"h^�*�,��ߚ���٫�@�J@ht�U4 ���� �j�&����(t{UL��3�q�q#�e�ǧ�2רwc�P>X	���Z��юte�9�
ĔI�V�3��� (F%W�}�u f:��;��9�YGy#��\@�����8g,��+]�Xt/�bu���E����T��R��)>�s�����)�r�3,,�Mr�v�J<�|�=��_��^��jE�����2�얀W(*����ઔ7�dyN6��h�2DR��Cz0�u�1Fŀ���>� �+_n��{� ����!?o��tP�� ���N��=?���M�ׅG�7pc�Q���q'>c1�ԣ;]$񨭐=��[^�97���6A��mҋ��Ca\W�#����♽��R�)��}慢8�[1����o�g+I_���ia���� ���p����B��˺���]kK)Ei�(I+x�AyǴ(Y�]	���}�:tXs!�և��������!h(Yx]�O�����S�+������T~G�)��r�]�j�X��g���7�']+\���H���/�?C49�oiG+l%��7syi�ޞf"�����wa�WX !B�0n߸��#%�Y*K}s�	��ƾ��c-��ձ���{*l�<�V/����͛��/�t#���۷�{�O0�5�EN�+�H0��\Y?rc�Gs�� ����W^ɣ��!@�߂R�a�z��GwWOaG_���<���$�����a��y6��g� tM�x��&
��3D�@PߏF!������B��B�=�@/�K��;@��uD:���*E���3����{*ݘ2�'W��+u���?.�n���1�1<�����w��7opK.jq�Ԕ�hɎ5C���x��"����4��<ρA���gׯs�{�
�;jş#��^�S�D���3g	t1>�	xx�ͳ��4�4ǒ�T9a!�&H��==m\�#L�o%3E8�0��+����iZ ��@��>O:U"�_���oT�⁷��^͠���bH�(�ce�W|��ۤ�i�Ѣe<R�Q�E��/m{�e�[����(��S�@�|���~�������ZiެyI����nta�*�!�l�F5��EM���t��.��������ִ���z#��q7̠�������������g��]ӑ#G��X�uq������R����Rf���rv����e^X*:��*�F�4��ӻAa�8�!�ڦ���i����y��@���H:3��(<� ��1����\�<��U�h��<�Z^�pF��إ��}4HB�A��$�Ժ�sj
x��KXk>�%,ؙ�����`�ò�{M	�������ܞ�)�[��������a��G�i|��.�H�TbkS����9x� a~E=��w��(<+��w~�pw���A�w0�S)!�JS��圽:�Cq�~��U>�XR������f�K
/�@�Z8?ӮuR��^���^8�x��<�LPQ�3�=�jS���E��	x!�IU��k��V`9�0Z�V��� O��Q�d�e������d�<�A���\PL����S]���}��͉���t#��=�1X�P�I8�
�}�Y;�Ȑ����2{4I�����Rbެ���ߚS�`/���V��^ K(�&9MbޕS�D���0Z?4$ٯy����)��R�[l����/ݑ8'��5����ª��H't��I|)����}����<`��QSO�7��M�[�v��Z�w�]�rsI<��Γǿc��;ȉ_^r�/^R�]�rg�h�o:f� �9*�v���3HE�c�#)��p���~�}ad�]2�n`�?����?�)���o��~�����l���w�C�9�{!����� H��h\�m!���i��~'h�9��]Z�ϴ+x3z��*�vbx���Ƽ�i�l�G�<͘y����f���3�>�i|zN�;p=2m�:߭���x��e��.,�3��c�|��>�!?ѵ��>��fT�6�J5��1�K(e�X�V{-���Qt�+4Q�R�W���x������ؙl��T�ش.ǲ�7�ݕw��r�P!N:0$�O��ʖ�tX�Jv{(�����y&���X¹=)���}��mM�K����̶�j�v������I�3�3Uv�[�A��͔�P
K焕갼H	3P���*��>Q�)���P�B�ǉ Z�}iC`�1G>[s	�}�e�u%h�9�g<���3��[ұ���b7��X�n�/��i.�U�P�1:�� x���j!Y���l(B����s.���\�����֦����$gG�;����z�Rc7N���vv���{wI�\��*�����my%�^k �0 H����B���։Nrм�<x䞢���>��o�a����+�c�޷��vg�H�<�KQ/-,��f�Dl��`:>�v��G��|�)�<��� �G����B��sȽ Pv��¨�v��{F����8���I����QN	o(�7�F�ab .��k_~Ir(�4C�(�YH�Z� �kP
� )0�����Ώ\(�Q ��uhe��W
��j�#�;��w����� �-�]8!Ȝ�]j�Aڧf���p�����#hQ���sT�V����&�Ԧ\���_�׎	S~�X��,G���c�O0���u���IH�ܴ
z0��3gN�G����gJ�V<K��;��U�c�+��!>�^b�;�B���L\�/��w⦺���o�y�s��?� ��姞�
�I2UqG*���3����3��o���|����B��u�Ե�_�l������)��d[qtn]����+��O+��9���:������nܺI��۷n���b��3�/\ 㒳��܉K���/�3����f�(�b,�k4��3��r{g[���h��Ӂ�S*�O�z��@�Db��=����&�[w�ѧrTr��ߕ5b�����N|�X�Q���x��H��6
�M�T�Y7 !�s�HC��*=�3HRK��JڡR�Dh�3?���so4qLi�Bg5�J�[�{ZMHPd��wو�����f/,Mqht�>$�T�'�S�	sN����
.	,	�XaOXTH����6�t(j��A�b�)���H��6Y�<�����4JC0>� �=2���=5y�@�
�Ѩf����?sG�eW���ɇa8^'+5<� i�����fHJ#5�T [�����b��O��6y��VK���k-&p.���φq,��r4 
^��E*���}�j:�"����27���I���.d�n�����%"� Ӌ��z��	�E!�ˀׄ� Z�䨃��6R���1�VqW������hhnP���C�XuZ�ҍ�)�W5�0��̕�MB{�a;q]v�g�)���
^x� P@�3T�YU�E�:��Ĩ�e�#��ta���˚+��׼��-�S6SpB*^8�謲�H�Z-RqY~��Ϙ?E��8Xtǎs�Ϝa!	<=��)[�2�Q߹˴0�Ƅ} �g�޿���}�z�4�u�8�l9�R�9X�@��Ó��6������0� ��
+�I��/�u�gQ����0�}���5cV����<�	��"N���s#�ً?�g^ܵ5w��9ޟ��(P�BJ���G1�#�*��s<W�
�*K��L�ä���b�'�2}W6|q$r#ʬ�Z��w��׼�m.P��iYw�v.��8KF��7H�_U��J������\�>|��
>b�5�9�s\?��C��_��d>wk�������O"��1��y+�%���ó�cpc��bs���G�1�;- �"�����}�O?�ԍ�K� �䳥��!G|�"N�¡�0�llK~g�T� ,<��.��s�>�z�{����K�{��<�;������A{��E�O�ύ��б�&�Q� �[�.�I��:%)�̘��MF ����Iz}S-�������;ܛ����f.���~��q�+H�׭4gX���Xy�+�z�'Q0guINGdM�N	������p]�Ԓ��3��$#�	 �{YK�M�ؿv���kKv�S�(�{<�o�V�W%\�F�/�7���+�׸S��!��n�Fm���������S��0�O�"x�?�t�A���՗��� �a,�n.�Ӝ��:!�i��g7mH�\�(K���U�C�6Ë/~�T<y�����0�T�f(|��|������q�y�n��0@�QSq��}��P��Zu��]������ǋ	�X.�j�y�^��7#��u��'��6s��Mt��J�Z�s��X�"o�ܩ���RG�}���}��
���4�M�y9�>yЌ��Gq�x|G粣��ǣ�P�����)�r^g?㊟���ط�,��vv��A��P9��<}u��� �(�O�Kً���a^`(���S<�X�3?�}}��	*���� �.]�D`/�5�=߀t�"}�R�	UR�^����Ɨ���c��P����(�"�|Ң1|@����"m ����h�\߱	��g�^LF�c�k��<'���-���莟8�E�Y�7��m��=����/��
���{�1��ȅ���
e,lM^Ӝd�1H#{���"��O��K�rQ\6g��Atk��d"_ 4L��KNxO����6M���e���mU�*-@��j+��*�g��\�P�(���`$��m�`7� 3G���~�>x�5�u��2��zC�t�Dcdue�<t�i L� U#�n���>s�ʜHZ	�'R�P�()�<w���@b���`���x��*-�3�0�s��	��o���;��;w�<�u�cG���e�=�#��/k!~�;���N�ԓ�S����k�̮��m*���+c #�{j�H#�F�����,jZ_�"�Jh4e]-`e��Z�G{��xK;�z�/-hH���'44�F�ceQ���: �]g|�ֆ�����k��O�#��o��e4"�ƻ����(S���1�dE�X��4ԩz/n�=�:}!Z��46������%�E�MX����9޶=x`�����|G��=��Cc߲F!���癠����'�r�4�)Pk]{�l����ޕ�f�����nnl��Ơ�y����M}�/�D�G����lus¨f%ꭃNr��o��B<���杚ڍ��V��H��Ki�jw��.+���*A3��t2V	6μ��,2x
R�o�����Ϝؠ ��V���D���%X=����15bsc�jdRؑ֨�L<���h+V��~|'����?����Đ�7����������ء�0(͞x8�ݝ�$�^2�,-cR�\���?F����j�d�s�9@Ƃ1��(C��~��r}�!C�!�'r�E/�*~��n^����6<���xxS�=�ݫ�����_BkdtN�W��x"�.B�����#.�'���F6�y���
tN���=ݮFk�&H{@�$�@���~�'�;��r��5���j4�������ur�"��$�=�����u��T�`�P����ԟzY�¼�{y�����g�@+3�.�D�m.�/�m>��Hx������KZ�Kk�qR4��c�਼&E�@kΪ�3OF��Sml%쨄Y��ö�Y�f�4�ŉwg��!�%
�����hW��0,,��	<+��������O	@��������#�wA�5H\Ǐu+��w/]d�W��M��}��5��dցki����)0�d�K2qvo��}��	���[7	v!/]z��h�9��4t�ZsU��6�QgUb�x�[>����R-
����"����6��}�9k#�sx�/^��3����s�f|�0>�v����.���
�jsَ��;�|�����0V�E���x2�0Z��5Lо_iPt� �
b{�q⪎K)�8�X�/M��_b_R���_(ݺ ;�vC�`�S�*������96fwUb�TM���x���<�F�Vj��ƔbQ�)��D`׶���o[�^C�D�ذ�t�
ơ�#�q3��MP��%�V���ˆ-e���,l�/�&DM%Tp�'��PNX����dʥgת�-��
Rv��Ҍ��o�Zq�2��[�M<v6RŁ�ε��rżPRe,�� O��j�:%ac��8�Ss�����i\���.n�q�줬Ґ���Q",��<�C:�����Y9m�A>LT��g�7^C��s�P��ok�e��]\�Kh!nx:�_GiZ��a��z�\L<M	��A)�*�/�*
�Xf'���O���x/
�[�os���{�o˞1 �E�+�b�s)Ғ�:�����x��J�>stq��]_��!?�\�]� ����絵�i��9�t�z����eSt�	؁�R�<��&3���ȼ�3`�F����Y����J|V�
j�ݪ��{�{w�Z/3Z�"�Wu���b��y7��|�;ǜxMg���K��:�G|�g��e]�� #@ܿ�2d��b K���������~s�?;?u�k�S�ӹG ͬxˈa�f���YgRi*\��;}+�Z4���=�#|z�^�F��c�����A~3"��H=��Z�Q .�w�H��̫4|��"xu�~�m[�]�`�hN�;�kk���ۋ���5i�c��&"����=W���nh�=���}=�{>�� t�.�]6�1:�⠟7��\ Y%0�]6����r�߇,����'W�������wW�y7��'�S�~��s��#���4U	l��)���&8��x6�"����.
�"u��9�8F�ci\!u��3RF���=�g澬]G�D$�KO6�a$-"ޯ�IN:)mh�M���9��v�Lt�5�������,$p+��s%�Ņ��x2���8��`�A����r�
@���CfВ|a�[����#�����A�sSxZZiz�9��cGO�������B�����5_m�����(3��k) k6�14crbC�wSQ�1$�w��ɕ��v�SJ�W�P޿�l��]��1a\<	 n#���h}ܔB�Çܙ�g���
;�Yx����9�u+o�����z��z�
�R�Q�_(=4�IĠ�B����x2�*Z��	��W��N�w�ң�C^�׋.x�O�ܠg��(h�� �3�ݺF�z��r����b/Pg9_�V�yM�@�V����mUj�Z��\10ܹ�q���L�X֦6�j�COi�Z��=R{K7A�?����պ�YQ�K������te�!�!��O���>��@�����������罂��pW+��g��������4Н��<��wx��A�,��Y���S�3ny�f�[72��P�d}�u��[�=J:$��Q����t��슠��}ʅM���w�f�	k>���&(t�r��@t���L��(��w�W<�2�=wěѯ�hl@�4
�j�T��P��]fЧ�!3/$�Ԓ�����h���ʕ��I��qAY��	��;�Fb��M���1^��E���y7��� s^�0���3m�wR�Z�o�#��%��������X\���W̳t��x�8w�,�	�# KZ�c����Ҡ�.����+;Uz�ڄ�Cs0���7���0N K�+
���b���6�X�����������I̡�/�)�vӼ�\�`r	m�Q7a�D?��P�B���S'N�}�n�.��W�a5�B�UDJmN:�����h�.;�hڂ&�������]���\ੇ<��0��<�������K;�:�4�,J�[�BS��ϸ��G���B�'N���S�+2O�[�=./�e��]����N�mT.��H!�`�f2�)��~2)�w��d,]���U�#�ބ�Ν7��໱]u?�-z���� ������w2Qс-7�s��.vA��P���as�	��o��.�s�MBi�ps]���Ξ=�;��E;�W�Ro���Ԏg��T3:� ���C�&���#b�`Qܽ{�$�_^���(�@*���R�(,"L���$5��5�P�єX�Ԏzu�..��=��>޺}�t@W�^�����w��^|�����X��7�$`N�b\�cd�X�4�a��\A��_�K]��`�d���C
0/<w/��{!
�S��o��Ujc,p��̣���DG-��T���N��������޾u���=p���a�1W��4oY{��u=��*򶧈��I��]�P�� ��� ܐ� x>*�'o�F���7nѰ3~J�ZW)��<s9��h��?�<�3�y�g->y�Z����H{K�8<�+����"�^�G��T�}�r�=�=)꘾�O���is�bQ��2d�x��W�{�P���/{���O=M�nъ7o�cǎӫ�Q#�����A8f�To��Ф\PS�ӓ��p��8|X�%��`���9��	20h�-�!��ۈ�G �1���_��1��c��j�W�7<Lׯ�E0��i�T�zܫ�ʪ�\BK��i�)J���t�g�B}	����*^�.�T�vM���ѐ@�o���L'�
��ҍ҂���إӒ���E�㛰��˗��ӧ�����Kc<�����Ґp�����"��öaj�B�L�fmQ9v8,��T�ǡ
'��<�H��������A	��=�DFH���'?������5��b+� D� �b�P�����ێ?KM
�K�6���"U�������	K�<� �0�qƠ��`AC��!��w�t	�.d��(�έ4J��"Z�s�����[@:�݅A�V�Oq��7��PVƣa�����J�7���!���E}�!�V���O?��}����\���!0����?\�C\��s���_�X�c���X��,��-�<։�Jg[Q�\��*�\��рx���t ��*:�ͭ�e�KI4܌9�_�`>!K����mK3 '�I���0�W�B���7��K:���32'�V�CN��Nb�(�t��F�<�"�R��7q��k�'��^r��P��y�)�
^����M�o�]�\Nz�8x��>�͸oI��N�$!����|�65��	s�߰n���w���G(	`�����n�Cbi$�Si��%y�1��*<!�z]DX�Ԓ��.�������/�1��v<�f�� Y[xK���������ܿ�g��;ɸ�)�Y/��>�\��o����48>��S���"��P�t���P��8%�ѡ��,ؕ��L��j, <��㝶�^ww��g5&+�u�P��<��jf�y�=+{]��\�U��-�J�\1��R�$�k��}���1�j`�HcC�26�P�R��G�9��5K�1�0�KO�zi�A���斌�X�ϥWjz>����r�0~�03��kst8�3�:�☶�;��X��g����o���-\����_��?t� ��AE@P��*Uڂ6�V����������ѐ+�g� c�����p�<!��@+�Ԃkѐ���y�2�E#� �l�El�I�a� o��Zk�)a4K@APSo+��ң�?�e2�$E?�tq2TjT
e�So�xN��8�4�;��W)]!J8:�ܑ*ch��ЋK�>k
� �R��(�L(^���b��;��Ҩr��;E����VAxvkx1;"qD׺���Q!Z$��b��\��Ӝ=��,D
��^�X4��:>:���D��Nz9o?[���%K��N/��O�$�:@ư�y�,=N�1 ��uC�<^g�3�-g�t�X{r����V
;�I0����{R�}���N�۲O������렖=~�2��'92w��gk����5��&��MB����"�P/�Qc߃��9]��#����ی���
#�7o�匹�ԉS���'�7J����gD�j���|��.d�W�ၦFW�}�u�2v8?��œ*F�y�s�lv8T	C��LE�do�r1�z�:Z ���t*6P/{K�5U>3�T�%��3�Xp���Ȍ��9����f�Cr@M�r�^��I��6��.����18 �;q�@�-/����D�|���8L�O�r�LZ�b�����)/�����FBH %؈��&6���C���A�)�(�F��O�!��@ae���P`�:�TIȀSJ��W��E��Cv�3
����,����6�!��r��/��,��R�i����FC ���^�`7��~� 3~x;(�g�{N��!����]c�M6���VG���$0͡	��}<��H.���� ��c����	=�J�q�#p^���۴�5���Ok;��C�c�[
���@�R�sR��y�)hr�H)��W�I	�/:L���/|�f��c�B{���m�u�;�Ø{����2����{�pNŜS��w{x����}(�?�J���eFR�O�)'�������,��bLX?(�}K�̱�֍��
�ɆBE����'�óE�I�6����"�c�Iݟ�)= í9WU2��Kc[ ���u�^W��.�%ؚY��4�^Z+��j�N�������J'�v��(M��	x����5��ll�,~���"��6�m�Y�kjQ�]�Q�r,�IR)��X�ر�
�2�v�:��#eR�iHXY�B�k�M�S�E�u��D���ﲸ�s���Ӓ~,H�<<�(=��s{����������s���0?��
/��P&��s�d�[��z ����s�����qxu�1�9�H߱�� ����?�Y����\�G\����|��G��0n�4��g`9Ý�F���Y�H8��SG�8,bA�[e���Y����{?�?�?�����66j��ǟ� �x�޹���9\XXH�R ����ڤ� ^
�S�� �اB�)r�x�������t��p�Ѿ#��sm�`M�:���f��N=��s�z����Ǒ-�Um�` ސ0o	z+�R����~�u�ܽ����{��}kDI���(�"	Z�Ix�1�q�]U/ω�̬�`���J�`���*+3�Dĉq�8��Z�={.�>3g�R��h�f@�ޅ�F>(0ҹhQo���t�f�(�ظ�ػZ���WW[O����26��1�RK"�˽�xwn�q���۞�����Y�V�;d2��4�h^?'<��_x@�kU #-җ���UclU�/znav�{I��C���7����b�~��<߹S��qJ��H���q�Л��@�MpO��Ͽ�����;��ZECBQn���%�H�+���\K��QȔ OM`.�#mg���}{�;�>-�%���CD�H��P��kѤB��x�iD9�69U�H�-�	�� aӇg;���18� N�>�jq>öV�wV����5���a��-6��"3��!j n���"�q.��c�cc�G�y-��֒���y��"%�ߪ�I�
vْ���j�[7oС��cD�PNΉ/��f�%"3�$����P�W�
���EE< �+D���P

nD~qq,A�!��r[�����]�f<�Ec�<F<�?g�����5;�" 4|Ц?v������/:}�"��(d�mF5҈"��<�ӎW��j�������O�AFM"���v�  x~h��h�b#�ߗ��e�:u��Yز1pb�?�N�8�x��FM�Ѯ	��8`�>y�{��o1@G�U�+_��X�M��?�1������� 55F�Z�lM�l�:I@���`�����6�L�i(�T�9����k�����[~����D7hf�f�6~�l����W�Y@���ޞF;����7T�k���/ݯ~�+��'14�y63���c�`f^�K�qG�鼶��DhE���G����4�d�wÑ�x邿����߱�
���8Ygy3pݵ�s,��Xׯ]W`�͘�G�qF_ؿ/&���~J���lt<�"���c:�~6n��)is��K���+�0��X�Z�jI�7P^v�(-$P?��hk2iU͡���Н�^L�(EpvE
�t��I� 6q�pȮR�]&2���:Ӣ�� �2�cށĳe�e?f���t��`<Y�o�H�?W�k��Á����RՌ�~��C`48qn\�tUF�v����1Ȋ{,=�BP2I45~�wK����θK�.�yK��쐶@o:�7��@���;�PZ�b��)Y3	��ܢ�B=����~���E�%x�K���/��r�/����ر�TA��@?S�61�-Z�1Ѵ.��<!zOH� ������R{p��	�M��ŋH���n"�(>�Vc�m�p�dC��`�z�gyL�(���:��u������;���ss�\xo#�+	������R�[��V|c�O���,OW��l���dz�/<DF�mC�z^��z�� �9P���y�s���CLٯf'�1ι�eo?4-�p�f��W���?9W3���	��hZ�{z�mٺ%(��jiq�|Y�pZ`�)/����rŅ�S���bn���{E$���c4~h�`���vCM !�&漥Wk)��4�H�I0R�8'xܤ&�����v����4��x=>�k?id�,m"y6)�ù�3
�\�(P(�s⤅O�g�������S̫d�E�xd�P�ݼ'���b���TQIdG
ݴW)�h�w�^�$�]7Z�)�oI;�I�)y�8��x��w�����۹B�٥�[kidW6e)W��TT���](� �|@�	�@t�􎑅Hةv���W�gKt�s���D#]jR
|������.�c%Ay%�E���@Gm�� �EL�����^�o�gb�}����������F��m�����/~�~����ׄ% [l��$%j�(X_�)#�������
��Y�s� Z�]bOǞ&|�E�������V�t�2ڌ4�(�q!�Y�9�'��7�2 [.�p��jv#�g6d��q=��׭�������,>qPEv���2P��P�L�ҒP@���M�0Vl{փk ]�Ь���@�r&�Q����8#V`V���B�&���O�������Z��'5��7�)���5���[��nG$<���w�G� �"7�rpv����0���nk��7h�W�-o��b�"5�B�F�V���r39���~��%�=%�&���s��
��2K+(��.�z`i)Ny�J	a@p�m�Gѓ��zuF�#���2��S���[g���"���H�r��Gz��!4��	�T�xW�d�߽���#%��6�}���Z]U��DC���`3 p�6ǈ�����4%�� ��b�1e�(�q��%"e����Ä���c���X|��w~��Ɣ$n�qnV�Bou�T�9&�h�<bb�v�b�"���/cZ 5\����0,�j��Hō�lmX�j�}(u��Y�*P]t���(�S���/b�����Ad<v8hFQ0�����!<~�F�`¥ޱ���m|�`(�g ��M ]�@�i����r�P[&z�n����\�rE8�~��&j�i�{6�1����NW6���@�ڽ���n��4�.Y�);��m����h�)X\��'i
6��� ��A�ϭ�E�:�E<llq>�����?��d�I�'��G�)m��qv����:�=I�}.��z�ia�c�u�l�F8�-�؊��9G�X�8/R���':�2v����~�p��PYI=��J �M�.W��y�m��-�N�B��� H�y��k����׶m��l.{'��=l�߼y�^�unԘK�@��X;l}m�Ð����(е& �7�CV���o�8A6@���X_$!���:��g�f��ِ�Sqvan�R>��ڄ�H%
��B_ ��d��:Z�����b�-.C׎)j�K<[�q�ԅu������#簵�
�]#�+
ښÇ�����>`���?��F�GK  a��X
�3$;g�(���W5|K�`������7�P�2�v+�]����bK���܍i�O왈޿�b�բ20�n�s����f�0@�g�#��������!�G
�ڳ-���хÊ��/�;+�wpÞ}��9�j�\0B�m���$F�Nim># �넻:Ƿ$�³�,��XU�$�m��� VA�*�Z�Ti�����M]O c��1�`,0��Ō��T�H�S8cv��Z֨6m���蘇g_�T]���1�@�&&����M���s�T:"jw�=����|P�$[�7$I��o%�Yc41�~��Ȕ6" 7 ��������k� ՙ}H´��4�R����d(��l4h�:6&zo&e���E�*Wj��%�G�FN����?�R����3�ܩ�������8�Dq���"EK��H�}r�QE�A!�& �V0Az"�� �/?S��Q���Æ�K.�];w�u7��
	۝�HXPgZ�4,�R7�\���h�_?����3q=(�����?t���=��LS�]��T��b���/,æZ3�U4�x\��W��K�cɼ�����@�Ǽ���y�gƆ~��Am�����y+s����-�-��7���{�[a�)�(g6'��tMz��cT��4o:x�0꛷la$�����hD@0��¼Hn7H�g�Zk
��8�۽�I?&���,����ռWJ[����H#tͨ5ϯ��f�lԑ>s{��\4�8h�o�CC�R����MM��酝�B����ꍃN�0�$�m��=�� xn��R���ɶ;�o�Me��B!���\�>�5�l!
ܦ��E� ~bR�3ޘ��[P��ڱ˭�tʯ+p�-�-�b�R_�X+� ���j��DE!lL4�b�jp��O ���ǟ0���^Ti::�K����7�$8>x��$�1j����8��,]�r?dr�YE�)���8�s�~s�:�~Z���L8��Z)d���h)�A��\�)�y�Q��H<gu��j�*:��t��������({���2~8KU�0�Fƥu���֭;�~�����S�ıTH�������(�,���W_���i�	�>��C��[�&g�հc���h�3�([ۦ�Rw�Ҩ|
���Ln&:�	��f0b�u�uE
�Mȯ���F ���-����B�L��� <���~)�վ:�T�e/��"��%7>�%Ȭ\�, �Vz�,,�s�r��]�"P.�d��.E_�����t�ݺ}�w�^:��fҋ(�I����1��kwu��v�9��8`���`��>��kA�JtoU��Y^�gOU�$ӹ��ػ���
��UZҲB� V��YAU��Y��]�X%�6.��e��BU�nJzBCg����Yݷ� C�x���g�s��t�ぷ�zU�0	`�Z�lR d| ��Qr���%Ǖ*�w�0o���k�w	]���  �Hkܺ%��@�W9��H5�u�t�3�s����{w	�:���z�*���:L��,2�c-�(VL#���"��}ĵ�}b'�5���xA[Qhk�JR)$zF��x>�R�n;s����@Yh��
�������S��2;<pFT��7�O�w�y�@,�k��>��-��Q|���IZ.��Za�֯�I��6�]���奄.������ �D�;φ����k����l��S�йW	K�;��Z��2��,��5��84l����N ���i������y�q��[-��f�+��A�"�ᡢ֡5l��*Wv��I"�����Ո�҈��Sҧ8@�SO>I#��<��O��N�{SI�\|P �?�(
V�~�!�`<�tyR���S��l�X[&�/R^Ҫ�#ͨd�q^8��lQ|��W_1���2>jU6�'�����9)wcM�������n�Ɇv�Z��d��^ٜ���7�`��nif`�3������9$�0/_���{�O?�V+�C��G}�N~r�}����'�|��ܹKd��5^�TX�g�O�%$u�+ �r��� H�O�q��:�m�6u�ؕ���,��hj���ZI ]2=��R����*1UT[˔90Gi�,t�tےg�ff
"����8A! ��4�ncgm����z&�N����3������#�,����<=�)'75�)-De5�T��!�+sr�M�Q�x?�V�s�}��?�� �Cy��v�.�]��>38ˠ��>Dm�J6�P�YsxN �,��JF��e@��I�y�.�� ���Ņ"G[j�и���Js]�P&�O�ׯL�o�p!&f�?�����9W��Հp����s�Y���OJ"Έ�Z��ީ�T�b��������N2)�-KϏ��j�J�y�,XF��܊���H��D}�
�J^_t�� Qݼa�K���j����`)��0�,�~$"-cރ���R���.5�Ł��Da�#��H~@9��G4Ւ�<�����r#1�ۉT����%��Q��J�;����ubN��C���2�������ga�<�^#�EFUtZ��U��eTĉ�Z5"�q��Uw��5����l�T� �T}��`r�ܽ����死~�	��,�H/-�Yj�y�SSk(>�.'�Y��ӻ�fZS@��%��/i��EUC)^\�����s��A o4���W!�R�krOS�5%�le2.�aI����._��������_��;���u.U�T��;Z8�B�\�t�Ÿ�;�x&����9�#`��$�d���
x�F�)�l��A�@�C��Vt�F�%�%�(�5�P8�\C�C�����ñ��a�`w�4$���
���5Xj��Q��t��AJ�?b���R���f�iQ0�iN�@���mhF~�X�k`c��4���sU7p���N�(}`"�U|��q��D�49�h�G20a^Y��q6Lp��]�v��E��v�������˯H���}� "�DW�e�	A�o�5ك3e�P��U
���2R�ʡ)��drg��L8rXBpaxn�Z�.g�_&u�6�B��4����)�0�N@#�I��ڶ(~��݉[u:�EC]�	xe��:�K}�	���aG��pp�� ��F ���e��ao�Q9����J(�������5�Dzm�����@�.$�̇svt�t���2g�$81�,�Rы�ȷ��J��=K�ŤUu{k�����.�[pw�ގYn�t+�NǄ�8�*�V6U��\P�Ȫ�fC�՚�W8, ��9a��Dn����t�-�dI.���/�ç�5]lf7<Cv'7''��L;�ծ�t�!�z���E�6N��@Ar����mMT꘎-�4�HO<Q���㿰Q�u�c ff�c07�j�EZG�v;�wj�B��{�V��jc�S�a�ą5]]x�w��
���(06�ۓԋpo�<	�\%��
�&
R#{��v�ӻl3�უ����<��i�ݢ
�tO�����M���z7���3���=�TY<z�hb b�������J�Ft����]8Gn6D���KA��ط"��+ �ɩIr7<��X,2�'\�F�|�qu���qAJ�FDst?��S����L��h���[T�P��lf�I=j~�����C���MQ�耊"��^���e�+�A# �݈ؾп~�\�R[�C�;�F!�$��%7��g��أt�D��7l���ݯv੣�؎,��)Β?$G�ƿ������`>"E����kC!�֬U���U!���q-3�M�W�{�q�ހ-�p�+�B�$��'�1@�H�7��Tb��l[��C{�6����Za��FQDq����35�����a�{0��,����ˀ.�A�(��<p�}��;x�w�'���wY(>��Y�گO�v�/]f
���<�fz��9I�G��~u��;�h��={��ʺ!k�������G;r-��sH��SN�X��oi�-�<�SU�Tm�!o�a���T�������3�ko��_3 �F��Cd7����:S�V�WW�ڂ�]+k�n-b{��0�̓�^u�S:A���eWTm�p�����n���\E��_�Ɍ��g򫭽�8��K2#����ǅ�@רa��5�J�JVE��1��PGd�@#�u��o�f���8p�M��%-s���@|� \+�����Ǖ�%:n���w�iu���xߢ��!�a���䐙*�V�7֭��ā��?"H7�KY<S��/��f.	Xԭ7�-�b}�;˸wy�!x�ܢ�gpQ�^k��i�b����E�9kt^��I�lp�\x-2�Wc���� ,)��y4�Q��ڵ��� ~�z�I�vL��dT)��m��;R�f�1M�aR0;���ݮΞ[�L�� �|YI )��5T�'�Er�Lm�ă�_0-�s]�z�����[䛉Υ��Y���TZ]��˅s�'|��� m�n�t!o�8�{�����s�ܺ}��Y�e�^CF�8��7S!�?���Mn��dh-,��k2��M,.�^g>�ܲe��\��4�~Z�ͤ��,P���k�p����Ħk��M8��QeA^$�#ida�r���İ�lȐ�$qɋ�ּ�F�-W_8�x�zC�iW��V�n��W�� �D<�܃ձк��-��z��c�wu�X�NYW��{���k�pSS�e;����W��/Oy'�{T�n�25���������*�kk�re�"�Ƹ�~�B,FPu�?��ݣ��%�S,���?#8#�w�O��T�lt�����?��'�$"�!�f��N�)�l��\���s{�W�V&�-�H��	'���ٵ�_/�Ĕ�Rۑ�Q}܁H�E��	Gt|\�4䷤�+h�~�}�\~&<�J"�+=WU+6ʒ�jT,,� 7w��=F�������;��7�݃l��۟�X�Ŝ9f����-+���E� Z+��qV������ �+�6�H'��2����Ż �f��	�[���1�������j���:#֍4�0�ʼ6��Z�����p?����cG�S۶����|��W�B�[�f$N��4�����wP��~RY݁*�N���"�'*'� rOj�����"�e4��CU�Y6�> yP��Κ�UA���y�mK
,u�m�5�A�f�rSX�2�r�9���ƛCė(�I��H�]oظ���g���J%b3���f�Q�����tR$M�,k�b\�J�XĹ���u"��������e��Mb)J�D�(��&�H���W9�]zP5�Wz�x�;��"yx��Sg앍�<x��Ƭ_�N��s���%-Ke��3#�� 	��4��¬���<7}<,<<��pK[<���Wi/���a�2q,j2̃����|����f t�_�N���~��� (@ �#��$ j���
%�Z.�DnA'��%�ݴi��S�����@h�Wx�h��H 6��P��	�S={z|:Ʀ�B��
u�a���s����=�ox�W��T+�#�l�F���/,�L�V l�?��nZ��f��#E�
dQ�E꜑ف�@��UQ�_�<AKU�*X��,/y����;n���.D�Am����>������sV�/�
��ʠ�i�J@m5��󄣄��}�����v;�F�8n���s0S�������U�����$�x�����-W�qC������w��g�/*��őmus:��H�G�d�.���G:vI�� u�pU✹8��u�c&
�`o�E�L��s@�ۀ+tV�{�6�Zx	��&����8� ���|�I��C�C�'������="Ϩ�6��E��<7�2�n��W6��Y;K�O2^�ۼ�MP����3��>��,�\�j�II��k������w�u�Vc/y'��w�I�p.P�H��	����;Di����,�Sn��i�^���Սu$0ʄ=Kq���t��s�_��^�a��r�sCq37���v�n���{���X�B)��z��TU(�Eҹ��Z����变-�R�ߓ_�e*�LOO�m�}��g��pv�p���9gm�m�� &��ǩ%v=R,�	=π�Q*g�h��tw���m�m�J�D^'Qhi�lU��8Q��P�0"��Q$��^�!^�����l{�9�C�����,�drְ?��ΓF��r��x�y��TC{�db
j�g������SQ��rA
�v7Θ����8�9)DVg1ڥ�84#䶚�#+��5�-�3m͊<��@� �a�i���%��E�o`3<p '�M���L����%g�u�|R�����Z��U�|4��xD�)F%bjA�<U\z�ťy�[�wQ�3��1�����96���;����T[�I��G�HI�`w�#���zBk�Q�ߥ桾�M'eɠ"�Ģ�T'��I��[���z��@\GQ����bF�xvT�%M7Cָ�ڂn�8���؀�dϥ�SY���-W�`���""��LZ���PFQC�6�ZJ��c:N%����D�Ћ���o��I�}<';�������?�����E�٩���t0�!��bt@^���o޼��ih3��*ؕk��%�s`��� "�0��x����VW�� W��#�x� ��ڳ�g馁�'�e:ҕ�h)rʨ��ډT*'�6�b�1���
��>8yp���z
T��R(_0=0_ݽ{7�� ��;�n �RFH��g�[�K��C����D�9��[�Nhu���R!r���ك�YKD�t)dΝs��\�z����m[��������.����ۼ�m�@� ��ԩS���uȚu�z%K�����wa��F Km��g�/�q���j�'څ0�6!W��_f4Dҝ���x��1|��:d��VU�,�(@�k�9l�d�a�P�̩�������E� ���4*΂vnd�h�?.j����sl�^��@��z�
3��a-Jr��x�R|ڪ䂿a�[Q��֎}��5�Itp�C��~�O�~S*E�ȓZ5�z���f�e�Ɓ�.~�K2�d�`�d��q�'k�k&(~Dj�\��W֯I_��^����0V�*+v���������a�3O���e.K�d8��-���O�e�:�v�F��(�7�2�xs��w�'{Nxo+y�FQ�@��C^����jޞ������qq_����)���n�^��Y�����j�D���H�#����ܨ��T�3�s�~g���kdLb�n����5)(���K��3z�+;R�Z�o��J>7:�3G����~��$�at&�ƹ�Jd�-��Y��pͻL�\/�mO3Q�Z��͛�{D(r�5����XP��i����ssIt�dԣ�.a�����<�TZ��|t�Ω4bQ?�� �����=�"��W��.Im�`#���
52ib ��h-*����ه�X�C�s��P��Ҭh���|��།������ܖ:Ab�[�J� <�+v�?/�CpB��f���81���	�v<�#�i�U�Z7(�����QmV�.��Z��jj�Mc���7��*�S����lSޘ��{�ʘ5�X�;��P L|�{r�Q4Y(������ ����U�(%>ڼ���t�����{��0>��{(�9g�!*�C�8vy�����<���XՎ�C��@��m��NZ�w�}˂�S�O1|��Sl���`��&�:W�&z�m�	m�9WE�cA�,�`U���m�LN��)W�Ս�7��S�������T�X�zM�g�J�q]� '�\\/��̵V�J#s���ݎl��J~��M�?�it�@,�-γo�~�iX����B�t��7nR����~�J�J+>� ��)�_~\�k�π����͵J�g��F	cv'f�#P�@��P�"=1��ݏ�O��o�6"����a��
L����ȍ�h�Y��	3�-�RP������,��1�]��	�Rc2�vM�m��� �o�E��a �@z����y�R��Ri�8[A��}ƣ��I�<��9��+�}�q�R�k+ITq mN�,i�Ϝ{�y�K��Ї�_%�Huk^���A�r�U%��C?1����=jTCאeѱ��Z�������ks)�77��L_�fg��l���J�L�^����v�L�!�E4n^��,�/D:���K7;��!�$#W��y�L�ks�!*AϷ�)�,[$�C�)� �Ҍ ��c���֣릪�@s��h�y5�C+�7h ���7����� �[۝@m��u��������2R�o�������t���BEp��6�u�6�^x����_c��]�s�@��	�׉s�6�Ů~�\#N���o�����L�h����'�i�|2�:����h��\��Vb��'�w0���`:�mN���FA>�gp��Ν'M�Z��pR�t!�ϰ��"w�����=���3�lXi�k��bS���de�"��h��>w�&pn�d�b+�J�m_�Z���j>'D�!���B��m�x�֫�X�`���iSNq����.E<�q�RŖڃP��G���h<��|������K���7x�X���@�ϣ���Qm����s�иV��m���ȩ6V����7{�$+ �g�����A��v���v-�((�����O���@;x��++��=f�6���=fOyfgN�)^@�[�t��G|m)�4�jq�Ƴ�,��-T6��9#Y��F7�Lt��d��j��=��ݪ1 @忶Cv�1�Mܔ�fت��DBLRF�C��6����`�*�16���l����0ꞌ�!�XXf�E>��U���u)�G`+�H2K�+8�Yrˬ�{����>�|Y��X�s��r��J�ԣ����|*��C��|r�����k(k<���k�Ms�%���c?�� *�느��d�����"�+�@�<�xXKDDv`f`(����E_���sl_m�7�b&����"C��޻o�y����Z#�c�A,�ҥ���Qw���v��ꭨ����j���x���������s�aH�x�!t���,W����NuȪZdw��RY8{�A樊o�~�OZ�
��g�ha�O��)
��M,��Fy `xمl�z����o޼ņ�}5z�H�#"	�a��*�=h!�	e���,�lQ�rT�D7_�s�Cs_k��Y�61!]7��J�����;��N��Q͞�56`i�R��^��d�@UA�����{Z$4P	>��nY�� B���*�ꠧ�\:gS��
G*�������[����Fe?��X7�݊�!i ��g�1��!Dͱ�Q�[9��7md�e�Z�5"K糀�����8��L�{�v�;v����R:������z�����~��,��4�<��%���,�tV��R�\��A�g�e�y)��<.�+��<ص"�p��%�����X�2SV�goNO�ܗ�iS ={os��!Y��%{Ah{�1|G���"pL:�q��i�R���tO�l"���Z���N���/ZQ]S{���q�契�X��U���4�|�saT�Y�:'h>�9'2���M��р�~���F�8Lp0�ܟe4��BJL)��mކ`�x�;��$�?c�4Ϋ�S؏"%0b�@c���͡���c�x5���&b�O�$O jޙ��4m�#WO�VɰT2f *�zD��ݬ|��hb ��&g�tU�)�=����AU��6���G9	:�C���>��!*jGnJ<�p�O.b��tYb82C�#��}ǟ듍�RJG��e��})f�	�¥�]#7��suP{y��57O-r��q@+VD��|0C �h���Z�a��1��B�1"�fӃs^S.F������xg��]���iK�^��>�`����|��[�����Y<��D\/1dm s8�D�Ǯ�,�����ύ_t�F$=��$�;x��aBt���! ��h�@ss������a�֯��9 #�����ρ�"��kQ ȅ��ܘ� �,PP�J`��J��
�2��IӂyÊT���<)��k�جB�2I�`<F|��s�2#|�N`�b=u$�Ў�ɪ�io��5�8S'�R '�>�������xO^����*l2��1W҈���{��	�������ӯx@���wH�1�|���������~�>����G(�[�_�N��];�-����^y�%j�b����*��
3;���>���1�F�1��"j�*�� � ��u��#�{��1f�p,�]��]�b��p�,�Q�D��iQ�EAfㆢg(z�����'���L���)�$ϗ�1�T�!Bk� ϊ�p���$����E���tjMfұ	O-��(���_ɑ~���:��$۱ÁȲ����<��)vl�|G�]��m�����'	,�p'�D�eܟ �0�:�˔�lv;V�{���O�/���jHX۸H��?��]���z���Lf��b5)Y�q#?2��dn�6Xg>��c��������C	���~������ۯ��{��^�$�'�lTbP��g��w�yǝ���ͫt��{���~Ws8W v���TWY��U���k�M]�O�^�=J��B���ǩU�����,L�G�JtqI�����彑9;���S 6�xS�Shꊑþ�Փ�^Ū�,T:[e��l�x.Y��+��ύ���ݝ�DZ�{K�Z�b�q��{e{�J��cLS��e1���p,!S�۠��D)B�	y��X�#���RGG~f�IS�p#,Ny��xl#
�nFm�8% ���ܸ7([�n%��t��E4��d��*)P5��y8���(� GhU��\�Ζ��Vx�XI!�y��o��R�5n:K�@Mhf�Q�ځ��"�ך��4�E�G<{9���~&��!�ͯ�M@�b�7�B6<�ǡ����sz�'�Ml؅}�F7mC0�zT��B�� 6 2 t�i��X�^��9+�3M���i�s����$�g{v.�hqP�@r�����J�li����?0�zi�ajR�?¥��TK��@�ƕj�?g�\��ӏ�6������{���>� �X������_�Ѕy/��,�����E�oP���Z��}��]�pу�q��Ş苳qDw�ri��1F�~�H!d�fgJKT�`���⍛=v�\�?�@������&.-��zT�x�H	�~���,� T.�
��Tӥ=�4�D�i��6hÒ�^��Q^�y]Y�6S"�؊�y�-������y��]o��}}��λ�N˒:�v����/6����%�'�W��!�R[� B��D�̜f� ���p�(	�h���k���s��|k�Ě�pHM[�v%:�	��p���g�y���u��u�g
��I��v�[\��G�ӱ�	w���D8/ ���}�������<:���9~��F$J��A1�ӧO8�3��ߒ �( �eJ���h�?���=�ϋ5����� 絧l�$�~"���K/Q��Lp��<Gt����P���-WA�9����?K�)���*VڤT�e���q��c�~���y_|�%7=���0?~�?g���x��e=cn����W��A1��E�̮^����
����o��^}�u�F��7�uffi���N��L�sN[��ihMP�7ӥ���n푍���VY��C�S��,����P�H	�z�� Ee�H&�������K��Q
u*V^ �Ƥ�e7n�V�?�7n�����LT��@/�k��
�����J���,�3{sD;�bF�U�X�n���˿#p�h�:�.7�Z*�Ċ��n3��vԈ��E\$-;�[�I��q�uFW��Yd|���ʼ�ڽŐ2?W�O6 x�H� �%�_���ol�H������(m I�Ӓ�k�[�r�b ޢ@YxΣ��P<�sf �
Sawk�:���g��h	AV���D)Q9r��EB�
�p�J`ԍR�W���Ȳp� �C�gvv޲m�v�z��(SIfƢ�6ޚApU� %�C�֓a���'�'�U����\k�i5-(KRt#��z�w���\�9.al*� �5o�H�v��-t��Q�w!�U������NB���d_hE��?�G�+
ذ��������ĪI]]��.`w�����3���@6�E�W���� ��捛���S~������D՞�uv��de|�����أ�4�����X���w� v�lA�`[Y*5�0��k�!��vX��d�iR⦒�[p�8f�"Y~����gn~Qڨc�Yf���n3��4�1ٮ�T�Eg�7�C_���fQe��ce��,rKg��T�\+� �� �Þ��a�r����QF�8{E1� v{떭��?�)O�XG-xY%�ϙ3ߒF����lo�;�׆$^�& ?�A�o��<p�{*���?�qW��{����/���짬E�uhKrj�w���=��D֭(>����3݂�)��xكA�B8���V�����O���s��m�7�#�Af[�ܴy�۽g���p��"J���/y�~�s�*�O�o[7o���F����Ň�SFF��}�\0G@C���x9|�6z��?�z����Й�i�޽� �@U�裿�o�m@���wz��D�w���}�r��lgV[�����qN�&��Fv��?���B���4���O�qW�a�HR�B��}��d��- L��9Aak��>���_8-r�ݲ;�
ٔa�IjQ�@^��D�����L��"MJ͢{�� ���Aԑ�!�� ��O��@d�Ү`8,�:�!�(Åɷ�������8 ����=vl��n�����Y����3�l�]�馐�D�W��#�E1�g]���k���s�A[n2�����1y^�#�uH�V	hЍݏ�I�P'#���8?��u��(d�����&�!����?o:�1�'�g�%�\9-$
)@W��v;pmml�k+,��Y�Tji�|u��l����*�s�⿗�����GK� 3���e!T��2o8/�@�G��Bw�,�����t�q��ޭ�wܯ��u���[�msG�a	:@=)j����>w��mR]�����l]��&"�K�捇�	4�}���S۷����V%��:em����?L0��ң����1"��eC�Ѣ;6^�δ�� �|�.J�v)5ΕT��!��~��)�l��M�aW�j��[a�`5���z����x.N'��>���Z�=����/EZ)�H
�X�q�FTz�Vp��&v�*)Q�J�1Ɠm��_����stF�����3_����O�Y!���[o�~�b�w��WP�Q�-�L/��o/"���K�?��{���97�}~������l4�F���o~3r�=nm��fc��b���D�Ф��#�R�C6�%.z����>��=��������n��4o���/Y|h
A�?��;z��/��s�������V�mw��&���C���{�>��~�w��E���4�H���D��>Ԟ������eƏ78�{��g @;2��YML�ю?j�4��2�vC�8	u�N\���_&F	����z�l�Ԕ��� {��#�_���\�#>�i����С��Mz`6G��s A��0��w�b�opG���7��ׯ��wn9Y�Z���������
�7l�H�	�H9IS1��v@����9N�=�G��O�M0�4�C�s�v�XNOO�
Y��A�w׼
^�W_}�t/���-ڡp �5>-����c(��9j(:9v��7��#H�˄�76�6n\�^{�5w�O�m~|M� ��h(����Q���%��""��7½����9����#�����JR�֩s�h�j�c���2fa�4��vݏ*���Vn4�u��WI��6��u�[�5lٕ	���� �*�I�ȗ���M�5pcU��<":�Ce��B�qRl�I/w#ǂ��D~�Z��y�`��=��
�1Nd���3�eu�SZT �ՓM����bdZ�F:�tfZ�g�R#ߌ��^_
���M�B���1�#�h�ͅ�oU�M�_�<� �����{u�D&�;)���
��R�� �9���Bhw_�t�6�ݤ4�a�jJ͡:��!ػ�_}ͽ�?�Qb&Z�n7���o��<�����ǝ>�w�v5%�/����z�7�Jt�ܴi�;��	n��xa�bP"�䇈}V�e1��%�-�	<_D!����.l��7�Gb~5oTCr����*�	��|l�R������]��l^+J�k*���5^`�Z����S�M�t�J��V��lf��(X��ӷm[Ź�9�
�v��i>7<34.A$v�{���C�Ӗ-[�` ˞;��Up��8�L-��u��3e���}����= D��?���G�q�mnz��w�eЌ�uҦ'�4���F[�87�YYw"d��ݮ��B�
eu��@3J~GX59��F��͛�pi@=�_�:(� ?��Z�yG�	]A�V��p�����c���K/���g ���� %g|r�Nx�{��s��6K-�'<(��}���w��]�0�(�����u'?��]�r����f��c��i^`��v��2���\�h��O��kЦ�AL�x��4��Da���G��A�7tr�A�-��'?!o!��0}���d�!۷w�;���΍�,����y��ק�ǟ̳cY��P�b� ��)2lx���%�����{�Jr��jk���c>Nhx�/���{�/ ��EZaa��{����+��BO���L��8�@��o���	͍�eD�N =��}ZB"��� Up��qNZt��x����'�t�)��;r�{��_P�]�(^��Ң7"w�L��g�h1���7��5j�p�����G��!�ČƂڸ�f�h�����Í)��s7�Ԍ���.��Q��Q@��Ѭx���
������y�1SO���0#�N �8����Ź!��8�F�y+�%�zg�9F)˳�Y�=)�U����r��`�%��VK[���.3QiK�<���Őu3�T�u�I�Q_��;/�t=�א+p�uãbD���^u�R{E�F�����dq�N�.�:o�]����w~��y��ע���/�����&�<�,
��"`ػg���/���x`c\�tΦ)���#���6p��/�"_���a��?#Ջ���ʫA������z�g��VGbX:��]~����wP�y��302�Z�+��b�_6w�l��TGh��8��m�c�#;�V���Z�(�7p�\U 1�i[��f�ѵL��.�A���3FZ�H�Ќ!����7`�F��4�=���;Ꜭa���/�@8 �g�)ұ�	C�����sg�9m�^8"����4��s�o �a����'�\rs\!�h���V��9�a�:7���P�*R��a0
|�A�؏�O�҄;�!X���:ɂ,%��b�z�t������S��
��d=�`��������pp�ݸN;���ڵ���}�%ϋy1�)i�f8wpԦV��s��ƚ�kd��"D��֒%f++V��-7���5?��!)�,�tѭ$�Lo���4pp���z�g��_{ ��?��)�3�������0D�p`��3�#h���$�8��� n����M~᠊�vqq���#l��H��{�����mr;#�W�ÿs��6O|M��r�xA ��߽k�;|h���*Z����믻C��G~28W-�~�J#XM�Z�B�����\�t����������ګ����Fh�p�������|� �ƈ����?���yioz�Y�	������ �,l�2�t�񴜔�_s$��P���N�_�`�[�Ŗ�J9�y6|M�cl$��i�a�[�	���nԦd���N�"8BQGi���1@��!�Wg{�Q����
5<
�0>��e��XK������`�Ɠ�c�֍m=�=`8�H�d��)�^�5�n��ڊ�)�5��a�'ֹ:�sEa��Z:��0`�3UR0}�$��K�#;-���2�A�S�&�~���z?Y�v�cQP�H��ё�Q�0:u#��y�^$�LZ��p@ i_���$�b����Ҁ�MƼ���@y�5�$ n�9H�bO O�drl<��;֖ku��C'��Pq���>��G�`��nFpMO�G�P�.��O��D<g�;΁�C��gVWܩl�]���m3 Φ��G����%U3�#0i��E��-c'sF�����M�=m�a�X(D����X��Q1ľ˜�BA�Q�R����y<Ѐ�o�BQ��V��B<|��bl�izT� Ǔ�< Ğ�6�w�p�H���������2�]��F��|(�Rt��D�I�p2�: x����"�y���I�����R�x��G�VmO���0��) ^�	�&|�t>l�0\��5x�ڶ��<���@��m�y3��`����t몸�#:S��`χ������'���;R���{��9># �'��.*6��{�r��}{��K�e�&)�>~�&
�����+y�RH��I+X��cQgFDםE�}�j�+䍬3E���U�?�?��+�y��0>��sRoq���ܺu����P;��~�� ��	-���b��4������Ç�t���S6 �	^ƞ={ݮݻH@E�;���;s�k�F�0i��ydC��"|_�(k�b.��C�t?N�yPRp�Sax}������gmNf�v�}�YR1f�xO�����z�۷os/��=*�h�����*o4%�«%^���S~����UV6c����ET�UtI���x�?v�����n�7 �>w�yt�B�8N�N}ͨ.���ϸW^yٟo=?����gbt�l.2��D����܀�l���H>#�(���<��`�D�L�����cZf�\�saNԢa+���t���u����/MѰ����U�bY�κ)j��ZWFi,��dZ)�j��B��p������/-�W�S���`S貽)�}�Ri[����v����F�2�D�R���H6��%-ō���$��Z��ժ�G��ڜ�蒳j^�o�H�QL�WUA�]�t;R�U�k�'�gD�y�F*�^���R������"Ŗ�"�2d*�:����3FA�gMyQ(��N�ȡe� +��91֥���~�w� ���@z`�G@�Ȱo�ɜ)�Ҝ���E	Dp�?F�;gOi\;��#�~~������R��6H)�V \2f����r�GXw��njc��_����a���t7�}��;ה{�T@�k��:�ׂK�,�ɠ�%��� *�јt2:W�kbr�m��
E�<����8 B�)p6 a�>⃖�$��IF.��b���^�H�8����XP��s|Ȣ�y�
L�v[ڱwTEE~�.�zH��`��R�PP<�����}����(�{�.;�![��w`���Q����{~�=���C�0��B� �)S:�E��4���ٱ_|�c���zB��/�$�c��1�	��Q7�ϻ��y���0Ʀ�;�L���>�} ��'(���1�B�[ⵀ��q�:���;wq��Y�3�l@0~�`��TX�أC;�y�H�;�I����'+=�~�L�/��aX����7l��HD��W�ʈׁf���w��;������BmݾM:�!���ɓ��`,^_p�.^h)2K����z���Ku<�U� �n�rs�K�J��޽{܁�x#�X��D�.�<�9�v��o�y�ԙ�0yMް�� ���� ^L�+W���|���\��v��A�̉�2;Y�����$JLD�Ф@�<�LTL"ٰ$\ߡxu;(.��Ҁ�:t��	��������'��w
 v��/�u�ֲ�׏�,�,�����a�BƋ��X'D�L �
&�"1���#���x�������S!���~��<c!~�٧�C�rE���R�v�7R���n޸�q���M=�՘L�II5ijF8�#�Y�:��E*���'�T�5��0�]��C�|�xn���i��19�>����[IT���{5r���1�B�W��,PB�T�B�5SpU���v#O2�U����7�
q��v��n�^��8W�c��~/�i;g䗦��^}Ui:4�5�Ţ��҈k�H���
m���ڼ �*څ���e�g7�aJ�^���3�m�6�3����[��*C��|㳪�R����"2.&��F�K��c4���烪��~�}���m���-1�<)Q?������Lإ�O�%/���\�Z$�0��i��_-�0���3� �!6�kׯ�'�?�z�m��RI�Ӧ���YW�d��`]+�s�$���C�e�޽������!j.�Is5�L�tsLljc�:(:��%�7�Ni~Jt�riۍ`Ϟ=���4Y�*H[p����ю�s�F�����a��K*{�C�Q�GW�O�Z��)�7�q��t������1kS�*K��[�D��][�,A����ú݁V�=h��M�v�<�ءM	�\�L�5�,��\��<�D-mIN��%���� ���E`W��a^���X��<ֳ�#�fO�1
�jR���3��eR�	�̛�>G��b������5�	n��d.m�M���?�H9��o^o/�{��^�J�8�x��d ��	�i|I�춹��� ����3���*MxZ�5ɢ�S�YD��r7VK�����N�&�Q�'<N -x��vAn��?�C  ��<r��t!2��O"��c�ǀ����*8c/]mN!� v��A��ET�L���[�!�Cc��[�S<h����.-�C��C�$
�п *��&R'~�=w��yzҗ._bkUDTPx�� =��ޭ�T��FBt^��e ���ĉg�i�kO�>���?��mZ�1�~�ƫ���,O�o��NZ��{ņ��CH�{�uݾu�]�r�׋� � :����%���m�ni5�9T+}8��4����d `H������q0ͦc�e>�����ꨥ�3�P�ƴ�H��4R!�kI�i�k�.���a ��i�P�������i76����06 ���2d�b�I�f�^p��/�_SL;��G�k8A�UK�ce��������3�(�e�r=_��g��{X�	�\��P.F����Z
�&�F� $�FJ��g�V��Jjoc��%���@�1��
^�T0���S-<�9-7�]_�mɽ{%k5脷;��ɏ.X��c�u��g��%�G`ke�Uj��	N�ڦ4>���3�aY<W�8F:�5J]0]٦�eI�*d��.�x��h���Ct��V#}�sbla�$�'�)�s<K�jP����o����~6��ܢƳ�x�RX�t���ČK?�4[� �Ji�f'!U�5��eq���[P��4<dqvN�rmB�;�@�jo��	]�/�6��v"��\ �f?0^1�Ӣ#nm�{J��&*BO�Z[d������n1צ��u���Z���ɓ'�.1��fA:QY,/�=�׀K����܇�9EAcz�>����V�.�1��Qx�R�~��"�lX�z�����v9��Ƴ����`����S����s� TÁJa.ѹ+7ݢ�bF����ר���1��ݤn�C i�F�ǃ�Ä���SЀC���b����B�p4RXX�I�w��1N
Ȕ@څU�w��x  ߺ}��k�[[���$e=|n�@߼Y830L0�(���M�,� �̎��Y����Ő��cI�7�0G?P���£�� krV	O�7D�nm�+���L1�y`��C9A��6�
��G��$'O~��z��a@�{��i��Z�q�T ��HC�]GU:7;4��Fܤ@����o
��_s�	��C�߱@ ^��`L��<\�� �[�̂�(�TTg��\c<�G�*�;�1�*^=����(�� N�v6���X����RX�#����`)N,CӚ:�ĨYy���}j��̵`c4��^�i�|�{ͩD��-)i\�Mw���׀�}!H��q}�9C�ё<�m�ZK�f~�{��sgϑh�&��]�x�f�m�7g�aGBD�`����kx��.�.�~�Z����V�*���}�L�Oѹ��n��	����L����Rp�y���]�\�
@t��$� '�`fv��K�%�c��1��zP�4|���*F�&�wb|��ܝ�СT�AP�Y7�ୃ����\r��UXQ���]Ւ"d3H�%G%�­���lR��%ѕ��[��=�[ҬEbo�XL��[&�_P�H���
�{`��c�_"ȅ��T�|��7��Y֌ɟE�rt�D�3��195���g�{�M�=����d�|��)w��e��Pc�׉�D�0,D5 � ��A�K\I{킔Jt�ݘ̛˗%����ژ7~���cf�ส��y��"�z�|ּwd{n˦�|Oh�'�#���O�-�#:�(�q�p�<�c�{�n����F�l|�ˬ��O��V�e���DOw䲊��f�V���W ���hP=4"���w�����n��iʭ R��-� !����f�ü\����'�A)�`�O^|?�?U��}�}跌b/<l���;���%&���D*o˖͔�Cٹk'�l[k�`	��Ͽ���ANnT~Zt"p~��C҄\)T�+�4�
�ؚ�Т7��	X�W����~+����<�K~C^E��a�3�c�.:�� ll6n��s����N�����?D��*l s���Ŭm~z��;unTaͲ38�R�.�l��y
�^�I���U�1	���M��.wX�(�V[pI4���&��*s��VU"�~j�&��ےϳX�9�Ӵ�mF�w��777������#�Ŵ%l>��XWD��ϥ8�u�Q�� ��OE�N�*��4t��?J�@5�۱8�X8b�a��bä����4S��sM;R���xY��t� f���☊7(]r�s�V-m\��4�q���H�}�V�lKhL��/�\X���V;mu�'xM�T���b�;ðu��cp��]�0W٤PȤ���ه���^b��Y�N�1����G����A��@k���-
R�����Ǥ�w��Li�T:R;�����lݵ��t5����P�Fj��w�<xyT�_�v�b�e����eHWSz@|�5�g�a��ƍ��`�^#���G��L�n��5c�Q̸�=ٸ���
�	����)�3܎�ض�% ��$���1�jY&���f/�6U��V�+@��/�(��J�:"�	O~z�5?�~
ou�|���%�dU�/Epȣf,&�	V8 !�
�����o�s7o�⸠S�|(O G�Q]�`��?s6�_��5�+��Jm�����G�!�5>!w!��
�KŅ:��cG�m��0���q9��qr�;l���ذj�Ir�a�\}�<�>�Qy��Y65W
�����gw��`��(� �����d��ت��A���΄��V�Nu�AM������9;J���[I��?�����'8�~!��נ��޽;�&�$5�<�����i��r��Dv��ھ}�[�z��H` � �.�x�%���p�h���nG�l$�(CI�H�c�AFm��l0�\����il֯c��[�J�t�� �B��BJi��f� �$�$]��Sxh����Uu,{��b�s�KQ�tUB��D"�]�Z�����7^"��'�{��������<��O�8�����6m��>����H\W��i0���[��Z፶qTd=F!�'6�P�g�m&Z��3����DU�Kߟ���빫����{u�XD!n$����*H����g�E���Xďk2��b��zM�������אnε���"���T�!�A��V��:R�1��e<:��pzq�Q%+5��]V��p����R�<�xk���<]�^+́B��Do��[���hɧ0�
�3����.h'@���UԜS�g9��1�#��^v���*�fi����}ϒ_�ۧ*.��s}"�F���@a\��"*eY��P�QS���c�X;���Z���ԏ�i)��UC�Œ�,o� x=�\�y��y(6Ӣ��;J�n��ԑ%Ω�+�To�*�q�[Jq6��-/�b�9�"�h�

׵���V��LMJF�;��Ƃ6sQ�;g�X�?P,B���oϸS�O3��H_[���%�t}�2�t�l����u�A�&�m��|����F).~�9�|^�<�B�/��Rd� �2a񅽐-��b���Y���M"�lwZ"�<�sȬ���� �C�t��=���,k"׎�$�#c���]��!{��A�o�����{A�:�v���$�؍���%=�������S�UB�0��l��j1~�u>/�@Q
���tA]	�,�&�&X�����m�N�=�����'O��^�E��T��TgIjl?Oi��ց���u�k�>�6o���sʙ$!�>�՛=��ӂ�H�
A�^R:�� �� @:� ���tKG�:��E'Z���c�y��Dx�&�ɢ/�v�Nr�]�\،ئjb?&zL�������t��}�LQ԰�lI5xa�s���,���'���{ܷ�������.T%Cp����H��ĄH��*X�݄�>x�^?ĝ7{���or���=9i�YP�փ��*���M�.dQ�s�D�v;�e�
�n�3*���(�["?H	�ˌ�$~/c! ����h�q��5���/�����=ӻܯ���V���q�4�{ S�i�w�.��H��g&�%���1�;".�R���5��;
���������P
�Ӫ]���t�� �׫�R5�YP��� ,�BC�b�e!�L"1��zd�"1bh` Dx^��֮��H��Ǎ'��+�x(z��榌T�w�5���z�9A�2(����Q4���]H��r��b;s�ݡS�D�(3�"�w�`�\���ҩΥ�7ō�L���+ z��΅����z+a;,M,�!4#�5��7��G�jVd!�E�����Q�E(Ii�{ȍ�8µ�A���1%��$RG[E���������iF���w�3@��P���3Xnߺ���׿v���}f_z����¤���O���ws��;�)Q���9w��9��I���K�ps`���]�q��T��P&vC��9�I��F�P��Y���~�r����Awo�t����:���zlt$4��p����j�/���P���؟���Xw��m^OQ������Y��4ې�_�[Z�?��%N^%�s�{k���D�Y8,b[hG���^�W�4}	a����+d��f:7ɡE�ǿ~�T���,4�Ұo�>f	���\�A �(V�<E�_��_X�ou9a�7���Y�o�p_}ʿ��\��`��悷=��	��/�e0��:?�>��S2q"+`����.�p������#W\x� �G�!� T�߳��?��M1Џ �a��~�ը��2 x� �焪������*�a�z����Ľ��k�\8�c޾b,.^��,:��3��arM3���Lc\�?��+�LQ�9G��w<pq����42D�Z�g����	仪�˽�֏�*�P�����,h��%?2��)w��^�Pp�kvNeW�_qX�g9z���V� � Y<| YPΜ��b޷o�s���w��E:	�Y��N,��F\6^h��+�$GVN�:��x������/ԅn+��M�Ã��cy>�!�aD����[F���1?��N����|��[�S�r@Sn����c��.vV�
�;W�wO�.@lL�ۇ�N�:���~��^��T��l�h�w���� ���{Ш�ņ9,Rl~��g_��xcI�4t�紫�֡��&��X��U�-\�R������f�]Q�?�X���N�(Vioם�4E]�7��nzϢ5)�{f����F_�d1
}M+<��9�pH��~p��"@[/�J5rk�V{����Ϣ1C���9d<�B�E0N5��0<q��*M�*h�\�u!�tK��񈛾m��i��-�&�`
0�@c�Ti6#v��1�t*�[t�'w��,�}6Sr�] ��AiD�GeĆ�ƜK��@F�D;�y��I�"d��&q��3��Q�Ω_ߠz�[���0�@ې�+���N�f�0o+U�]�l ��A��s3n��=w��u�~�Z�!�]��T�I�Q�4+(�	s������8��<.jf˘2ȁ	
ұ��D��
����wv^��ƾ�{�^�&��i2�>c%�$��s��\u�݄�o�m�f� ;�'W�[z��t}ٛ*7l{�f��=�C(�5JHje䳤#�v	�U��E�	�/��w�����j��laܱ�����5�W�.ؾ|��ʡ?~�Gz3CZ���˚�\BD��H�۽{��I���|.�'P]D�K��X[dWA3�Q�E`p��P�cp����K�.��	�^H����
H�p|��\����?��<g�t�<q��J �j8V:��ѼF�?T� |��u�c�2�"�[\X }����?}�+�mP�7���ay83K�������e8䤮����Z�m�����k�3���F��O7�Nf�	��<��79��֎�v��.�8x�a𳘊u �u��6�_����+����̅�N�G��̈ �H]�q�����������מ�禟d,��@��8����*;Da�c�F
��>�8b��5#��=d�����=njk��w=B��f�dӝL�s����f ����%�rx|�O|>�Y |,���io���(��߷o�N�^,~�J @�i�^[��p-
��P;5m5l��-�0`�-�*i#�<���#�� �,R�8��_ql����Y�o�Y�ɢ�g;)v>{�m6�c��YtX
jo>_y�"�;�܍�V�����Zې6(WKU��!�l��c���m�*�~փ��MT6~��J)(���樂�f-β����k������d:�AA�qmRα �Vm��&D�uD���ya\�3�\�a��[�z���M�c�v�V�|��W*���s@�|�&ok���iY�=�[
1���~1��ԉ,��噭�7���g�h�o�;�7:2��iI.��R���@4GrTd}�oqM�y!�g2]�}�{z���N �-��@�}�95��:��S��L�3���:����N;\C��pX���
����e���nH$�(�%p�?1�+��2��FS`&F#�U��K2v�d�js_�b�H�k�\�\M� ��<�ӟ��qGf q�ƍR��?l�����z0�8�xMֺ���PUB�����8 �[6ou�{�)g�4�P�%��<���;��dg�`;����,w�	�u�5������z���hӁ�z�J�*J������GS�������1ʹ��� ��C�`��QDy��3NF��k�f8B
���7������k�-c�&��4
����sw��m�1�X Ƞ�@ydcβ��<��.������a��ih+�eYdW����~�!P;tL��)�>��X�;���ɞ@��N����_����Q;/�.u=-�u��ua2Adz@�����YXo@�������O�i�V
�윶�m�ÁjJ�}����idf�\Z�nw<D_�H��*P��%`��Ƣ
uw�Z�n�{���D���W_}��$�.�u���ϭ4�U:I] M�Vٶ�P"K�|U�p���?�񏔌�a�w�.�^
�@�ǵH4�%NS˃�����oW�~��e�	apq�(������?^I�����~٠^��?�̳�a��t���,�+� &<s\Uk82�,Xs�찔_�(ÿ)J�9?t�U���e�kېJ�O�졢�,�T�[l�������R�id�)wX3s�$m/]��z�uS5×e���[�ը���'�B1&-h�e���t�TF���(�&�YK#8�@wY��<䜆ȚQ5���d�!�$��A$��1ݸQp��؁���"�_V�H;���>�[u�Pp̣�K@�{��(��K�kh ���[zp�[5�u�W	ǲ7蹼3�( ���`���\�Y�b��a8w}��_"���щ�XB�l�/^f+�B6bVd�'���K}l�
��w<�]K]Y�[$�Q� K:	���c���]��)k+�m�3/��$�h��(-̦��F+u$d~�X�Y�m�f��� ��ac! �Z�Ϡ�!�5?�?�<#�xMW�% T��E����>��YUZ� ���0TTH��c�fI~!:�&���g�=��S�O�������-�q��e�/�\��{��y�nȊ�sw�h2��+qųw���N0�� ��k��L�_��/�b�{���KټH
U���u(� F�f�� �.{�&�̍{g�����Çw��?΍w���s���N���l(B�>�9��=	.�*�isNfLlJ�\Y��[��#R����8ؖZ�M�sA�{׮�L	��v�\��D ��7�_���M��]�TUj�F�@H��G3��u'q�����~��$�Cl���0�$$���ZSwW�����a�OU�N�{x�nUW�ak���[iq�=�U`?^�z���t����O~�7,��>6�C=(mx�Eq��<��mr�Ie�j���b<�0�O<w�B>��}�ث�jQ��aeA�#W׃G���U���H	
��)C˛y�2�I����"����_�ơ���+�¥g��'۶��W�x^t82^@�n԰��98�$��.n�tP F���2
��xf����4V8m�ˉ�A=6�[bW�5۪x5��Ҷ��nc�T�V���PC�n�_�$���{�*|BN�F	���E+�Ӈ�<�u%P[զ|;�6`�B�N'O�VL���6 ���:I+ȍ9��<�	Ʋ9����	kW��y��H�E���5���Ma��T�������q��!F�d^�v���6�V(�I��8�S9�p�tp���p��K�u!]oPB��Ϲ�\��Y�4 �u�Qp�Z��&��E��o���w�#}��s�t��(��[�D���h4ڴ�(���F+�F�`���ER�B�Mp������J��0<��(=�T\�ݟ�ٻ� n2�h~i�����4��ٻ��c�11�	�Y�yԄ w�J-�Y˺g���l�Ȋ�!�#S�3��z���o��o��.������V����?����dp���'�����E*��G�el��T�^$McF0m�-`،l����� ǚ�x�n��Ȟ�����\���#̓�����F�y����tʜWy��&,�Y-�ilF�$d}�ɧ�d>i��V R8�,���w���c�4`�+���7�A'�;�p �
s�N-���xf�����=�Y�D��P�^��N����R3%�h��@��&��Q�^^r)��m ���
���`��}�8Q�@w�@�v��eC��pMp���0���*�)0�����]�z��l�o+�!F�JI�$a蒰���Z���X��"u`^L�W118ZYΣ�¾dEIG,,�Y!uS��#�Ab4�>Ѕ��^�ET!>��S�p���?���߲K_Zv" �������* 1�����8g�'d�����G(^�G ���G�W�{��cw������o��.0�-?��֋���N}q��|�z�O�r(�BU6^���:$ls�=��V�^�X��4aM��|�3�=~�x>
5�F?/������E� X/<B�[�D=۾�W`����#��ٷ�3��Y0���빹:72�K�Zk��]^��o�\�5L��G�Ot]B١x�ץy��dTyq�#o �L�P�͙����/� ֚�}���Hrk��͏��wN#ȃ����)F�.���ۚ���0�:�®kn���F�.}~����u�y��I��Ϲ-�3���6�A���3i�tL����اXT��bg�n�e����S�1!�s����8��.`��R�5��e=Gҙ���V�xJ��O��Vy�C&�@� {rn%�P�%2"#���O���(΍2�l�m�Q|��'������=�>���j�L��&wB��<Џ�xS׳�P�J��>^�f*�`aA:��v�Ho<�hy�W�Z�����^�~$z(�$|��O?��)�%��3��޽�O��of &F��Ţ3M`v�}ls�:k�"h�u��c���^�e��a/d''�W�Ek�c���5B��v�hf2Z��!�o����i � ��5��]�;��{�)#L#ԣ�c8ߵk�?�t��!�0�)�3��&f0=ve����Br_7 �.�{i��'��]�B(�\=�޹��2oEFf&�VZ�sn�.2c/0g�iW�f�<��~�qy^"2\��2%�����[���V[���u��Ǝ���@SK.>h�q�5��d�2��y��s�J��N�L��`=Xc��.�N��>���7V�ҥ	4=�����"�  ��g�p��q�!#u�=��6(_�׳�r�}�Q:v�/V+������ɓ��f�ɭ0-���<pX�,vcY�yQ ��JO��j@�
�?�G���#���@�R(�a̟��Ek�N}�^���`E>��cU^.,�4�t���׹��a���}w]���E�6"@-@�R �t���Ol��9Ϝ���z�2�zX`:�9Q�i�]����6}}�kN[�f�Qh��Z�y�y �����You� h,�S�l%i1 P��J��\4�ozϘOc��J��"��pV�F��N�"�Òk�Q
f3��p�݋�B�0�Y�2��?w�r�uF�,�}ؾ
�����"(M!�F�6��r(ѕuVR�H��.eС����oK1��Sa����Ĭ#�ST%�wz��� w���r�B�OE��G�_���V@K]?�Q��/�l�����B��l��D�@P*��iQ���B�y`<.�[� $tA��Uͳ�`r�(�k�H@�X@��ܐY��J�u�s�&n����埆��N� �aT$�ݦ�K-�r����	�&���r>�[Kd���o��6����<�����G� ����{�������P�W�|����M���sm�U�Z���\�7r��7v��q��C�t'r���L!L�׈<��`T`�Z�2���3q#�`g|���GCIq�4�g�S&���B��s+X�
���#H�RV����h5��u�]!������0c�Xr^q�Xj���Ӯ_h���z�e��3\��t���l��SƼ#�ˏ�5���	;����v҃ r���`���fD�Ģ;o9�������Y�v�Ui���u�s|������?rZ_�`7&<�hebN�5E]45_S��L��:v�mͳ��B(i	��b־��dC�i���� �ܨ�v� r���9�&��f�j����� #�&���X]�$�}��$*g���thK:��� D"8��$�/��d�$�`w%E$b#�!t��E:ȜrK<A��9��&�,���9 Л�I���_��=����2x k|o0�ˠd�a�>��+l���p<�i	h�����,�g��V���}������&�ڒ�Y����4N��2��9	ssS���R�c,���M��!�[6S�K>!���J�X��o�k�Q����1�[U�̂�<�]���W8���q�s�9Sd��dZ
#)SO�����2��j��B��mox����g��
�^Q�a��@�0�A�	2��N�H��ӐT�,{�2zcЛ����fG^G(6DK���]� �r��Ly���Qڳ� F���.I�EP���P3�d�Q��5w�\d�9�2��K9"����J��-��2:V!}
�Y0�����U��6�8���2ķ���0��O�I�R��u��xM�����%}4����7�u\�6���̫O�'��"�J{�)�Q#�i�hiҏin��R��{&芌�֜繀���	���|Թ7yPw����c��3�<͟�e�T��m~�'nE��B������c�0P�kđB�)��l�كm�������}2K�I�m�s�+<ɛ}�/9�[_�꿛cā<�0�&ע�� ������{A0��&+������U�D%j���n�F	�ᖞ�HT�Ƞ����;�Ÿz���>΁A^W� �l�C*l�\�����m�$�� w΢ ����Uy��rvZ͏�.�t,<�P��9GQ��UPCp#� |��2j�##�%��C�#ԑ /��U���i��/�8�	�;�g�prYػ���.x|�!a�j���3H�~�ڲ�XT`}Ki=n�B�{e�L������{�ɿ#'ZBDI�O:6~�
~���q�<N\��!�Ⱥ��ڒ1�����f��3M�	Uà�!�P���4����rx�Jx����$U��'+�NI�A�iZ�YOv��b��Ǝ\�f��8��*���l��X}.����=n�Gɯ��w
S��5��i�慳y�N73�����~��2r�z1���x�?�J��r��ˏ�����Ja��<�6nyd+/��bQ���?n��$��R.Y�y�e��ݛD�nx1$/\�����v-粢A�h�)�,�)V'0]�ٜ;����D�D�o������xO���sij��[gK��������r��k��G� �X�/�wG%���.�;ٗ��B:Λj����r��wR7ZjB���+� 8X 4��\2��x�=4T��̙"+�ү�ޅ�c�k������/��Ч��@A�9�pt��<bӖ"N�D�����J�΄*��Ìti��7{�/;|po; �N������[�t�����|�����᳐e٦����-���ܷ���7��Xy�{���.jG�y�+�m�:T�h��4��ɶrv�����<��CmpH�$���p(]���
�5�������0�� @�ps���_��C!�7`)��A�y-��vM8�%�����=�h��ĀW<�������$��B���+���F�Z%*�B.z�|�9��XŤ	#�]N0_XPڞ�
���<�V�A��o�r�S���`���84�^g O����;#q3�;�Gw'T1�Sw�Dt��nj�м_���=rk�,��^�����eo�98d-��"��ztmŀ(a�>���0�z��'�<�p��{�0��-�q(`�?O�<��fԁ�M�W�F�CU�G���l�kī�k1���mh��{0�{���7���o%1�n���9��6C&_��
�N��������䜮�Ůk�� ���(i���0��cyS M��5��[;�5XJnU����."QBWx�=~�z�eϜ�'��V�Q \n����8}��o���"����^~I g��(�3������0��F�<<�f\[~iE�״Lt�hؕW�րps5+�:��+{J��t�P�z�87����*/�.7�y ��̷ ;��kF��b�Ϡ�*�|trkfQ���>�!	�;KI���<���}w����X���n/yV�7��Y��9�@U߄��:�P������1�����tg�wz����Oy�n�x|n�(�n{��0�}�4�G;3��S3DWj����bc1��Gw¨{P�/��@�	�i��/Hj�`�=6�� �/Q�u-J��I�q�&�Bix�h��[G�4�M��~�;�n�{P����,�ب�l��{U;KyJ����ydȮ-�����a�u�*4Ґ�|G�<V��q?w���|;w��joQxV)j�g�*��=�rB�^<�Rq. ��y�6�߸�UtݘqBw�"2׿*h�&3�y��3��Cij-�A��4,p�������V�
=�_cy����;%�I@�k`�y��b�*M	N�A�`�����֍�B8rJ����J�k�^i|���&N�����K��~7,^3���k�۸���k�@-�=^�}�9x��|��i3Gb�V������
�KW�!j�XB�V���5sy�n���>1�d���}�	��w�ω�vF+�$~�0�����rt���1�3��,�9�֗�z2�����(&�!�4������:��<k.�ڴ�;|~]�����������c��f�h�삭�Q'N��w�}��حU�Hrl/�l�hK�0���P��tD�.�Hn=��=����ͣ�@z�Y̩���@[�G0tJ�`^@)+�[i�Q��T �A�T� 8=�{�i��%�&����K�����A�"-�.(�Fʁ��8+������f�|����˻���}�usLu&-k��3�y��b�s%����]ks����ѧ��vek�=����4������̽�3:=�z�
}�uUYW�fb�m�W�!�F�H^\w��������Jd�R����B����̳����F����s�$�NdY�FTp��0�\�Y�fy$�uX<+R�庴�b��E!�*O�-��l��I�B�%���k1�` ,��� d�h�$]�9�[4�y�B� M�"��O��~�IV��^��M��y�
�"���� �iB^`���)%�c���u��٫�ND�R��=��\44�r(|#;<��)�W��_8D�5#�<Z2V+�Mԍiy\I���*����<��{�0�wA����P��W�g�� ����e���%�	�r��I���O��׸�w�Ëyn�?�75h�i�M�����g�֙n(�}�XȺkr���.��A�+H�ӫ��<����B=9�_j#&S�p4�u&p
#�w���ԻQ�J��q���w��pJ���,������$���u(k �k"bU�"s�,[!��}�� �
�����"rB�-"_;�����R--���Nh�ӟ������3Sƴ�G�:D�ЖTj�r4˞7���U霧7I�K�́���9k-�xȹ�R-.^��p�=�f�;
B�ͺ�����+�� ((lL&�<D۫b�K�3�&pNp6���\��.��(�}2`ߔs���GZ��|���lP���>JA%���>^VXA)�A�5� p���@G�a^�����Lh����������G�vP����~�qa	�:HS|Bρ@EVg�5e�"2<����M{(c��<㢢��X����ω���T�(���V�y��o�D?Z3�_8��χ��~�c�����>��f��;��r2��6E�4�be�o/����y��s2Jq:Ф��hO�Ǽ'%�ر��k�m��A������w�R��U��=�d��]ٹ���`�l#��de��2x���gJ��ߗ{/׈���>MM{�v�I�p�^�dty1��G�0�x $/�:&,9��/�%SK�t^ܻK���C�ߨ��!�Y���W��Tt���W� 2���w�՜�Ʒ(��~��'X�I�g��5��zGVP���g��c�!Q��BXsXY�isC�������ߣ�#W�Oz�Z��n�"�kP,f$�ρb=�o�'F�X�&h�adP���@�Q�uZ�6x^�F��=�GՏ�=�9k�?�.�֛�G� ��G˕Г\kx�I�����Rb�" "����ǀ�Jÿ���Ң����L�%㺾&se����˲m-�H��9�!5���E~|#�=��F���q5"zj@��j�<���0�����3�:޵�.�Ή��֚)�H�ͬ�G��g�52���\�}�O��'3(�5�(�����Rdl�2��1 ]�u�]�P�)?b�"/(��u�(���#�	A��3�����ōN�LW�Ǔ2�&2���dJ�t�w��:��=r��,�G��S���c8��IN9��	�'��ȼ(���e:��ϵ$���(34Dv�aB�;w�/�D���s�C�~͗@/����p� �e�Ș����?�]�~E�O���7n���1úӟ�)�P��:�ț����;�G f�"�A�G6��B�gB5�e��w3�[�i���>�~�R�o��^��s#T�0���ӹO:�*7X�ӻ���	U�a��g�� ���ᰞ[�*����2���iL�z�ȵi�"g��S����%�-�x���}��ݣ>�q����a�q�"���{��Ab,Z�r� r�����Q���	ʍW^��j�L�D��Q�c���u�/$��Vt�0-�a����T�J���
�&wb��s���	a=�js.J��wǤt��'t� R��10i���r���)#j�]<�o��M*��.���p��Ί.�����Bv#���s��S;K6��d"�}�����Y_]�4'���}���:�X�Hy���¢�#6\���:!�Z%%7{֩5�cf��x����*7s��Y�٫��)�,��[;����c>��`�R��;Ѱ2��^�m�߯[�x&0m0?��_�d�6��67�����kW�o�fkR���p3D�	�$����kI�M�Z�x�q�c@�X�1�P�kk*x��hc��7ɱ$��	�gF�P��8t��iJ�H�,�?(�u�
kK��Rb����K�d:�ť=��G������~�a��L�,CxN�h���^2`f�:�;�������s��B��̘��AY�t�&R�U�[S�dT�.�t)pj�̐sfpI�L�vZmN�t�c�����Q������9�@.rv;k�@�����W�.y�{���9:�m-}�9߶kPv��Rt����ou�������gXqSN������r
����0|�6��h)x(��~��%�_K/PC�
��`�/rg-�t��5C�{�M(��[ˡk���Ud^�>q�F�*����C.))^?�W�M�y�����kE�Ӕ�������u�\�Fxu-����U��{��{����Jz�9+����f���Bbÿ7���7�N�����F+�H9�u3&����+F�ڇ�`��LX�.qa�9d~J��&XÝ
i�3��{%eE"Gҥ賤��i�l?2c��S�'}�3�C5�m�{��v@�w��N��xF��ҲtFM���)u/�l,l>0_�:0�"c@���"�J�YS� \�N�y�Ғ>�.5�ĉcў���6:����nj�:<�4=���f���T��%�����̷�T�\�A���2��"������w����	�8��B
��IW�㏵�����v٣>�ra3���ۣG�O�Y�k+W����[t=�+�!io��z���d\���Ԇ��]t�����cl���Ŋ���EuJWB��������ף�P���9�*;p��6�x��@�S�&�h��_,r��Xlz+��+���ٿΡ�t��y�Q?N���L'��;<bm�ͼ�m%����tK�ᮟ�6KyL�۩�����Vή�r�D��h�:�h\������w%���7a�C>��g��N]��Bm%}���i �Ƣ�J���@�3�O��(���M$����-������'�m��IWrz�1TH��p�tIp���FU��Q����'�Z�2@3a��V����
:z/�YOŊY÷�@��1�@o��hj{��l��wڶ40�r�N��=l�0�6e�yϊ�(@�	5>Q�K�n��gޓ�ߺ};)�Ŝ_X�M�=43���qs:��kḓ� [�����en�%�ae�FMşl9�X����������5E6w�sy?��F�Բ~F�3:A|�*���V�  ̧�Հ�䴆l�pQ���yN�Y�����:o�2]���UҺ%�mJ[Gܞ;Hg���L=Z����P�Y20Ԍ�xw2i���2�{{���Ө�6u�)�ތ� @=�9��BA7��Ox�Q#��;��AK�EM%�xX^c.�)ŧ�I��%F΍�l���!4����Un�{���|�[n.~�w஠X� ��.��ΝK��������s	�#�,�pAe$)��;t���nI�7��g��4�=gEޣ� ��%{���͕�.�&�da��Ѹ7���j��d����[��:j���d�L(0u3Dwt��N����/�/�e�2֊w-�o�3`z$*Aa݌{����7�2��yM�+�`�n
VB(s���v߁d�����_i��g��C&�����V�u1?���2�]���+�T�C�"4�VSƵ�������|n�xe�-b��(As��/�:*	o�W�H� c���(��X��ٌ�pU�N�$�E�G�r�*�JFW�St��O-hI=D���X�m`���u�N�g��u���3?7��{��s���FU�j��##ӷ�m����Ҧi�k
I�isÝ��g�R~�ެ�e)��c�
����k�I�]%��n0g~�XAڦw��,���s��RH�]�ڽQ�����>��r0�F�޹#CAX�(��n6��1�4��)(*�2���1ޔg���M�s�|Ut�\Y��tmh3��A�z=���w��b�P���f|W�a��=GÎ3_��v��JS�%o�i}(d�����Α��f��r'Yj24��-�1�s��%z�����:��ݱ@O<�=���t��1�(L�ƃ�=\���[ݺt�[:w�kvFAx���N��:�a�-b�[ZfTSV� �6 7�B��~��W��s<��%�|Ϧ�P��O�;|��{ g��FA�1(�K������19�ޯ���.	��<w��eJDsl���I�}υ;�i����ܛ=Ϙyk'�}����&����轶O����1���дT(h1
U���ԍ�-�/�V-G�9msQ1_����z3Mx֤��N���厊���Q. �:v��)�Fj﵂�n�Ѣ� ��0{�B��#U�Vl�󘶶~h�Y���� Sl�uDn-XA� ��dε��/`s@�<!럩%��7[��dè����U,��O@�>Tr� oय़�w�(t!�t� �Y�7+�ܿ�47�������2��(��q�u�����*2��)��eMΣbt0h�*��#n���ۨs�	�ηf�_�u�k�kW��/YK��'g}��x��ύY���>������L�;�h�Bt����D֝��u.�,��!�:�� �5rO��D~2y�(��\�6i��3��U�5�˖�D�DN�7��+-�mv\���_|q�����և~���XO�ܝ}ځ��%��"�`�]��k��z�]��0�:���,�|�	�kP�W�������bo&N���5�Ɩ���4��(�~��\69�� ���?�4�,:^��7u~���$rS$�'�r��Kx�[-���?5�pz�/�E�;3�B����u�`���:�р�@��
�h�W���ʰq�1󰏴3�`�ܩ������,q{��m(ѶbP��:3ll8Zd��y����=��o�~7�]7��T�i��ɳ�ENM����")�WY�Y�OKA���8��%�,d2AAg`0=��n�<j!�v�sBf`O�9m�U�bǅ�h<����SOҔ,W\t�|�]8?w�UY��!̶񒗢�I�.cZ��~
s�s��^�kd���1��b��@��@���@�N�3���/\�Ŋ/�����2W>�٪s��ұ��y2�{�7b�>�f����\e9�?��� Ww�Ǯ0J=�&x��5!��FΗӎw�F�y�� �QP[�1�k��` ��]5,:���y�����
�<v����S�t�h����յ� �^��B?����/q�։	/}1h��f'��[b���u��4*�����>�J&�w9���,\� �ƧQ�e��;�ߨ���h(�rB��rr?]!�y��4b~�ã�}m��S1���e�	��p3��*��=ozw���ƌ��k���1_�8'��c�NR;�s��.���B��q�͠�\�|��t� dʰV�Z��ty���*��څ��ЍՄ������S"��1c�{��)�o#(����|��������㴔�
j�	�z����y+����hʽ�Z4�@xx-a���� x�����ôk�2�O���1U�St��^nAe�[��DR��4c�yMs�k�n�&�y��I�u�6Yn�Q��0f�s���<̠Э�5	��:�z��uih4�&#c7S�]��B��쥝�Kt��!ڑ��p�Wx=w�i�I�c�rM{�S�HQ��F:��4����3����>�?o�V1�k9zߩϽյf]�GjEF���w<��DHb��1��+��]kn�9�(L.%:+��k���3{YY#���!oY���f���Ѵn�=�~4���LV��賀u��VUw��/�����i!������W]G}�T����F5R��I>�)��/
n}dO~�Z�-2���~��;^Ym���Q�8�-N[���B��Z�,_�/�:A[��,k�C!�� rF/f��9Qm��SP(��oT{�~X2�T��i ���)�+�)a*�#w/���~bZuȉ�H�ӝۇɼ���t�����c9���p,�Ã@&������竖�����sƒS-��&�����.��g�P��YA���e�ۮ�e�|4��.�0['V?�CX�\�/-MJq����ڇR]�׎�{z�Xdo�1��):fNq��I>��~,+�>��S ��e��R5�S�qse�;ҙ΀�=�݀(��ʳ������v*�eY�%=G;�5A�oǚWl�LS9�rz�Ml��`�қ����9�9]��_q��� v�2���5������H���w�J�������g����? �>���:�Un�����_ҙ�gX^��|�ڷ/ݘܐN�^m�r
�ei��D~k]����E�t��/ѧ	����[�c>�F�eM��%f�X\�nk֤�� 2��5)Ϗ���#=��;�5�4\�#G��?��?�=���W��������|�AK�c��s��Hn..xyӘI�B�9�gYRܷ�������ϱQg�u��������=���<�F��ن�������ڄ��8/-.��n��)�W:^G\�5�:�H�����0�v
yO��)솣���Y&��;��٘��M�8�?ƪ0덻�F�7��/�����^��r�@�hJ�JW�1�&袓���=�1�������N[�*�D�~O|ؿ��>��|�#pl������Qhl��
��!�P>k��6�eC�t��z��9�Z�@�O�N��=ߊLr��ޘ�\���cQJ&�e3I�C�������ZB?>/�!Z�~�����G��
��C����ʀ�2�f}c��� l��`��#�5栐���sx���Ҷڌ��8Z�=~�/�;�����߇��`�ܾW	�[xP�3��V�lK��-{ ;��@񯭯r�w][��O_^L՟3[�1�9n߾�^+y�J
��Sۙo������7:����ϫ	;�Y�Q6���8k�npX��yW�@2����<�5��Ѯe�`i� �[w^w�Uʁ{� ^?��ȹ�im���CVװ�Dl{g��X��Ya� �(c�2Ģ �׮^�ΎP�L��#)�ݻw�D�3���w�`p���1��*�~�٧��,�9�=d��y?�kׯ�7���	 "\Ϛ�oգ��y�~~U_y�-��Eq&{M�./�k����߼������%�qV'�����!t@���{f�u�i��6����~��G����t����am.�56??�Д!��(P�yzy��㮈AZNs׶n-G{��ȟ̆�	r�ݡ��zˁ0�� ���N���̌C�n�MS7z�V
?�~V��۷/͕t�;x�:p�~ڹs'����b?޺��ƖqϷ�"�}��G���늸�3Do���{�=���z�����)6L%�@˅��~������se�:���?�>� �_q������1M1�EyJ�!����+�˺�O+ޝz�b�5��r�ˠIGr��j��m�@ު�8�����P�7�[V �z�����+�4����&��ߴ^�5�3�{ꇁ���,��bFH$_&@{����y���ϸ@���wJ>�`��x2M)�s�B�l�c�
&����x-ih��n�з�M1EBy~���G�yvg�M�ݱ����F�m�>�{i���ͬS4M���R݀Mh����4! I�T|NW�����������7Q`2�M��F���O�cQ���N_�.jG����6�쑵��M���Ά�oZ��ʍ����o�ȍ���50��%�r��5\�]T�0^��Q-'��d,/�l7��Fr�[���H�(�ґ��h�q���=Y��3�(�I��#���	��E��x�k��.�iw'�������X�4"
������t^�0Π��5����ҿ�^�*{B�{��
���}���Q//�z����))3���Q3����Q�r�ʷ�-��7ߤ�?��n�Ww���6G����ty��/r<S��4 I��~��@��k��ܹ3��_�"�GC�<���=�Y&�w��N}������{��:A77�.�;w��,SE�Z�����&��Pv�d����coMw.LyV/~~��ښm�r��  ��IDAT����͎��w���y5��^��:������<D/<�S��ݳ����hW�/f�ᚊ�Dǒ����v�������L#���Ⴜo[9���w,ұ����O<FO>��w����\�P.�l��.�A?�kyF�����F-F��gz=��S�Oq�#�|M-���ǽ�] c�0yUE��E��� ����	�*�5���f�W+b�� Q�e�y��j
 R@�������i�Lj���n�^�
���M[�&���졩��
ѽx�3H̓�����f�u:�b�������&_��^�IZC^�~��;2��]�h�Ӕ^t��։9%�#-'[A��/}��t}k��i\��↲��<��������5ke\R?�3�tRZ�����Hg�=�.�����<�FC��Z��"���	EBZ�՚�����������u�k�1DqX��h�:�T"���۟�ph 6@ɿ�D�b�n`Y�t��(��ER�K#�ue ��Lt�u/B��7�����2ɖ�͆�LGf��3��x���o�+F� �(��t���j�d���L���<gA����7f�FY1X�4�M�݌��9�����h\��ن�?_d�GƄ�B�k��J�r�C���2�\�r�f S9��q>�\ڱĝ�ևbF�~G��/���9�������l����&�������e���1ͥg���e����IgϜ����R�L5M�t��� ��SO=��g=�����ܤE��%e���o��w��\��_�}4��ݤc	��<H%2&�.r�:�}��)�������>Ǟ��?��#1&K��J*��}.8�u����
�ۜR�fvd�}�T����d�t�>����_��;j�3�0� �����|M��G����~�[7�g�I��+�t��v��Ԇ��v{� �۳/��47���zx}2�]{v�D���t-\��瞥�}�=��r�U!�z	��q���[���}{5]c%��	�`Di����>�?�f�B@��0��+�		�}�I�4�aj>EF�u���8��	�Ճ�H�S� ��YS��:�{���<�^������K��+鏱�[�yٌ�g�ըk��ZE���O������xVZ���|�N��I�DB�%k�t��^������3)���)T{'�1�8M4����n��@����,a�r�N�.j�Yٔ�8�
�^`�g�F�y�u@�1k����^��ِ�/�yXL�`���og�(J�"t���E8�8C!H��6�4}��C����KF���۴���K��f*�q�O��g�r�r�qJA�����``ɹQk�U5{̔Z�+��W�Ak{�Q.�po�7�S�������hqNd�8����k���:Gݯ�F���� A�s��Tҿ���ŪqF:5���2��T�W���j�MFdы�O0?�R��(*�� "V�ŵ�2��O[�>������)T(��6��xv����߭���^4}!}a}mU@� �%��a�k�-x��h>�B�ȁ(>�d<����D�X�#'ZЂ5&��z�Ay6Gz3��������c�=N���
�A�r�ρ�ma2�M>��Q�N:;A�u��
���#���ƹs縉��"��_7or�®�{�?LO%�%��EOo*�M(��"�E]Pg�'�oΟ�?���fz}�ɧ,��oh5/��.j�"����?b���c���
�r�P�8�����&�-rs1�o��:�����?|�SE�i�����8 d�__�z��k?�K��'���:��=�%-'�$�2��qa�9��[�8�\�b�Ш��&�+	]�q(G����y_��E(�r��7K���QG7�����϶Us�=�ag����E{��I��1z����_b�=����$k��]Z��`�p��{�:�׷��N/H��j�w�ߗ�7J��������Z��CGQfuH�^�5�!�<�(��O�6��'���X!G v��Ǿ��;��{	�-Xv$�~Gx��w���w�"�H���<���/��/�)�Lo��6�-<�@y�YOieI�UźU�L�A㌪�q�V�w��`�ȴ��,T�xG7>�G����Y����q=Th��G��AC2fIb�%������r�����sb���0� ��j���wc� S�X�I��]�s�g^9Z���!jh�ñ�CH������! ���J�B�d>�$g}�a���@KФ�+^b?�>�S�Y��t�I��b��c���-%��g*�]��z�N��
�ʳ�z�$5��Ja�.*���y�y��$9���	����y�{������k>]#ia�]�1��U:�P[�SYH�6�
�JdĚ8�+D��"2�:-���1�rU�G��&m.Дt$�>R�{�3�� !6x~X[!��pδ��:������܉m7ݵ?�T�@�ף����;�퍇����J'�c8�i�W�fԏ���&�i!�w�x%�S�+���UY@��$-�~�~����⼗e��ێ��7�+mV�1�Bc2ψ�i�:vT��Fްlx:��i��=L�x�f���	;��_3�{1)b �^x�^|�En|0�j�b���AVv�yr���k���ȃ|��Ǆ�&4���Ȟ�t0۷w/=��x�}��$������I��r`��ü�B�����1����i�0ؽp��_�a07�c9�u��I�V���ы����O0V��z��=�@��w��Û=� �ѣG���#ӽ�LzSt�r��)x}�w���[�� �S��f�h>:�p�6#�Ͱ%�l�����r��O�}:f�8����QU�������fG�3��x�A,�(��f!���1#-�6˸w?H�3�<��ࡇ�п0�O28���|��_�H_~u��	�8�,�w1�3��l`�./�Xǲ\H���sgy�c�����CD��g��W_}�^z�Ŵ���EГk�����䵊�~�}�՗���8����>����C,��Y�)r�`<p,��OX`�!bp������my͵�ehƼx�~v��e]m��6;��rXo��q�c�O�B8>��	(�&���3��<[s�y2�,2�@�",��h,(Ώ�|JߋӅd�;v��|�	:~��V�+��^k�pM�"��"� �4絤�"jn�,�ZHZ�1B��ꘅ��}1�C�L�pJ������eS����EŅ]C� ��y��iBn0F�+r�,]����6*�ZI:��7��$$�?��2�$T"Bkތ�'�kx�j�>؅�;��&�:��)7�Z�jLA�-���synm&f,�������.���ӼVcð�X�r�Jz����o|�>��,��
o8��5��U�@}@���B�ߝ@ŕ$�W��L
/��2�`���k���>���R��`�	���Բ�˟e�:OQ��[I�"k�֦��\��;6��P10�i�-��Bo(c�VV�ҩS'�,R��V��݁�]fఎu}���r��岧�vZ��ן��WVR���޵���(��G?J�'��6�8�!NT����go�NL����F���s�I�SI�O(i�T�bɯ��A���z�ɧ������ɧ��.��&���{>��?�d�mW5 FYp�r:�����Po�G( Z]���Z������'K�����D�ǃ��q��Y�0(�����������%����2=��s��Ǔ!�'����C#L���1do��7��Jf���q�d����7)d��=imlJ��i�=h�<�ڔ�#"����$`�1�8����W��ʵg�6�ss�7�}�up��3��si.}�1��bъ��ŋt���́���x�{�]��i'��[�3g9��7D3���\:�\�P���7�|��Y֙��e>iDR^~�e~�#�{E�ɓ_pa�ʵ��j���<���{���ĉ�7�"�V�fͫ4h9����:t��>��c>7����~��Ӕ�cL'��+JA�L�EVk�fK�[,9aA\1��W��G��$�p�#o9E� cD�F���~�V��sҐ�r�+l�����d_b�(��qH���C��^x�����&H�y�:J��as�j��������Ε�cH?q�:�~��M3���MFH���2�ޣk��o�
/�={�<���?�W���d$�Je�����HQ���ң����f��6X��P<�P�q�s�8jΜ�h�}n�z�t�Dc�ȟv��Ƣ�G�[M�]�1��/�T�JD��SY9H-U�\�tQ���lX�8q�nܼ����PV�a��Ϗ�}s�\v���\��Bז�d�k�t^3=0n9����y�􊰡"��3V��7���=��]��zv�
>ԓ�@f}}�L e���*����Q��m�8�9][��@�r�rA��%4�p�Q�ٶ�(j���Ms��Ao����|: �7��O��~��'9�����h���h�2p�D�Q�~��h�Ni��5�l��{ｇ<�Ix��*ϗ_}�~����G�={��܇Qк���mm@��q�%�tP���:�'�x����t/��>����\�7����6��f��87b���� �P��hʀt���Cf9�9�)z����OЏ^}�~�?c�5����Ba�TӳxC��$]0>`<����B��c�$�Y;I21j<3X�~�k̾#�t�e:^%���!lSq�lW����
c��ڛ�����k<���l��l8�3��������i�����s"�)�{M��N�{�ل[^�4xoQ�8L�c�g��O�Fsme�>��c�[t�����@� �l�����ٳt��y�-����&�y���o��F�o���q��ɨ���.�=�O��O�ހT	<�5-Z�4l�b���b�����R��~ ������n^�}��fJ�Q���Jة�¥�YBM���j��pxBq�J��G��>�9o7o�bK |&Y"_$�w9�3ڿ�!��D!4��Op��e�4�ܜH,3#)7Z((1#�!��P?z�[T�}�i:gE�z����N��c�:�����1�EP�%��>������±�u�k�d����h�kAz�h���F^/��³?��J|ͪ��vj^l]��X�?r�l�a��&[�����믳�@���	�!L�)��;�N���8}v.����dUö����~MZ�QEY�ΞQRt��<�2SG�l��\���AP�xx�ԛ��d���ܽ5y�l��CU�/�K�oTz�=�����X-�=-rRx�!� ��hsJ�
>���gT�W��b�s�|Q�S8����78*#,����n���N{�C1
?q?�A�he~���:7v{L�9�p"�>�i!ʿ�$�o�Ѵ�)���T'���4k�,�
��g�~���'?I���z)'����z��x���vm�t�,iY[�:�����}��{��c��3�p��#���g�a���K��Xʞ��70�(�dA�y���Zr��3W�C �8pN�{�!�l|��eaj0/�v��tB^#��7n�ҩS�١�[�a��iBȋ7����?����'i��0wߜ��>��Sz��w�c���5^�^���L��?{i�ݹZ�.�P�����6�wc":|����Y��5�HS�`���Xn�
�x���#]t�O�Z�>R��_y����>G)<�\Kn- +�D2 2a� �iv0��F/����d ��r�a�L�ie�G�O~O2����i����78J��O�C	w ���`Dx�ŗx��[�%^���a�۽|.���Й ��c `��g�����S��o��:B����������s�q��#����^������7���j�s!}K�Ub�8]{8�����k�����%Æ�4�����Q�9�ҳ�y�\1�����4�?��^z9-���Aj�U��5-g�-��6���*��	�����.V���8��*����nV����?p���.�7TP§*���p��*f��[(��b@�v,���w���w��ҿw�7yZ8oεE��͒������U��A����-�F3LE�5��8 K�A[rwe�B%�7,0�JbM}a5�4f ����S����7�Q�JW��Q*�$�n$����d�(�>�z���3����*�����pz�(�����^��As��x-jτv��z��5�#+���	ƹ�Q�aR�|�#A7T:������BI�}��',H���?a��N� �]U�*E���\̌t�8�Q�5Q1�N.��u	���C�0N?��]�1�
�t��s}{8+���:����<�+�����nqQԠJ���Q�0I݁�S�h���1?E�0��4�P�������c�}�!����YV��s(�{�7�
��7��(ߟt�qc���x�@{Rˉ�:L`x~�@���!�0���F�oiV�2�q�}G�Ok�{���C���#v�[��(xR���;�#Js�v�U�K>��9|vO�	�K�荇�L VB�B�o����F�Ɛ������~+}��yk2�M��8�3���~饗� - �^t���oˌ߱���:���5
�	owN��
���c�Nа�%6�"'j=e��wp�rGYH8�í��Ź�� f}M]R���>�M�q��C���&f����1�Α�o�"���z*���	x�汹~�&%���}�xb-0�W��PS<����(4���Ar����w�cق��G},�a��-7p��y:p�.�L��C ]0�ೃ0Цv�&�kI[q���[�:t���pT��,�Z���v~������H�58K����ylm����S]��t=�r����ChD�mM=-��:	��[4�_(Yl�ۍ�A˘i�ֲ�i���aU<����bڈ� �`"q�.+R����j���d�1W��2q��A2�s0M�.��o~ˤڗ�\�*�V"�0 p��E�x��y�+-(p���g�/����t��y�4 ���-����Ώ<���;���ڽkOZ�k\�x��)�Pj���D�F�T�����u�*�Bկ]�X�]|^/�\6�t�Ti1���S�yQM��=[y�t�N̛U144��C�M�F��l�b��� ��m%lgD�/��ą��5cQR�g#�`E�R�<���$�.�VY(�XX��U���j}�X���3Çʫ2��ʴ��/�<�`dg�WBtJj��=�)�0H��ae9�n85�W A;"�n� F���Gi�⁎ݽ�!��%A�:^�sǜ�SFeګ�~}���
��ZӘ#�
�=�����c�9h�<gاF�.���p`�!���v���`mn�4&)��7A�X0 d �|���`(�J�� ( ��(a|�����y��5�9-gM����������暗�ʹJ�S=���i2"��՗�~�����cO޼q����Z��9f��:���w��?�oΝaoW�#�{<f�����/��2׮���){������F�"C������N�Z�\�K�V�<��5���p�h��#'r�����!����y��LGj�#	�����O�4�>��`>Ae=���~~����G}��b����}�p�xÃ�����t��1�V�Eo��-����?�ׯ�����+N� G�
݇�F0&�la�C�x���e�X���yP���������}U*sjO��WI5�kM��YN<O9U��UZ��U?����c.�uz���	�>Ưc��#���2W���^�?��'�D�s"���q�+��(@	�L?��S��㏧��!}�$}��.��<��?�Ȃ)���^��)�0]��@7^�����iM�FF*7�����ۤ�6d��<�uk���r�=�}�){��|u��{���hznȣ�$�]y��W�7��BWe�ӈuHW%�Ƥ�&������LF�n����:���|5�&:��B�Rl��ky*�0��
�, P���{B�����ky7iL�ꪤ' V����m+B�8��%U�x�^H��О����~��:���e��s�������ٻo/�>u���BE�rL�,(ɲy ��c���"l���B�V��������>�sc�8��J�u�נ@7(�'�� |�B�\x�9��V�A1{ǅø�V���U��y)��jY�En-N���AU�0<p��V/�ߒ�%����
٘�
�<���e\�A�z� t}Ȫ���>6�R�f ��Lz�
2w�x�F�BU3"X#�i�Z��~�?,���&{W��@�9�⃾�D��(�b�o���\�V�<���D7�ASO�^�_	�of5��'�ɍF��u�!2��f��y�ה~� ��_����$�l8�?��H���k%�O�U֩x����h������GVj%�3fl]�Ʉ��r [ܻ8Zo���@;ݮ��x���ڸ���Km�Xo��xn���{�ͫ.9���(� �:�(Ɯ@~t�X��t���8@N>�pntGW�4JaN��c�.���-<��!T̺�7��J� x�ۨnu��S}��g�! �PX�$�g��C�!��E�[d�"|���HZ���i��H� Ҳ�u��u����o+����۫����Q����rvS������&���<q�S�Kɿ��Pp]Y_�@��/ �4��s�u�72@^<���kry+�[�5��]�7�␮����z*a��xoޖ�%h,���o�7�����E��q+zH���7R������1~`����e�;XN�2 <�Ff+QU҈�αrm��5x�O�:���N;��_#���܆��āN���w�WB{n�l��$����.�� �t��JM�w���G}��ֵ�;����GԚ��цI]TлϮ}�;�w�/�M�%�8W�	ٛ������dN`���xm�08*������ �P0�L}��x�a� ����|��_�*�1���p�'��O?�4��'?��.l��_���BB�8����eH����1X�������[ZZN�����ᇷ�ސ�F�a�s9`|a�MZ�R@P���i@o��Z�*���<͔	��f�B��l�&C%���Yv/&��kW�e��	���sߛ���E�!�\ɡE�M�e��ߩ|�[YP3pN���$�)�f��SO��]PǠ�\�m�y=Ts��ҕ�}�+��@�Z�0E븧�
��j�\K`��u�MZ�0�N�>��-���>*"cW�BDΓ\{�m|˜��w/Ob�����N��G�d���|] ]P�h#��a���P�˅]D=��ÏvBߑ�5l�n�pS�e�g�w�}����3��G�C��� SH�!�._�N^~�W>X��C����M8�W]�ܛ}~OyB7
�~�gR�dEg�}�݄�����ڄ=�HeV���1�uf�V���N�Ӣ�s;��NA��t	
�v���W�3�9�~��̉ �?r��8X~��_qx��ˬ;a�Ȋ���I���&��7҅ь^엥�C��Y��ǟx��K2@��ԡ�u���%7_�`0��7ǉ8�J7I�|R���3]#2���F�Kbto��œ��O0�mu��b�K.�yMMY����6{�o����G�v�qGx��EZ	���7~���ܹ�˄=0��H�[d6���{�!n&��F�3?����}x�1� �X����>�3�UZM �(Z�@�'���8?X�̱f�p���6�ƺ`�����y�������E�2sm��2=�7��e��۽����u${��5�j1�l�M�n�\xQ'��ߛSʬ����p��&W��ag�<��c�����W�vx� �Сn����wLO�A Vx~�oY�y�$��bx��v�#E�!W�$�/̱G����_x���@���-'c�@�;����C��$�6�lY�c�0�"7<3���y�O���rx�\�2�\0�>�_p��t�V>�)6�h}�m�;�DU~��\�2?�R@��4/���XH�Ņn^�~��$��F�>���?%����V��; �в5��������zx�֓�EN6<Nȃ�����A�h�s�"H��r-���0�)?�V��A70 �`�
I�/$ac���xB���O�u�C���u��B����]����6�\O�t��4�� 9p�+�����9WVD�A���r^�H�P����F�؊�kt��./�:u
v�� F�P!U��d\#|'� I�8��QE-�;�'�h������t{$��k�Q>�<�aES�Z2��|�|Xڞm�G�oo���5�5ew���I�3�sy���
�jV���9�bͱ��Q[�	ە-��s��5.$ڹ��=S�.R��߸��w/��zMUʚ���Jc��3��Z��/�����O���)h�R#�_�>�3Z�t�/
������e t����\�*O�����y���_�U� R�$��7_C�R 9�^�d0}d�
��-r�e/��6�@Z;u�&���1V4��� �>�dR��=ʥNH�f���8x��Or���_����؝v� �=z�oS +`�QK��{�q;]	JJO�K�v!�1;�v��߅3��s\����@� �\� � �p�!}`s����v./16B
&�<}���x�M�7o�~���;n��{����9������.1��E}��h#�@�t,��"&0���Eό�/�a�i<`{�ƀ����i�U�OM������o��8����s�sV��^��5殝������*=X.(V(���:_~u���@R/��2�4%�%(x0�Ǐca��@ �F��DQ�ظ/4�{0��*T���l�����R�i}���Q�@XA��:X�ȥ¹��ĉ�9�	� DF���1^P��� �,�7|��m�뤮��� .[�1�v���D����G]��x�V����EX��o�d�/�B�ʯ��`�7,{3Y�[���\�ٴB��I^){c�h]�vʶv��Rض�*���kmF�X��<�W�\e/".6��CG�s��0���X��QS��p�-a35hr�u�d�Z�Y<}M>��B���A-�V�α7��«lXqQ�P�=S����d62Vf�uĻӣo��gӸ�8��ye+���?�w�v���˚�!P-�fE�AK�����)�>����J�:�zE��*�F�|��Ɗ�db�fP�
]a�(FM?矧����˝;�r��o��fcsv��\H	��w�*���s�.�$9*)	��z�
�J�5�iIW�-U?�T����.�����9ݭ���՜��su���H���N��������CMc�hȣ��c����A�t*�O;v��=��CO=�Dҭ�9-M��~��PrS�?�k��������]���|̏tO�d�h߫k��w�f4���(����ؑN�:��I�5����	Y#����G��Ψ�l����)�L�;9��W���(�Lg����,���� ������z�-:q�ֺ{��g��.��i0��_8���fY_��>���I&����:������ ���}^�t
�5��O?��1��'[!��K�^0���٨�;��	�ac�q�R��y�H#X�K����5�K��;i��Ow�5Ќel�4"��m7�ն�
pA;�ln3��U��(U�L����j�Â�\�#�h<��+(3vqXj��U�^����5��oG��Wk=|�v&����|�>s���}p�c@��+�O?���,HX»w��س
Pk	ߑ��Ĺ�gϞK�yt/HXz�s��[Ƅ���,>7�b�΍X� ���#?��bK*�%�
�{,�Q^��)�	]�Z����L o,Bm�a��dbz�:+�c�L���z��i.-Y����2	K���\��z�$�ׇYe�vN���妲@�$����a#�ZQ��,,n�<�d�\����*�����]�"=��4WH���t5	)�`�~��%�1G����{W��2��	F�U<�!P��dF����%� 0�c��;+��0��O���$D�����\�69R3�q:^�t��~��x��Үt8����x<H�y��A���F@�9��ck�v�ۡx/^��]R"�yw����)P;v�ȼ��Mv,7a�Z��޺E֕����'��p��}'���+���Y0@ s�a���O !Hxu�ք�V��|Ηm��s� ��T>�@�(KtHr������-��S�X�w�[���V�䂭�2$��E5d�Ɏ�@٘!��y�sᅍG���������hn�1s ڢ��
��=�=g���^����s�|ۚ��v�����2�m��ڤ��j�O��4P����*�/x�z�&RY�^������1|N�u���N�^Mp��A�um[��z���IP���h��_y�:���	@�|3P��0��I��O��n	n�p��$$�5g;:Բ-J�Vr�J�n~��1R!���&ٱ#CX��z�\�Fj:k�����=`��pP�N�5�ofxr)�k]^V�Eic�N۾`C�A �`�b*���.�$��{��%v�<�w�Mu�y�)Uo�����,� ?�]�7�|�-ߡ��-�pD�wt�[O��DX�+ׯ��׹x�}���m5�[�E�|�5�h~��ί$<�=ބ|Mϲ/�+�7��"����̳ڈ쎲��O|�Sg"rxv���1ǨL����N9�rYd���V�¹Y��$Њ�HV����1Oh9|�ڼR��
�cg��e� &h�]���O2���	4 <ey� ��|�)����+\��P�p�#t��g�'��z]G̑��� O.�4�U��VtHEx��g���$G��(łXЄmA@Q�����pe�&Q<�	w?���]>`�1���kcij��~���'! ���:ZI
x����T"�|��]˴{�.N^���vȘ�!w-���*�X��C�A��.X
�8�DtPA���9�4'-�
�Ļі���Ȗ�Q�Q<bĹua{_��t*@<��q<'+F� w�|���,��OQS �w�e����OT���B��@E-�0�~�M��g��Ox�1�L�~{�n^��C`<��q����aC�f��20�r!�O�]�xL�xᕚpN���}/	@��G�������,�g+��r*HCu�}�1S3ߴ}���G��ִ!B
��P��c�p��#��xDd.'��s�w���P-�+H�~6��B�mF��=�L��g�^璙F�#�8<�P$��6���\Ph�}�~�%��i&I��B��u����Q0�)ܢ�l�3�-K �Q˝1�Є'�4��=��7�<�jhk���  �X��d�f"�ۍ��K�n84��	�9�#]��%�2��.^���� ��;�پ}���N�0��������5��G��uQ��b6�%�4��6����K��B �y3�وSf��==˥U��<��G���<����e�;����ܜFZIk�m��!�C\��]�J�ka]⼼��k|�:;�V�ϋp.]�F?x�a��C����}��q%�t��
k����\I)@X��&8�N6[9�^P�L�����ר���S�c3��~��X^n~�3fp� ��=���Q��6��uJ&�:��1e)���w��N��b�YDr�m�E,p�,�fi"f�c�#�$���K��so ��?��0�h�P�ej�@����{�2�E�$��p���q׈[u��l2Zn�� �V�cqM���6��,�N���}/�^��V�Q�N�ibG"�0�Rd*]o�։g�Ķ ^�ٚ��O{#D��Lkd���紓a�So��-��v��n#m����q���2���?������,��-f(@C{:T�: ^�#G��W9$x�p��N .�F�|�?~��x�	&����'�������Oq�D���A�\�U�2	/�J�<�T�����"P��!����>M��S� �lq�Dz��
rܧ�k�,|���	�i=��� �S����u��Z�;PO�����}M�<��ϑUφ`yLf�X�q�܀������Z�{�|�©�&���ה��m�L"/P��g-�$�[hʼ9�����6��.��-���]���#Iʥ�%���0%��kb�Q=oytV������5����2�O bJ�"��� ���NI�=l�*d���@U-�	Z�9��Q	� �(֎|�-84��j"�̌s�@B�ˑ��8��0? ��z�<��F0@��d$�LB��hg�{����z��guN�����o����*� �Pd�xWV���>A�caA�D��(a[�wr4n\��m��A�|�T(���bTQ�[mh�|�ȌuS�|ȭ�X�*�1��;���c���@�YC� | ��xއ�:�o�o|��c�zy��
��ͻ��� ���`yȍ/�A��aD"�%�_�����QcO�>@��1� t���9n�-΍���6c�وE�eN�kdM)p~8p��S	��?I���A�,1����o
#t�d}��]���aI�j�zd�x�h7�Qy]x��A�k$
��B�D�j'���,�%h�E�YW��ѩ3�����]us���j~�`bf*],�C�|^+��!(=eG3N���8����p 0�"As�T�ؠ�	������a/-> j�ax^�#����st��Uu2E�*[��߻V��	g~�g��v/��=��3�GЌ0�=��\h�H��%�Ds�����n5jD*[�1'<�� b8���D3��䮋i=���h�����$m�7 ����.�ȕ�,�/	hb��y����X6����VT"~{�"'C���&ϭ%a�񍢅�an:3��1���gl|�]�����Fe}�| ��	:{�k^��<s���L
�6���a�Z #�B�c���h{x�p%�	!$Ƨ�ݼy��'�
�XI�s�'��o_��mx�.$zE\(�X1 m&��dJ�oNSt�UhZ6��^�;Ŕ�P���<��>"v߾�NT�:+�����1V�z(oRk8�uQ{ď9����¬�bY߶��rUul>�S�;����s\UoL
�[��| �����W/j0���2��ll:�:��Ã�.+�Z�A@v��`\�բ㈅g�Z��"����K�˸z�c����Is��F�u��:=��H{���>M ��K�Y�-�}���t�A �keE�Y���3ܢ�E�^�U��eY�i��H��i��	�A.�������/U�4� 0=�Q*����h!�JV�d�.+z��J��$�����d-Y0��e�n�ſ�m]�}��\9ý?�����\�@�k�r��V1���f�����a�/�<���,["Y[S��E7��x7�|F�\�׮%��S�s�=N�A��L��& �L����������79�����4?�|Rf-�fy�#zX!7��X�����F� ��g�ǵ�<G��?ȫ��eYH�k,2ت�}�N5�>M^7�!�4u�u�|�s�J��6T������MO�J���diك�N��Wt��R�>����R��R�'�48B�XR�Q�� ���{.��|��L�u�6�~r��wWY~��⋓P��&�qP�		�4�k�����?�޳˒�<'�i��G�����d�������:�O?af֚�$�>��=:�@� ��i��u���3�#bǉ��Vw��&�Bu]���;"v�u�EF�8���BS��W�W%�H�G�c����;��hW�����D����ι�	�,�c���<�aoU[�Tc!�*u�{���:�T��UG�@%¶����esNs���<����A\+�'��+/�,�o��m�V j�?qL���R�t)��,�z��e��E-���
L�1��|�!��&��_���D,C���W�^|�%�Z��oak'+�V@+@,����4�~���W�� 0K'����2xtWKوf����� U��%Q�,..�c�Xb��&���6���	�L亩d��j'M�EE�	���卅 0@r�a��P�X�z�1c�}���[��\�~F�p���8����m���kaWT�c_����+xW6�u��"��f��������Ѝ���p$�U�X$���Nώ������g�I�N9�E	!u]���fԅ��6ۇ�u����Ď��\{��q'6��&��]։�~�^}��G�d ~��90)���6���c��Jcc���!�\3	f�9T��Yǎ�
�P�̧��d �6�c'�˜_��xd��qj_���{aMm��:�&#+�Ѳ�<�l֮tFk���`���n<�* ����D$�7��Y)~<��m�
('�8��B�D�bɘ�w/{&qNy�4/zs6��9?�y9����G��)��c �P6f������?�q��Vc���8�H�Iȝj�K�Ya�;ؼ�����1՛� ���z��K mV&���}��)��T(dC��*5۾%P���8Ԝ�yž"���Y�˹�w�$�},0��c���^� �Ƴ3��I��X
q�^�j�>U������a��#���Y۱��zRl���Z�.��Q *@տC]�oW�t�����=�x�3����������#�uփ��i�Ki@&I����4�ѕ��������J ��6Ɉ�\���X��&k��1-�0�G�"m�<���۰W��к.����c��`�0-5�$f�	�z�;c0+*m.��t�m�7|fI�f+hd%�#?i.�� �	�$��1���Gʦ
���.\�y晧�o^3����؈:y�n�S��b����;R���׾�����N�!����� }�{��MM4w�$N	�G���`0"���z�c�}̣c54��KlW)�X�eʋ�=�yg����q���Ԣ�&2?���U^r3I����rJ�·�pn$!9�[-=y�1�Jw��r��;�ЌvsG���懞gH��ףD֜mc��;�5�av+�p�M�E�q^���tb��k�@K,�b�vX2���4 Y��$���� �R��"�{���~���/�3�i9��(7mj`o�Y�|̙�uǢ�>3*��7}�>Ƙ?��s�O��M�`��@W�Id�v$�q�� ��X�nf�@>goW�m��|���+�%��:��6K.�������b-:y��{�!��o�~�ony�g�$�T6�Xd�7�/6���oq)y`_�ka;1~�����"��-6�:Z��+3#�9���P�'I�wmZ�7ĘD� � q���kj$�{�Hxð��޽����#��7�mwQڥBC�G�U�dx�{l���[v�
��/W줹ib`�8���0��Y�[:��J��p,$.97�F͜�R�W�<���>��?�QŐ��VW�ġd��cu����󍽕UЋɍ���>i������;u�H���N�o���Z�f�{� ���g����F5�`�e���n1wt�kEVW�pM����eY�D��s�.�ܛ�`
�q�� *@�7�9�[I̜��H�.�8�����a��jX�塦�!qQ���{0�k���G�� ��|�M�6e�X��x�Q�xoW�5#��Nә"Ԩ���r?�HcteO3���-dM6��]�q���֮1�.�!�B�����;Vfm�[�� X#�p�rkar�h��XP�[~4NiG�4,&p�`�%{W��/	�J\?+$,����� ���ᕒ|?��0�`_!������G�(ѩ[�	�`�̻�#���C���K<��c%Y���uzF�=�L��D�q�+@hԷ<h�A:�*��5X^c�s�O�u��.��m���e\f�z��Zb�M6�2dpy���al$י���
��X��	�)8��sX�'�F�gƊ���i����lb�;�_��yC�_Ċ���$�P��RZ��JH�>�孨���-(�f�\b��،�<�%�lu����������%	@�\ǃ�n��J"n�����}x'�lM`_���/'����=]�e@,�,;\hp����7o���d�3	*f����or��';D@<g��������s�y����Y�|�5�I���ȭ�Cm����6�쫾��`Lb��| $?!�k@g8���@�<�Ih�n��+��|-�ɖM'��M�OU㩴�Lܔ� ��N|	��̓ä��qP#��l�ZJ����k�s�"3�"�����~{z��d�>��akK4\Y��:��6����V	�i5'�ssor�`�֣l���32�e!ϋ�C���?�$j	��N�uh��%ĳ�+~�KIԇ������בV,ki�x�$�"�& ���/���>G��<���L�&�'�!��$p�1�����i��M.[AdM�Sk��;�x�������}������7X����BմK/K%G�|Ne.K�.Ξ5C[�i�@���'��4�!��w,�8{*1LP�LD�e%�D�)�%�6/]J��%�����&����H�GR$�������%��kc=C�
� A_�}�{�L�CC�V�%��^-��R�`�#����!����y�(^UHuԅ`B��^�6����]2��Y�.�4cn�3�+�)���|S}O��[�TT��V�͵ʄ-�M� qM�F�V}����f`�	a�����E�;��ӹ�eZ�H4�����7�{՜K/�Kw_��^����n��}~����_�i����w ��ݔ��J�,!u(�fY��l�m��sI*�N	X���ߥgTS�lW�A:5	 �4�,Y��IT��#��s�j@`>���`b^,��%;;�O�[���{�1�-^����%ci�|���ܑ�٢a��Pe�5�G˟fW���Z<�L⠜`�%�(���z�pHwٰ��X{���t�;��K	���r�������8�����q��G�&C���������I�l�W5�t�I(�Ξ�mÂ��M�@IC�,�G���'h�T�Fe��ٺ�Ѕ0D��� ϵ�m�hJl�A/�D)�m��Vܤ��~6�4�=�}��;I�@f��Ĕ
q1�a�U�1|�a��L��� 4�W��z�S"���v�`'�.����r�=���ؽ���k����(�p�������N"-Zϻ�Y�1n+f�(g�̸Gʵ�eib*���x�!\�..c����L�@p@��0eNġ%�A[X�>@���/�+I����>����HL\וI�*Xփ��H?t�����.�q)�$�zn���+G�iN]i�u��U������Fs�K�\�r۸)&KŃ��=#��6��|��W�'o��et�w|=���E��u��.,�|%id
f�� ���"1�Yܘ:��B8����gzH���/D/�����e���~g���,��q�E@I�.���?~��[�-2���+S�i]������y-a��?��p�B �줤~�0�-I='$f��
�?���$�v�;���6f7q8.�%�J5|����[��0!��U�hmq��@��q�@��ǎ�5��B�5J�a `�AG �����CF)��d�%{@�0�nyƵ�X�&"���=�1H�X4o��������i���t�����HT1~��%��w
��p�?l��n"na�E-�D+(�����-�e�sb%�4�}ʔt]o���&#��e8s}mKbav?+�� [�M7+�ΰ!��g���5�"2���Й-��Lpo.?բ<f�^�]�8�� fH����>.�_־�o�@�tg)UԲnb��<$w��V�>��a)7=u��k,$A,V7Oߜޛ��ݵgr�Raqn�C�������܍��Iw�6��L[��mw�Bh���⩘^6X�q'hЄM�Ž�ٚT��ܰ��Wl�� �}ruQ��~e�fuh|�c�OU����zvAVe1��P2(�o�,�K�5��F��b³&$�mm^�B(���~�3i��6�Ռ��̸��|��34��n�CZ-Fa��o ��N��^��0�'Ƙw��w%-$�u�Yt�PA��nX;G?BX���6JG`����@=8 �v�鸳�*�J�>?���^��[��)��/&c�,ND�X�Љ.�����S"EUcd�)��K��O��� $�0��ypq�b������L�8b!��h�PH��3�f�ǃ)-�H��PJ�<-0v��D���|����o��눩�I�k)ZuL�d ^�V���4� ��$��B�������QR����>��7�$�r�e$��㼲�B�[; j���.r� _�
r�dU������!��Eh�1��w����@0��'$�&KO���ڽا�S%%�9�3������n�{##�aE�~4I�q��0�f�q�#���南�S֣֜1���G�[�v�@����O��/�O�?�XHM������Ϝ���]פ/L��jג��g��;}�I�FG!���;$b���bU��L\Ӡ��! l_$�� �_s�c��1ɴ!��M��	���ۺ�xŴ8�~�8h�F6\�T
f�(������t���׼�����N�cLLZ��$���-�	aЙ\��5	��`��dڊ����3�`� ����Y���A�}.a��a�ۗd���� �:U�����?���loonT�X(��e�H�]g��֘�7�ҲYu���թ�K�W���c�a�0g[�����%'���Z�q"U߬Jb�֓��]O�ڨ�l��Tg#+���C�VI<�2(��3(4��גw�:��&�X��U�܀-K��ۛ�D��u]s��03	�=���U��3�v&��P~��>q�������񼩆� ���C���$h���
��h+�?Ң�U�#�J �[@�(F!��٠��ꡯ������/\37�
BT�q��4Ct�j��p��-�b�Z*�o�f�j�ǰ�X�����)	�Xl��Ԣ�k>s���rHxK�F%9A# vP�l�&����/���zZ=sXgk�>��E����@�T�b[�����K�*��U�%q��%�Rɢ��j������SR\�>H���������5t�7'O"�����o�ϩ����g�&Y���'��`$��~��e�x�����}i�b�K�;�qpS�` �1�	�$)��w�]\��˱ʺ�:����kb��|�s��G�bẤ����̭o c<�[��"������w!�dL�0x =u<�)^L?��Ӄ=$/2���A�9,	��8T+�wX3�,e�lN�CT�*c�ßC����h��y qR���@L-CZi`�UA���-�u�7Ѻ�U�0^��I��y�|p�R�P�uM>��W]�ȑ���<�(�낊��9h���k.	2n@1�_�Z�s�Z���8?�?�,��iݚ��T�=�'KK��h�=��,�-����
�+���N:l^;�>���:��@��l�qt7��i�$��̲����v���S��=���J�]��p�Е�"s�5=l�,6�T�g�q��&m�	ۯ�cev����9��_8�xU�;cɈ���1��3e���r���҉�?6��!��u��1����*tï�Ii���2�!��a����'�c�?&U$�I�;�ۡi:��K��h2�Pѐ�jh�$_�V�_�{�:���EZ��K�0\O�g`����J�ljL��"����=ȋ]]� ~���+���\zKrb�������4�с��ބ��R� ���Ύ�,)�I؄�����c`����}�~�jvI��?�0��G?J?��υ���<n���5����o�?r-bג�&;�y��6���>��w�u���3���n��54,h6�0Rw�.(�1�0*�.��d��b�/礀�Q�<:Ub� �7�>$n��<�����ʈ�����亇�FN��FیkSIX��i� ��{%����I���A��u��F������l��W��%�.L��]oN����偀_�����C��SO?%j
��W>x���ꫯ
f���P瞖�E�(��|�M	��:F6���h$��>��t��E"�I�	�p/�I�������	����bWx�WB\�a�P�VȻ��S�|@�T���fͭ�8�e����͔�� S�-sEk��=uI�b�2��j]�0�k{�0�[E�`��eU�/�C�[��Z�h���fx�H���t{�+L_R0_�;3��鰒4k]��h�[�<c~�]��}�h�$ �T(5dm���I�]p������s�3�TLP�6.����J]�n��5��v�谍U�^'�C�������Z�T)0��Z���~���R�W8a4F�l3�]��tLb�Q��d��L�)	 ֲ���:Sgl7����8\�:����D@���ӱxu1|,�k��� @�� �;;S{��iwPmj���g-�M<�#%g�	fu�z��oF34�P��O��G������Ѥ��<]�ڵ�d�cͺgZ��Ae�i<��Y).��m�{����S-Rf`��IՈ/Z�U���sML0�(_���^D�%�hB���,R��L�r�Y�G�ټ�96�|�ei�2�%;X��
qᲒ��,3�����*%��$���u��)U�]�1���f7�]dD)X�+��E	A9�������~T&��%����(� q)^�I�����doh����t ����`��iSnҚ�T� ��[�u�Z�p?������x#��֛�����/v��\��_`�nL���Ӓ�*�����k�V��PH��_F���ߛ�"epl��&a���rҊ,%�x�e���O)�,.)m��(��0ye�^��ӱ�{�_x8Y�Zٸ�����F�18nsL>�߱PI6$�ZO�g����p������X��Z<Pw�u:�}����SO
I�jj.K9�H��&�����6���!������JTX�PF�_6�]�ɐ�C!����N��*
�� � �(#�*��"��0(x d���C�_<6���G|����z�a=�����.XYTB�J�����.q@�Xq�c�U��8֐$��`�.���P[�I����_h�e&W�X�M�R������.������pf�`����_����O���o��W�h�6 QqN���\���2���Nڙ1�p�R9$$��"�A�ǋ8������C�6Z��5f%���A��1�ƽ��ԡ%���Mfƃ��t�T#[<u�f)�8u���6p[p�%�W��k������\kw�Q������	@��$����6���(����r���>e�ؼ�w)���lp�=��/Jx��c|�0��w��~��$�^�N�8�l���=s��.�Ş]�Y������) �زܔ�>������ѶB)e�����k+��@���@1�������d	{:�@�`K��dFǝ]�����e��I�82�I٫x�<~BX�K.	�e����°��+d�����¨���xww�Ɔ�1��Rs��#�)y�p����x����~jg��TAvl �톕iE�)�77����t|a�Jf�6v�F)�w6��M�s�{N��gh�e�X��4I�h�N4��`(��Y�R�Z������6���=��k��c��]"<�,uR�`�������Z��=}�H��|�І:  � W�iE��ЛD�{�\����RF�)�H��h���]3C[R��J�aK�֒ݝ^�����FN�����!H	��]�<"�e�~�}�注t���Eܥ�q��GcW�tVu1�o$�9�@臶��+��g\�s�>78w�H!k��v0e�.��@��	�!c���=}�%��X���T�z�����ள�L6��J,��+fb��ŋ�ӕ��c�?�N����=)=����N��I�Y��=$���ׯ�'��5��w�}'�{�=���0�qO����u�@�
�ΟL��8�_��T���� ������F���p�87^��ȉ�ڄ\)��`Ԣ��d�y�� 6�̠����z��o$Mb-�;u��:]�y]0������jH�Ү�JgĆ��	m�����19�}o� '�P�!�h��OvR�r狢޼����F�_��=�S�,��{��iS:�!�Q��{C(��4.F��%8��i����/���
�M�d�X�͢�ߋXEe`W�`����0��}F'ئ�Z-&�B�1��F�Zٽ� U/E��B-F%���Ut�\��&�3������5�0Q���
HY�8*�\2�0�16d�x��es�ԦٌO���Tb�����u�~M�*����S�ܷ�DO<����w��E�GR宖!�v��R5v
�(k����֊��H2G�̼�.v�-r����U��p��Ұ�*GC&�ج@@X)c��Qc�k,_vw�,�!�76�7�ɼ�c��(��[H�?
�C?�q�&�k}*��˺��g�Fu'=��C�B#���uf�z��0�3�]�;�0�b,ᘎ۝6	l4'�Zp!J�ѕ��y�b��q}2�O�C���:�v�X�X[&0�%E��������ˢFx�1�}��VCi����b����U�1�w*&2k�eg������zkn4w\7���D�������f��e��J0E�)q���z��
��"�C��Mb�-tI��^��<c6�J6� {���T�In@��,�V%�7��$��zt��bX�J�ͩ^��c}٧&1��zfF{�b!c�͜UWc��uz�w ɲ�]3''����5T"䑘m���p��Ҫ�Z=�$���zU��$eg�8%�Ę�)��{ȃ>��d���K.D�С���4�����^K�=�xz��'ӱ�� (�����N���(Tl�>�j�`�����d ���]MC=[�$�?��#"�����-�f�	c�Ʒ��[�_�b:{���o�%e���%��P�d{h	�(VYqZ@�����(��*�{��@���x�̩�{��\+�����d��B%M���+����B��m�ۃ�;���,�vnk�$�d}�as&ص�������Y�.�zJ)��J�����>]p��82/9K�$��q1����qH��Q��6 �	H|8[�{ �` �0��9�b2X�7���Z��ON��Y�t��+O�a >��K,�E�qm]�ԛ��!ѡ��X@�>3v)~�1PB�
Pc�o*�X�A&�Zﻖ苀T�y�˦�[��>�G��^;�O}NZa��L/�_���3��]9s�C��M�W��i#9~���;3�>��Ǐ���^�c��z�8/D_�EN��$J�F�403\K��d�����D��mǌ�k[d���K��䘒6���� �Vo'�'����5F�k�5�kx���>,�>���8Wݟ�`���g֍��í/�>��ε�á�h��@�δ���[�$���1\芥[�7�����!�Fg=b���*F-��.m�J{A����v	*f��޸�\qA� ���ϧ>� ]�tQ�`�&0FS�;.e��
V�����$w[I֬$�h},�/�����ZP�y���\_�&�B	�U,��J8k��߲)K�� �,b熙* �-/mjar��ԅ����c,�mS�9"q]Q����%��v0��^J�S(/GY��<7�M��%>7���0�*chnj[Z�r������WflUo���]`�5	uU��c������~�RLKy�0��ؾ)b!����q�V�)BR���ϯ_�u�kz�?����*��4 �k� ���D�2ǯ���`e���6��-0 )�c�'(��+�/�ju#D����0��,<��7�Q�桠�+@��O>>��	;�t�}��+φ���`tq�(^�`�4j�`w�����~2�=�o����?�������r�)1����-�z&��p�-��y���t$�e��ɛ���YoF'M]��C�֚س��W��8>-���N?�o�%~'��Ԓ�`=^|�E��GyT*!F�,�K�/	���{%� :oj~��ߤ��"
�s�T �@�]��g?'��.*����闿�Ub����Y��T	�M��]D��\�T�Q,յfG���ڞ��i�-��ymG��t'���i���$]�
jV��ٚm�W�@�͂e��ޙ]/ә7cyY7�K�<*Wc)��!�q�� \��-FL?�x+&�͞[m���݅�� v����j���r�����6��lV;{��'8l�2��?̽��=��8�E�?�Q�tTp�͐��8�wQ�g��o��I��~̌�ef�P��J��T���ȵ`��xoʸ�]Z9N���i���6b-�=���@咠���!��>\m�	Ԯ�!kK�ecS�9��"r�~���SU�����4���@�()8���{i�hg������֛o�'�x2�D0]}�9n�Xc��� �L�E�E���}��2Za�pm�@n ���?����>2R��;Ǔ���TM�uR(�}-U�^��;��D-@\B��4��}�C?c�g�j��6o�5��Ǜ�M	B�1b��8�!��g/J�`��˾Ӱ��:��&� ��P,���1%(��4�QI�IBA��'��z�^U��_��&����$M"4b�jCH����!O��0.�(K�kJ������BF�����	���?�0���+�|衳R �o�����8�3aD��^�X-e�!���'��g&��g>���o�F���0��y$��'FKh�=��>��s���3cl9���]�F;�;a���7��5���u?���޹���D�#�wGHA�H��J����:�>sW:5��oO��wߝ��kҖ�=�<�Pڟ����V� �a9�3ݜ^[AE�I�I�ﻰOݑ��eC�A�U��$F�x�+�/`1��M�f~ހF.��Q�� @~��_�t:^�% ��sg�9���n�,ɹs��;�p�q�d������'����������?*%E���Iף���=��}��j���	�=�E�� ��߿`j+�1�sQ�
��5o�1i3��>7��.���-��X�F����&C��5��#���M��&���Y�Vo���n��{d^��:Q�#uL����rCbܯ.���Z�4;I1W
��HP~6�A�(h؂��ho>7����lzm�:yߚd�J�\�ksyEW��ځ,�|3͵q0ѽ~����?��Uw�wV�8�a�E��~n\/���ݫ��#���ce��3�⦝y+$_�`��븯3Ӻ�����6��t�kLr\Rh� g|��
:hrP�q֮�əC��(^��]�8���N͘H��) $�U�g�|6�|��h#lο��/$������?�pS���tw�������p�u5N�I0R�Gu�  T�^�1���5��x�q��B"��2ۅ�)!�lIz˴�Gr��;�si��Fc\����R	&$���+�������@p:��|=�.�ۀ@�'S��q��u<ձ���ͦ�b�Ç�*�I�=�g�R�!h@rA��YT\�;dh�T^ǋ���[�ꑨ�/��
ր!���p�ЧY�nc����+.6��'$Q�]n�i6����^",��_Ԙ}��	׾0�e_p	��e�5ɭ'(����K�q�XV�ѥi}C�+h��^44&���zRXc�1 7	#<d�}�����g��ݑ�ʻ%WJ?�z��q����NxȪ�2�I���k£b�mx�B�uo����c�����%���� 1�xF�G�<����W�YI����/5vo}�����'���-�-\X%>�¤d�i��%=��#�Ƞ�Dqa����O�5�$!d/k���HP��;]���!�^E��3)������}.�����t>Xbt4ӣ�<*Aؘ@�w�kK+��sc �%F�u[e�M*�(�'���{T���ϽN�Gbn,N.��2kG��#��p�����\Ltc�Gd��n9ZӒ`%qYZ'<��|��թG7�=��[�o���Fٙ�P�%��P�{L��=cˢe��O+��̲�d��Ϥ������q���Tr��X���Uө����%y�xX��֌x.xmys�@��封bC�U>3�M�?j�H��:g�X%ރ����],j�K5`�~�6�9�o�[�'Zy�>Z�p����UX��!%X�aX2��4�>��?���B�a;H>���R\ՠ�5~�t:���BW��ۙ�X��$�q�{����	-U�,�	���$����|��FAJr0@P*%6�Y���ф1�+6m�P�����F�{�r-6ጺn��M�!'���B6��Mk������~�iu��|׻w��c�ڲ�y�g!k�"n� !� V��q`^  3�} l΅�gaI
v�M�2ޜu֑��T3mmY[��,�<�b����˿J/��'�m�P�3�G#�m��H=C?����@�ņ�L��iJ������?���SMDC�������� �($�d�E�|��J�U�MCR�6Y����zo�7f䚗��(�x�r�|~̭!�ɍC���{?t�*���/�d�s�}Y�)|�^��cw%�V
D���[o�֫���+��@��mO@�=���V��׿:p�
��c�;��O)�P}��U�;�'���0V@��+W�ف�8�v�>9W�L��:~��b�y�7�Ok�ǉ����*"���o���`z.y�i<�G5'+Z��3�^��&w����J2�9�x�V�A$t"�Yݳ�l(�����.N�5��=�F�L��o�4�{�{_%y&`��j��W>~#}8m�`���	v��� �Y����C�|�_L?ݯ}�k�=|��g�淾!:x�6�2�7$YY���Cv�ed�T{g׉y�f��;N ��t��C��	��x闿��8]�.I���C�k;�H݄����m���3�Z��?�@v&Y�Z9�&�(���lܺ��uj��:�)����<=�5ڪ+G��r<u���1��`�5���;n���-ŝ-p���c�␠� �6"�Cmz˘���ǚm��H�+�Lc���@T�7�n���iE�������Ĳ�*ȅ��X�/�*B}�|�`��3	I�|Ca<4�c�U������ �m޻;�9� p�!�k�f���mF
�w��[������a�kPSl��&�g?�l����i�?=�S"'u֯ߘ���F�r��3������b����ݽ^0�ڪۙ]"?��.ȼݜ�q����v$[%7���y\����D�,6�S'OU#r��N��� ��9"`�Dl-)Z<vx����r���fy��3�Vo� r)�!_��A*�Y�;A����3揞$0D`�B�۷���_�R��?����OJ��u(ƌU9FOd��O1�՘gR�h^��,q\'�� n_��ky��%%;�� �6v�%���>?�'d����P)�by
�hk	a>uͩ��I�Y�>t�����!	I%��;pq���G�������( ��%K�y�M� �,��%v"�o��Iw,��2��`�{����d0��Tz2�[�@��o�>@�h��@���h�C}d4E��ח�����sm1�����K�2�c�5ʤMFdߗyhU�N����~;}�;�I��@���Е8���<!������*_\�u1�Ir̫#	�JB���������-}�K�O?xw��*�W^N����$���i�a�����o��o���u=sׄ��{���|T/uK��*�NS(��A��ϋ|4���B߅i.��
BHGU��w|���uK��]���ƛ�$/cF9�k|W��u��~ph�p����tljW�i�p,6p[�9s�d�>�T9�+,���ۿ��h�����|��p)=���¬����$�]��F,r��+�;m���fM��)�"=��C�o��O�g�>���y2&��˶Ǣ� n�Ǐ=�X����	H�.^�d!�)�$��.O$���5��Kt0�t �w����2 4 n�������E�Z��F�f|'�jٴ$�[�	0�TD{]g������� �f⺕1��R�)u�H��jՀ g<C\؜m��n���D��?S�؉����
�����{���W��ۓ�BK7��
Du�%Ģt����|�r���j6�*Y�:��.�W�oF�W8���� ,�5��U�RN�%��O�M������H�<v��ě�L�Y6�-Q������ �K5!D\�)UO��m����-o���q���d�b�Y�����d�gĕ��K/���OX�
�k\$7��!˲ݒ��k�V'�' ����{�5���8��T�1;���l���x<^�fЎ{�l�r�����3�ڂ�N��X�����h�(�gc�ܶ��t��8H�<�x$c:��Z����lb�")]�K���®���o����.秦��]w)�5F��x�l�L���<��$�-Sfc �!��>�� ���чL���#?x���Ğ ���uO��Z��]���4T�!�K]160���+��ʴ�����Yˑy���C@&��T��َ��3��ހ;}�DŚ�isy�u"- ���$�k��j���b�5Nۤd�1h5!-����.��ĸ36}��&�=�r|����Hΰ�8�54�j��.�xf��o���я~(��/��/��o�2O��E'�
_��W}M��O~2��k�0�g��Ta�9�����|���W����3��֝S����酟�,�ۿ��(>H����02��?�������~�k�?��i]wn�0�&�a�p�I�i�Z��վq�E0�����pXbh�^�΍���r5hI򄒆���ȁ�-�TG{M
�g4�	���E%�-��~6W���7X��vP�7�A��z ��MC�'�ɚE���]t>D�A{L�!^.ߗl�d�B���\N�A��_H�!�����|NbOP ���L  � ��"��;eW����;@�dw��1�����U���2 �F?��#v�,_R��Ǩ�~���r˜2�z���`@�d��L�8���6,ʟ(�ׂV��<��Y_��(�ńߍ���mgzۿ74u�����8���?��/D�.	��k�w�$�7��5�L�"�L@�T���ee�>Χ ~� ~�G%H[�@X��/(�:&�����1@� y�B��)�2]��cH�%�p/��ka�-+H�8����K�5�������rjK�W�OwOF��i^�����	H`��������!������!\C/�%��FI(��u #��)��6o\��ڣR�z�u��O%�B���SOI�"��¾%p����j�D�Ӝ+,˭D�D�=Z�6r$+|�p{�"%���E&���ѓ#�g*ݡ���u����MFP��Q�d��W�6�^��r�4��Lw����z�t?�������Sߜ�BCZPf-ǎ5���(�NƩ�*�y �A���p?\U��J�$`� V�}���e]�a�*uթ�NQ�;�7~��pO���o
�w$�Q5���W ys�����2�q-L����ݕ~�G�����,4e	ƣ�{&��u�𱦨Zⱍ��{�dO\��z$s췬k��i�}�E,�3TC��=��M�{�F+����x�Z"jmxA�`P"aoW�\K��� ��
���O<�`�F6��ӧ��B�9Ƴ�����c��c��/���3�>+^�	.�a轞��_�%���������z�J���K�����s��8���@�DLo�|eP�{��(�"��Z���$>��{�ܻR�����A(�7|5�ޝ!m��}��O�A�n��c�,~��i"EW�YhM�J���x����yyT���K���3��L:;���G[��"dP�s7n<.�{X�X���3�O+�`q����4(>7ݿ��#=���	h.�7:� �ν/�ɰ�K'�4YQ���Z��]��u��`@��ӒxW��RF.M�����5�x�O7n^���"��4�y�����9a������U,�3У��֐W�2�@ωX;�2k��vi���O&,�I%bT�����Yc.�hk.fZ�s�a��Q���ZtS��hA�4�$�>c����0�6Se������׷Y�)Y�krO ?�[2��T�u�MW*�,*��	S;w�Q=L,����V�0�`�� �$n��_1_uH�km��\QЇ;}El�4j���K5(�a�j��M�����㡹I��D*u#
ˑ�l[��	����Z�3 ��@ή(�܍�򓁌���~9]8��ԋG{j��t��)]?���胄_�kn�駾>)}��~L�Ga��f�D��C�e_�o}�&h�PD��TȦ6�=���ge��ƺ��$J"f���1�ȓ���n�;�Ɵ������V��.��\�;�^����b!DrH��Cr�g����Bi�W��i�8v��A:~Y��`�NH����@}�we+Ƶ�7s�ӈ���Q�=�4%��F��h��/���d����|S5M��x��Ǆ,�H��Pّ�z��<c���d�!��&�3ׄ�:\-e�í���}o��_�S��9뛵���m�j%���W��A=�H��{��d��p����0�?Y�a׬����H��AѠ*���94�b�o�wgQ�q�/Y���,����L�~t:Џ�H����gW��$Zډs���đ(�)+8�q� @�!F	��w�+�a`q��(5����g�N/\���v;s�K�ﴎhUH́wpH�޿�^�����N`����z��1�>�|qZ�.�߽�v�ַ�%cr�8�z��+���(E��}d����\(�ѩ�6�����bM{�s�?��̩������@�,,ٗ�mo�`Zo,��>�6.�]\R������XH2e�w���Lϗ�I �O~�ө�R������@NYX�(kw殻��~�3	������](-`q�Φ�;�w��s_zN�`�`�Ǥ��0�����#��$H�3�@G���� �8QdS�I����]-"q�@7(��Ef�eH]�G�&H�`�#��w�K���G��w�+.6Џ�,Lڰ�q�!KZ��n��r�J�� ���8v�l��(��u������qd��ck���p�g=�&P\0Yv9�G���*0?�F�����*thZ�E0zXD`T�,�����n���2Bcqam��2kU��V�r�,ta��8eox֫l��c�F����f��Y媶�y�6�`�t]�X��yX�+M$`6�V&��-�o��-����tsؠO0����_���<�)�����oM�	k�M���#d���KWR���p-hd��ֈg�zp��)	���-X[�)�8 �aaF�'���`'2�Xo����I�0N3p��L���2�(񤺼��V;̱�\�a'cWYޢ�6]!X,����fpY���1�?��mK�(�&�JI3��)�m򁬻/��e�X��y�y0�Y���>v�X����p��^�������{{��m�d,�Zby���NׅA�~�&������V�*Ūj��`�s�1��2�ƞ�j�`�$^�W��&0�^��*n���9���C�p��d���v�k0���̰<���؞��u�a+�z� �����L�Y�E�r�ɼ5j �=ԫ�dP|Ib���E =�>dCӟ���O��^ە��S���p�a��������� ^�@ʚ?O�?��?H��_�şO���o����?�Ξ}D���;��Hrǹ1��c�����R��~�~���nܸ�}�62q�7���?�~�������/�}���$�@ձto���pY5��T
E����"F˛�x �������~���%�a5�%Um��v�n�8nC�z��Oa��&� �<�m�]VϺ�CR��P��,Fڸ�,< ����O^�$�C�/����"��]��*�&'��}�|�:ʴ;�����Ѓ���ɧ���R���E��u?���镗_NN@��{�� x������~f�`�KL1�HJ�XS:�wS�!�6 nڦ�٢����YX7p?|�3ϊ����[oI��w��?E���wlC�lv��ɍ���# W���Q���y׌kۤ�X	�.Y}�3�䌗�Y��>K�e܂ ���_����9..a����}�S�����ą<{!Ƅݪtm�����z&G��r���	g�t(F6GT���W�I��$�j�~�}��>L��4��k�o$��$�.d��avq�2�~�E�V��rlZ|��qZ�����h�j�C��?o�Vvk�а�8�2��$�q,���Lۏ�	��1����"eِ��֛o�D@�5�nw���K1�q4xH	�fa�ך��z��1�uN����ӱY!��J���Iæ6c���S���d�C	y��t��p��OR7��^,&6��i9����N�1ZK��DU7�#��}�HH��|�)�Z��sf���0��o��U
q*��8v�J����0rV(9���t�4�d��xZM���܌C(Om�kU�F�d�2E�}�}��%1k1�����H��QJ��Vj��8~R�8
�#�_���_��E���0���w��@ �P��o���'B���桄k��c�$�n�Q_k��) ��Q��I^ϓ�<��m�Z5|�A��il.L�\7�¸�w�q��
�kYr�g�g� �	I��"�����a��1���^%�!~�	t��F2�u?~��0jT��z�4(�����>fmV�,'*����K/�$�R�_������~�-;� �����0��t^�~��E�9D4�h1ݣj�(���,�@ʉ��������k���yN�:!D$��u洬�BL^�"�O<�{�_���~#À�ǜK�p�|���P�~R��ɼ�"�5V�;�&���8v�ؑ��5�-�Z;<W���������O��iq�,qU`W�y�)�
�
P���~%=��Y�{;�q�P7 �@<,�*� �sQ-��\~�;G+n��c	wֹi����SG�>>��g���t�R.֠�^���ŭ�f���@<�X��*�~�F���{�BCl�N ��;���&�%�xU����l�Af�y���zN��D`[k�������XSc k�&q�b����`���6�8Z��s]Ϻ��&�v]�{�����Tl���l@}��9cNey�@��`SB���$�Z'�ƺm4ebV�uc�.%��C7)<Gجn��k���@̩S0���A3�u�V�5��'��a�"nJ���3����-�HV����!�����7�m1����>1�[���J�FbF�M9� �B�8H�	��P
�fJ��R����\�X.a,d����mq���f~���X[@n���@*a)����=�cY�{���(_r��/��'���,�Ǭ��0_��><�I�V�Nf�����Ǘ�#8�Qɜ���1\��%�;)&�	-1�9K�����S?���i�L}��L[f#�5�uC՛��¬`.��êah8h���)坠/�le)���7��5Ql��Z��јDD�v%^[C+t���\}(�І9!�ܠ�p�B�v�rz�R-~7��X��xtJX�K���L� L;�kvo�8��pa�<X^���W�Ǘ�
��|`�����n>��`q��.ߓ&�=	Е�^|�g��Mz��wd?�f�quxP�sg��,w7bl�I>7x�Q��3���k��le�@
�]e��#�ubx�\�AAW�C�����-NOI�ؗ�*'�r'��`��at�l��6�]'WUI�[d;u$@�12 y���ʊ�{���m[�Y�5�� ����'�T�%�$xm������DEĴ"Ǉ�2n�Z�����+!_r�I���ꌽ/N2�M@ە�����&l�`� �&4�p=`(���ߕ
l;3��lu��][�2e���\���*�F�B`�.禝|�y�c���n0b%�X����`��5�Уq{��$��Ґ��W5 �����w��j�$�/>�����^c4���l4\ {{�>`1p��jk��J���=,} P����/<'�tk�w�xIs���#�c׍�!X!�\��|0X��+����^(�.	u�(�^,Kv3A먃�a�&5v������,���n�n��-���8��>3o��j�#{�E�{ސY�
�$ΰ��X�˄0R�`���ir�;��{�=��� z�ŏ�7������m$�Fk�|up0h� � �I��	�K_�Y�Z�p�0�x(#�k��Iq�c�bH�ρʓ��E�F7-�d��Q}BFF�Fk��=|_���;"m���Fy'<ߙ	�{�}��}��_CtC�:��=wߕΞ}P~� �"�f�ࡗU�X���O�	X�5���q�Z�E�#K2��O6�cd��j��'�PL0@�M��
�;��x��.�=g��eu�UףA����Y]z�i��[_��%c�%g�R��a�`��
麺�g�Ϙ,�u�y�*��Z�*B�������]`��!t>�W������,�	���Z�KS#y�-�{��V*�MٔJ�o�3P������� �y}\X�r�,�oɒ<<Dpx�=�c5�T�j;��i�&�2�T�G̈́g�U�һ\S	���s�2�8�*�'2rH���!/,��=/c�����BV#��B�x/�x���QkW�!Y���n��T@�lwȖ`�g;��/��-�����N�ֶ��!SǏ��:-����O�cer}�1������t��ns���s�[8p_��ϕ��d!NX�J��p/_R�5Y��a�HX�?������4s��(>���2��52��!�1'�I�8&.�6��Q��S�.:�C��:��@�̫H�L��,��Ѹ:Y��}�獂��%��oM���$���7����$�
-ld���/~�s������>-��`�=t�+�ak�lWQz����W�ԋF|�\�| tB$;�U��: �ہ�hɲ�6�JwGb��Wr�[����K�9U�?���BF&�LF��;�;���f��> ko�� J�ԅ��ItXk�& ���`I��	���8�cׇ������ ���5��ܵ��jW*?FI'V�j�@�J�u��u���Z�ԭ�b
�AW��$�c+!ձ���>m���W@\�_��hn�Q��K���"1C��7K�6�f77w���q gY,��dr��^-��X����:�i��iU�=[�Ee��i=I����o�����=���B-�
�I��K�?� 7&/��oh�����h��6�A��TCZ����O m�g�p�T����Y�^ǚV��ٍ��-�=W�sB�ea���ɞ#[�9��A���Tw��m�eԚ��Eþ��0�X�C%D`|u����c����E����� ~�t��g�sӓ%�l湠���ݻ*���Rn0��^[�����ɤ��ϛLAd�
��3*0�6��R��Hy���r~1I�/���P6[po]Q���͸X�#f(��J9��7U�ժ-��G<i;U��p��z���uG�U)F$U�ߺ'�
�J�%'=��0�П�VB��%� ��ɳC�}6j�~v)��~�B&j�
	 �	" ��.W�E=X"�s�q���9�C�ô���*[�D�^�H�ٰ�i4%����n�>(c�R` �bƊuC�٘�k�p���J �+���1!W���}�k���EC�S��F`�;yT6��Fj�����>����~�����ZXD������8��LJO?��F;��{���ШY���Ho�����^�;�M��O�,�u��ڛ���X�žk��Ξ-�Q�̙�TU�}�:�Gˊl,D��{o����펹{1��`��:y��ⓠ�;)8_LR�#�}Qv�q���-��6�P�V7XN�,^h��ի2�D��2�%!U X_�-�r�`o �o�H&�&�iE'��3�8�)�"��b-ie���A�EV���$�$��peY��/,T\��0���%�e�S�'̳�vf$t�̈+�L�d�^36~���J��ɴ�l�H��<b���=�x���kW��x�/u+�������ހ%�����<����fH���
��	#��O���U�dpC��k+�兇hC��tT�_�6�VoNr�ϭs3'�Z�Mucs��c�c�p'n��%���V�L��v�������[�d _a��8y��h�GU'�!i��;��fO�$��kȂBE�e�ļ^�x�>ЛA���,�RBfjhӶ���"2���4���4��\AiC�l���������W|�a_�����ѐnȯЏϭ0ف��)k�p2�NoF���4�����{E��
����tFb̓�u{�M�8���B�����YY7EsvL�̴����0��$�I�Y��+0u�y�⧫��h�H�I�]�
9 �Z�v/����݋�v_v�,w�3��Q�Y&����)sO�|\f�h<"�Z�uކ�ȣ�[o�ٙ�Rºg�H��o蓰a�9���țF�
��>�ի�	�.Ew�(��o|]����+��K�"QnCī��/�+ �+7�4�n���HV��0&:��������KL�s_~N6E,8�{{&5��vlpf(�I��,�AeT	������
����F=f��Q!�v����6�B�`�Z���x{�-~~�IN��vf�б|_��r�l;8�
��`�էH����RY�fu�y��d��}{�s=Ch��G]�Ǯjf��C���;X�\A���x���6������źJ9,G=Cu;��]���1��+s��k2k�H),���Hk�\xgWc��R���P����q��}D�Aw����㎁n����b1�5�s����,H*�g0������9)JK)(pS�Ec�1���u4��j�,6�.ˠ�H�;©L�t��C�u����C~�O��h'�}_� �0e[R�����ɐd��	��z�ʑ+#؅D�\0�G[/$��x6MXa��(-P���c{c�P\L���[�!q�������z�s�� ���yB���)�q�"	j���Ch�?��C��P��L�ð�{�y�%��poS���9��B� щ���A����z�%1^Y�|I�5#�!�%LB��fy� ��O*@p�ޟ1�Ґ,u�o2�:7H!
��n|�����J<&@��mI�=E�����ޞ̥�����iq�h����c���c�2�ܳ��(����}1?$&���M$f�d�d�9�����:[��
�C386����v�&�B]v���p,���*����n��O���P�`=�����T�t�7yW��Ĉ%�8�{� ۊ�c�?�����/�#�nD�ށ����0�ߩXL��}a��<�N\��܃,����^|�E	𗸕-�!%��gu�����6(0|��e��+衆d}f�Z����;���+&\PDXn.d�8�f�����Al�Z���ԘR.f)����i������+m�V^��.t]�+��NI#**��}Ƣ�<��ۮd�/�Yю衝^c��o����
���f�	2�R $e�F�ݣ�Bu�[V�.pY�	�e��WI�zX�,K��/-hN�%[?Q����q�x��ν�~����^���Γhm�[q\ʝvbt�����3ÔlH��~cQ����aeQ��Qǁ�Z�⾞���KyӸ�f(+���P���ߑ�
}�_f�v�h$X5���.0l��k�'�	�������2��>�2�����a�5c�	����H�1��^2o�͊�c#��3��7X| T�U�)8�
ra����t6��Ŗr�ue���A�!�A�{�3=l��Cl��@F�*�6r�
�M+֯�f�g��5>Ҙ� ��ؑdJڿm��]e�2�p��d7�co��v�}����6�0X��t�Ķs�ȩ�tt'�+�~�RNy�9��sg�: ڃ�AW��Ju;`� (�C��w��B֝���GS5�=�*�����7�3�>ە�IK�ˁ!�U�]�׌�[�Q}��ތ���g�Ddف�֊1��ͨ��R�h�{��4�rN���5�D��c5z0�/��;T$���"��̉�Ȟ�`�`�p�޽��(�A`&�����D�KF����^+r��8���WU%7�&7�<[��׋�zm^�aе�	�)	���*�Gv^�-�ÿ��p��)4�D���B���\���	-��ւ���l�I?��=��?�F6�rV��僳!�^���)هj���h�͋��k�]I���k��"�Y$��ޗ���^����������k.4�de��#�/#bj��&
ۋ[�u���4�5nN���Sހn�l��^G��AOtG�f`%&��:�6���5��]Ƴ*=��d�X,�|2�	���m�Pb�v4����U�1.l3zlO��S=�p�k�M����ߐ՚0S��Sx���;�-c�"�9+>!1��2�/Td�9�d�#�(gu���3E�Ži2J^�.p3"��[�L?������ENK�^�F��Rf2�������$5!3�Ϛ7�A�!��A�t�b�_]X8B�M�c���k�۪c�U���Dl�m"d��:}�$�>hy�?�]��"���kȘF�/0�b̬t^�:Ǐ����'uks}��ėeUF3�?��(����k�9g[���k� �����I4b���ۢz
���ή��*7q=�HD���k۫���m���!������r���E��w����y�@��l%����lί8%b����ŏ���`����Q�G]�H��ρnۖ�M_��c�dZ��ȑ��]�dMV����V����]�>���P�{�B�
c�G���P�d�"�[��A��ϸ�p��ge9;��Q� w��'�bhA�1�������9�C��k_G�'1B�Cl{_�R��3RZZn)3=��эS�����ao����{ݩ$E/��;U)c�Frh'�����4d7��?�Z����>����5a�������'�ϰ��~�����t������&c�^9H�/�Ւ;zs�N��H�oq���f8K������A�K�<Z��6�k&)���#��X�-j�V���u�;��(�F�,�Q��mwmϚ���Z�87}'�0&���ھ8\)b������-p�Ə�|���2'�q�$�A#s�̊�~n����}�c�<dL�7���A&���T�ّ�}iC1�V�1dm�q��
��s��h��(�^��-t��
vM��*�%Qv�KW�5V�0�\n�2�W��-ը:��8��1�1֔z��e6e���]�7Q�_7?y��Ć�F�E���;+�����1㱒�#!G�9�h��ދ|h��nL3w7P%9q�	���ۢkN7��T$Z�g�@��sI���2��f��� 𬇖��ޒ=qHV����ڜ����h�I2��f�a��'M"��w���6���h�9o�%hn�l�H�^s�g������M�� ⾀�z���J���������I理�P�܀cƙ��o\+����I"�Fn1Nnݦ��ӣF�{I؆G��ŭ�N�>�Q|���"���-ʹ�H��RO��N;��c�[�0z"^�*�is|�#*U��V7(�.Ciˎުč�������
/��}����8�ϣ��`�N�)N�[un\�(2��F-n�H���Z��
�r�	�z\��մ��G-DE�'�鋪��I6��y��P)�.�ZV:1{g��v}�f[k���͆�zkUԢ���� ���%+��������X���6�Id�f`e��n�,c�	Ҙ�������М��K0�L묗̚g-��j$��sFl�O,�iR���2 W�zu���=)`����g;�����(�� � ���V��E�,˸���60���0�"�{�!k+��x���(�L�����F�� �̮�y��Q^O���K���^n�{ܦ�]�\������m(3 f_�:M�Y��V���k���ߛX9���&�-,�va�#.]�8]�D�j@k;,�����;8 ó��A� ^K+i�N'Oh����_u��4�6��tU����[��������~}t���c9V�4C��-� �HM�3�^���	3�[Y��m.���e��k�ĵmt5�R�2lڏ�Q_�8�s%0�=�	q��
d�,'ϖ��X��q_k�d�}�v�Rɥ����as>��V)0�M"eK�F�$M�?{g�	t��(�q+,r�����f��9R�9Ғr�8A���k��}�V9���D��\��F�c`����{��\���������Z���-�?_�t�v����>���*>�v��{d���tK���٧��Ǹ�i��U��Vv�k���^�j�#&���sQ@wXL{��*hn4z��Y75VxJ�gv(�/W��F7�n��0�l[�ߩ����p���G��&m-��Vl�؎�.-p�}cygѲٙ|���4�_�������؋�~�J�S��0�	��u�$d���yX�n#�!�ƭ��?��EW ��,���
v���vwQc�l!S.����̅.�R��� C�W*S�n#k����hV��yW�C�^kQ.�*k�Z�ۍ�m��vD�vj^�$��쳒9l	D�A���י]�d��Y������#zg�6Ma�qeƓ�5RusP�ƻi3���ђ�:����3���OUd^�9�e[�ZB��{UT�c'���L�)��w%�t�ǾڶN�g�T.��>�dz�����y7���-d�iu��� ���Dô�JC$ ��럔e�A��e3�7&�^�@Vq'N��y���)=S�1�N��.>�Ďr�>��t�>��l|X�U61�Bi�Q������m������3�G:"Ѝc��6�"���(HD�������wq;�Ic�SO״A}h���+Y�؁k�n�4���#����4l���H�I��z�g�\��2)�Y	�y����<��������Ft'�J�����l���dӢ;�:�G]���l��\��A��eLK�ʌcT�u밳���(�R籦�\t��X����$4�݁�4�k��-Q�u�X����c�����Q �����\�6�n�h&;7�z�!0w'���x�0�r3�l����EuvGe>|u� �)`��#�����g��ha`To+�'	o�bQG �G�\�S=_hu3���z��χ�����Ҟf���>�2p�,W*�5�\�A��� ��^:Y��\�H9\I)iXP�V�QHP�d������� Z����㩸�J�nT�A���{��
�A4�9�z��+���$����L���r���J����|�G"L���E�ɡ(�p��ή�:'��/8s�R�c���񟋝c�i��ϡa�i,��[
�u��4Jt\�u�z :�T���s�s��;�}3��U�⒯�vi��c5\K��M����}r���M��،����������ɫ�"�� �l�>��j���� U=_ڸ�ٵ8銽���n��������3���������6�f��ou�����O��}操��k���RS��=C]�L����%��9*��o��Fg�5���T�R�����X7��84>�I�5v�$D�lْ�B���C����ܲU	x�0�J+�������D�$� �@S�����"z���?�Md2�,�<�y�8�o7���׌��q����JN����.�ʩ��|��s�* Y_��7����_;ƒQ�5 ��T����`�pz,V�����-�wTPZ%��tp�")c�+�K['��Ku�1����,��1�[�sj$�?�Ǐ5����S5_��VC%:�L�ѓ6F�W��O�8����c��R�"����	+�*��1���v��C��:�8�kLmY�A���0�0�u#ͭ�������p��ڪ�$6I�ɩi#V��ngnl��Q�Ą�0Sd��k�*��@e��ա���q�u��$o]����/|
1g����/����SE��8�pNJj�1Q�U����d=l<;�Y	;�f��饶7ץή)b���a�p*����H��iqܹ�~ϒ�&�E`DK~n�bA-�.�\�*-��xq�p���z�] ��\���`�TR������)�O�xps�cB'�`X�漞-����Xw�膖?>�8Wj{��Y��͵-�����p�����x?n֛ �A��sĵ�ֆo5�>	Qu�A��nt��npGI�Zq�*j�b>L���(A������z����{��4f܋dZ���!dI�$K�F�-)�P�)ɝ)�`V0�<!��o�c|n�gg�����Pʦ6S�]��׶�e���ݮ^[�|�V4+��zԻ����k�z2	ק����&H�Ha��^tЬ��c`&&7�vq+>(elo�%�W;�is��Ji�n�A�V��7>�!�M�#��
�V���ע���� � ������dW&�O�*K�lݤ��f�
c8�n �8ϥ$(���y�4_P��R��݌��e!LL�*5n�mNZ�$p��m+��oV���ys��䒟�ݰ��~��D[fee���}L���3`�ᰞ6+ޑE�43��`�q�;)�b� �õ�=[L��Z8���Mե/��aY�����ji�G��N:\j�~�s+����'�^K��Z�����x�5����kk3�ݗ^�=�4i���#6��i����T���u�N�ͬ�&�ŵ��j��ތ�o67	��՘�7�ym�s/E�k`U�̖D�%[d��@�{v$ц$�5�d��"����Έma4s��|>���gғ%�7-B��=(��VҘX��qL�N�5�(�l��m���F@��@�Ҷ���m�2����g4��>��v]��<!�u���%�Ξ]��ؾ�:N7��zu����đYd���ڷe3*?>[���ފq�S�{'̩��4h7YS@�l��#���z�vͰߑ�6�<�b�KhkLPz`HR�����J�+^eM^��/f`�wW+]Oe!�L ��z�W�����W�/ަj�JE�EdP{!�\�x�@�I��zmޝگXK�%;v��$U��s��X�n��Yy�������@���aw0�n�� Z�Tߘ_�1E�Nj�`������s��D��\�\1�m[�I0WuT`:��W'bj�]�jhi��&
N-N��b�ʴ�a�LΪq��i�v�or�Nnv���d7<�=k��'H¡��C�5&�V�V����G8E7c�th;c�Mw0%
i��{Q�8�R�������Xh������}1���z�Tf���e�;�}�l{��o�a�[��3�.+>�6���t��'n�+%�$l��n �dCH������y�X$���Y�,��k�E��:��``����}{0�\�LM� y��� l�/����ܼr8��Y�
�o}T�#S�b���e���,�%n���%&_6�F?��b�m
��1�֗�UEk 3Ü��-����B����jx2$���0P�Pco�f���2urwci��=��\��5{b"8���z���>*2��R��D�ޫU	Q���s�>��H ۑ�@u�$!��{
DH�� :zNnp�?�ެK��:���Wf�vv��NJͦ��Z�y��ꜙ���^�sz)��H Hbߪ Ծ���nc�]̮yxDf
JC/$22���ܖk�ݾ�u%6�x*Y�VKۯ�8au�_//��j9_C���&Pc�9qye�6�x�g5O-��8ti �#��FZ��bM��X���.�����le�J���/��Q�$��G��<tQLH���H�2��V�GKj��9�@gߊEQ���u~�B]��	X���:)aY�	[_�Gn�U5s�(����r_C��ݨ��EYXv���������K�Q�:�#�����c!颍Y�K��B�nw�ٷ~�I
sɈ�m��l���slg��7�F.T�7��T��d�}�
M�����$�+�ì[m��́�Q�3�<�yN5YG�� ~�E&��ì�ˁ�jH~hѺ�W43�o$�Ө�#�q\���~��W(< ���U���s��8�x��V�*h_�v�24�²ME�ǿI�����n"�G N&S��w��ד�=�������DY�jC�<�e�ۜ��h ���8�I�JSǞ��t�w���]⹆�-�^���=W�.G�=�^Y����k���=���<z-=g��t��8]�I�W�	q�K.훕�R�����zǨ!sedm����;Ь$rW��� �q��5��@���{�Ym�|]�����D^%��f�.
�S<\ϚfH��Y�h�w�o8�p�D��Dg�ׄW�5gY�	�S�+�p��3l������J �a������/�.fj��W�jo_]��q�~�p͆� o�.��,��n�_8���aM��&+Ұ�>;}�4�9s�Ν;�.���^���]p�c����A�jy�	��B��7nq%2Ь��<��t�ִ0��:3j$Qy��D�F�HTC�Ź6�� /I�A+ڸȌ e�a���|����7�~�!_��vrqԕk�3��(���f����"�ƗWXT?yk;Ctsm�<�cQU\����=�HB_��7���cho�O�>�x��Ղ�%g���Oi[�����*'�.�~\Z��A�qYcw����X�j�bY�@��$�f��
m�����X��7J�斚���ݐG�Jr��Њ�ƙ��t�������M���m����h�X��Q!bݧ��Q(_��U�He�����|.5�e�m	I�6ݖ�Q,6�W����5(�|�J�m'�2�O��HǤq�.��l7�Ǽ����)�����
����kd�	Q3�c����IC��-�P~�������ae9��y�GuG��3O9r��Y��ה�+�[�`/y4ؽ�|�j�h�924����W��P��s��=$����09�_���X݇Cʷ���(�5T��2M��R���_(���`���^���<�jF�����W���W�LYL���Z?�Z}pG^�٫`���~�jac�~��Xc8!�-n[BCv�2�`-�$�@
J?[�t�x�%�v����i�CV|��u׫8v��=N�C7���v�k�ĝ�D/�{_]��9xY<�y �Qp�g����~�.?��S�-��xOP�l�
P�}�.m��VU� �ϟ��Ҁ�{ow�]�v5�G
VE+�5I:�g:&K<��ZI���n��5ZF�Cж\���M1j�&uqR���Y�axC�s���1�
q��v�%'y���r�~o˴��R#�n�*9gJtُLF�fZw|t�
j���z�6>_�{��Lߣ�XDr<�eg9�B�4F*_@�X�F��_pt,~!�Q�h��4��L���i�9{���}z@'66�*2�"[Ym̲����hK㜩,mg{��ݿ���P@@���g��Hg@�4N�[S`g�K4=~��F�8<����W���j���ss��������hI�ΨA�
���G�n;�s��6'UT�E]i�U�lc%Z�I��x�Z:Ѹf��`��ҘI8D�{#�5���ny�f��.�Ju]DW`E����~E-(3�R���%In�R�#����ƨ�䦹Tb(nN�wBъ�,�>�ˍ,|�40�P�Hh��Cα�+H�ڥ]6e�|Y�s���îYd\|��E��X.��כm�"d����r�J/���r~�ރ�f��n}ר�~��\�Ϙ�Y�LN��v
$*n�Xd�`Y�*�;@7&�@��K@����.nٲ�<~P���J?���-p���/�e�w�h�q�m�{�7������5��E�P��=[(ެr�k0dF4ˮ_6H��_�
��s�3>�f;��ĥ�JX�L��s;u䖹R��"rE�,sm��P�J����=���-�Hzm�iv���
�6¥>b������'hsK�߹Ỵ�	V�
-YY]��ݽ���T����b_E��}z��7鷿�-ݼq���b,1���G-�o
����Fy�Y29�c,cY�d
N,{y�X�k����$oO9Y�
M���(8��㍍��k=�1�EK����,��9P�'���l}�-�E���ro(Ŀ���7���s�U��g>�m����ƽ�.t��?L�Ս�BՈ��.h{+����<ad$�b!���*&]��'�^���ۿIg��_���ܺI/��"}��o����=��h�D��hp��	����2�ݦ;I��r��o,ԋ/r����5QX�8��j]��,��xc� 3Pv}�4�F3�[8�ŗZt��i��?9��R��2�a�����\�-��zmy�%�=�B��$/}�e�I�F��]P�%u!���®:��{��T�kBd�>�d���cN�����o�AL��qOk�k��&�� l8<�<	J���J?fq��Pv�P�w�]��}�%Jqߤ�wn��d�<|H׮^�~�s.3_��:��HL�\Wxx�"��#���2�8�8����8���;�W�=2m���ZNk�Y��;�^�I-������q�T���v��������=UF�B�{t�SF'']l��-�aHYᦉT��Ჴoq+���X�$dC����&���g*Lqp���=��c�TYd�g56�E����Q�G=a�f��+��w�r�k��؏�)"DK.��=��z��O�Nٖð�h�|(�����ߚDk�g�]_=&'W��H��m�
�{���6h;���F��7A����+h�L��Ƨ�g�ғO<���V�`���m����d-�N�<ŗ��=�q��t�}�~����1��"�X�i�Hc����K owg��_�iIb�Q:����<w����[t��IƯ�(�����7��'��v��0��twZͻ���3	i�MsgW�C�$���XjG�R�Ƒ>�%�u̧	�d��nJ>A]*�	�� @��I`�+1Z,���Ѣ��4*�
˅)*�g�E����R��+�Eƙ2}�e��|�U�aqV�+k�yk+���f�-�V���w�|IO�`�nWu��P%��9ˆ���V7r�7{6�i�4NzJϴ�&�/�Ȗ�����e�t�rZXg�b��B�$G�|������>[�B=���pc �ܿw?W3��K�jL��H���L��B�`t��s����-����]�V�E��,�v����X�]t����Ֆ������W�LB�1*��i�ﺍK�n��1:��*��(E	�jpL�-d�9q$�<F��Rrp�AS
���4'&�� ���8h�d�%���7`%`�Brk�d�(�^|G���4g�%��.޷�~�n'P}��M����&-$T�w���K�:��g.Ԗl��_ˁc��������_ߡH��X-]���y��O=�~�8E����0�7s�f�հ�Ȕs=R�m�Y�U_˖�����}�Yr�%�z�z#ɴXN�fnr��=��xE�������!�sm�ު;tN�����Z.>��}�Ћ���<P�\��Ԑ<7Z4*�L�����]�`�䔻�W�=��! ��K��%�/����#�d�v���3�t�b�'���{�
"pq(-�3ҽʼ�H��!a_���g&�k�=�@����C��d�B��JX�" �w'����c1<�H�y���&��ij�*�a�@�p���, �Ѯ��kx�ʘy�]י"i�����}KQ� ��>ga��};��'4nd-/--i�O���y)4~��*H�Oᡯq A�Sm��=�g�B6�e�a�,-��N�`d������'q�L�	�=����oq���z-��k����f���L��L�-�#[{ͪk׆p�����9.Wj:�7؉�Mv�BA0�CĮ�m�me��D���s��01�+g1���jJ	�����c��3�)�1���%[�f]\�Rŋ�u��-�y=B)h�&}�:?�Pu1+a*��Y�'��X�Job�e%�+��Ҭl���sf3��k?�D���`��@g�޶��nn����F�nŖZ��hx�)�-�����Re�]���'�RW�I�.?���ƍ���^����
E
��{ �ˢ��:1[�Y!�Ѕ�b���aG��G��ek3h<�)��ܯx�E��+����]�Y�ܪco�c�R�������9^�.����e,�<���8x@k�*�vSzC����OY�ǘ���w�
ݛ�r���V����c��y�|I(�?c��z*SbcO��k��*��V��,�[�撱������PhK��ʞ�F�1�r��7,u.�"Ι�a��K? �ʕ�0b�7Ş�}���ۜ`l���,s�}�+52Yd��*���	c������9��ݿ�+q�������;m��*�O(+w�<�'���?��d7�_�^����l�3�A!k�1'7",��d󩖬h��(����RV*�e`*0�
[�Vцd��mh�l�9T�;��\aE���!OԒ݆�t6�a�'2<�=����⽪[�cBw����Y�Oѳ�Ԉ~�_Z��ǈ�w�P��-T��"W+KD,�h��g��2 �L���)������	���4i���w�k�8���,��`�)�+�y�*On#+\��)���r��F�QT'���b�![��Vr�lta1��[k[/ʙ�6O��rf|}[�@؍��,X-x��=,Մ�m!�6�ς��9�x��h�9��⬬�7�������s_���y�0�{��	�D���y�Y��/�[1`[[[�ӟ���a�#X{�> ^�R	�����tDTە0�O9�1�K����o�Ƞ�%�Xy۲6o���g����y�2���/%˱�\�@^�Pb^c��V�����I�GS�f?���
�-;\����.���E�{�G��a��缯6��_���}�������S[� |H�����Ӿ������:+�,�e�y&պoa��ks�A����9{���uU+�hy�?��J�z1ϣYz�&�� 4ِ�#{	��r�6b5���9� �!oa}�a��`�@8�打4݇>A�O�����}]�y\MloB['7isk�V�e���a|�����}Ր��fTr}�1m��)�[�_'�~~��;�1.��!�z>ۂ�b)F��.�m�u�('殮��}���c�E��k�
������h�9_�3Gc�Vo9���d��ͮ)�p��TXQ�C����L�s�o㑔sK��Z�����fnܵ��(Es۶�؆bR�Q�i���vv�-�Ɯ�����iX�pN몞XFpP��-;�~�N�4,�5D��Z�,������.���?d.�x�"� -]�!��b���sߧz#�]o��}���`�.�lU�k}�}��\}�mO���Tv��z&����h�˿9P�1M�P�ӝ��x�����D7��ɨm�Ra�&|�J��d탖/��ܻ{�v�wؒ�X5� ww�G��! ��爿�>���'��\�z,��*W�S���cf����:$�[��{��˦����6a�q�V۔q�Nǂ齔E���!}?�v�
�ݣjR߸U��7xH�q�rǉ\�%M�b��`:���Qd��u�|(���?JJ��O}^��!�4���:��p_�BkS�M~[��%�b}7Kǈ��%I֮-@��ļ��__��z�6�ָ|�?z�V{�-�4�7�߭nE��P���
7���-���xU��z�=���W�S �{��˼���R����o�����n�� �np��ү�X�ܲ����k;M u���:{�s'���<��3/rIle�{]���u� x�E8��=���wۨR�Dj��ْ?p]�ۢmZy�q��0����#��-	nLk��rO[���J�C�=瑨�ʔ,� /w�����(���"�l�|��"�m-�kVi���(�X��u��Ӏ�Odǵ�*M`�l�lp�,d�ru�b�$X@٭G�ȸ��v\�@�N� �c	���Y�b�e�����F�&�o�>��Z�-X?[�Q+�l�����$�~�T�Y�L�W֮viȸ�IA�M�}щ�i�b-j3��TH9�
x�.�A/*�\-�A�cnc(՟J�L���Sk6I�<�)K�a���1HOIwx�-wA�[���B�[���l���8��`��Q<��7Ial��?�*BW2��~mjR��F����vv�[p�h92�0�䬛Q-M�r�UW�M���8
x�1)�� A����#r
�)�QP���l9w��I�u�8\��.	k�"R,��D���q��]�O��m�G��+��s��n`�we�?'Ӭ��_<`/f��l���],z���df�Y �o]��=�ni���c�\��{���<I��,{V%�,���gf'����DY)w�(S��g��`�(^3�`��Ί��pp}H����cݟsrT�/՗;���ؚ�>C��H�R`��s��dY����ëջ�9�n7��x�}�3��U�"WWhwo'�����~����7���2�m��n�v��Խ�d�%���j���g>�}��
���$�a�IB�0}X�r1���lx���/�^����� a��v;��ֲĕ��9�!//�0Yٍy_Ęj�5�HѮE��P�g͓
����4��{���������j��AS`�X� ���h�ev��g�����:Y�2	:Lbv[�:*u�C>�U���7�P�Y�i��)�l%T�b{ ֱ��>�����.v+ ��-c�,���-rLpה�C@���4I4k���F= ��fh�9��Pm�?�<���u����mWN�2�]kV��{6j�2u{�kum�鳑nR,4#��~��Ä�������Y(�:�%�eg�ڝ?!�s��-^N%��ZQ;����I��с ���59���Svz�����}�$e���k[��l��u����ѭ��{��s��Cx9��0�譿�m9��:7EI���DO3*�%f#�S��%Q)WL��u��2�9��]�cIj�X�.:��Y
3@F��eE���O��[��X�A���ِ��D�\�d�=
�ute��ʳc�|��y�ڢ�&�rBeVNC)����W��1�����"h�ǲ����6ԟEv��|�xњQ�*6m�T��P�@�3����j�o��G.^��~B���.���,��BF��~]�߫���D��w̓	<��D��r�6_7�(kH���QaOЂD�˖��G�f�!b��h�+���.w�0��|�����-�
�Dc��
:~\:���5��|�l��Y�����%���m��ew��ﵕe��p�n��V��;��/�k�FAY�;殔��12�6�F΁��x�+R�c:��+�J	uM)����;
�ҡ��jbʛt�a@�+*���\U�Qo��Z�[�bl:������>AC)|<���x�hő�	���G׬����T_S,��������;j�=��63��YU����0��Z���p�~0q�u��|��~�cc�h�1Ѭa.�`͹�>[zM8�6�I@����'-���PZ����Y�����󋕼����(�q�Vyμ���m1�Q=`6��9Rp o����Z�&�'�0�����@��A薱����"n}"��Q�4������
�U�G~��M&�4��*6p���%�8�wVbط�<�@���V~q|�
xS��⯣6t���;��C�/�՛�Ra�������v�J0��T¾x� ���ӡk�� �d	em�<6o��o��TIW�y�`M�yQ��M��?��xT��1�T�,yY�"��Y���`,7��7�ě�owjY��h��Ȁ���pO��s����� �k+k��$r����*�욒?�U>WF�2Ҥ5�?�������V�x�p���Q%��ȃEb}}Ġ�(����Y�_ws�Q=�-����a��A3�y��a�K�Jt��`'\�����뢣vi�	Jdր����$	�X��F�3�R �p@�._aM�qCUE#�6�&% ���ksG�����������[H�m��Z����}mQ����{G��#����UG}��(|G��6c�A3Ϳ�l\�E\���`#{������K�̰��������O��?�>�۶�rQU��nMu>���ǜH9���)�3�=��s7��l����=IeX@�7�C�m��ԤF�'�V��h�F��{�M��/��̬�rHr�R�c���Ҹ����`�d�����џ�ìP��C��0�n�zl�s�-n�&��2�*ܦ� z�%P%�?V;缙 *}������:w{�=��A��:������x���+S[�z�VQ-�V�G���Y,nr>��Zⶽ�O��v@�,@wn�t����j����z>t�ր9�bWeM���rY��"�.b.�Kʋ����rX�SZ���0&;?,�[:C�¼�
:�'py��=���.�Ѹ���wW,�1�K�saF�P�-kb[g�s��Y�٠���59�� H�����3i���Յn�̽#�1T���[������e���o.C�x�U��}wQ��JR��Pl������y?#H�1u�ƫ�n�ii�,ȴ_�`]��FY0�;���.��2�Ǩm�0����8N�,�V���_�ō5��||��b����n�Տ����BSe@n��#�}w�g ,��� �����9:�9�<RGjY�q���\�>��y��JX�%�W�SA���������>38�:s�����~�;��?������?���T[[��X�^�3�us����r1�P@���P}��E���M�@��w�PV��R�B�kȉ�M�X�HJ�*E���3��'��Ov�I@�ɞ�T�"ʱ�Cm7<@��O�Δ��;�d>#k.���w��)�������wap9��'٧��R�f�}߬�ރ�f��x��X-X#� =p1��*�g�����Ʈ���1"��<�8�|�^�@����^�!Ej��������{(�Jf�g�Ӈ�V9����>E�>B��A��0��d��{����F��Hc_G��+�!D�^<$�?��?�<��r�X�m^���l�l.��p��}WV��a�kGh��ʽR��,�F^W�i3W.{c`	�~U���1��q;�<�
�]\?�9c'2�0�2�fj@e�&3��?L��w��E$N�ⷸL^���w�&=T�\�D�f�OH�C��.��SO=�U�^y�e�T�����j��H�;3i?\!�\@4�D�$ӂ=�����}h��آ�l֝�]y��+���{߷�3�?�)Y�m�1�Bw���������8��'L{d�P@!5C@:����˗y�"�
�EI̟��'<��߾}�+��
��x�̳d�]�ԣ\@!�ی�.�\$c�X��:aW}|t��*G
w�Yt�uEx;��Ʒ�v���
=��3t��Y�Nrbg'�۽}�L����чл�C7o���~Y拉9��e���O�pI����N}��7�+����qv�s�B�.��c�\�JUt_�tC�U:�}-��\�M�〤6��UΊ۲K�ٞ�yݑLJ�r)�F�+�,m�EbNT�3��|��Ma[�4�bԋ���F�p�e��� �o���5j�

�
�z�/�\�q����fHMY1�c�H�g��>͛}w֤�C�H<l�[^b�O_��7���˘�a�������`�<�V}��}T���w������r	��!����/sI~,' �E=H����B�+��Y/U�SSx�|��PJ���!�n�+᩿b���h,ah)'hH��hCV]���-k��nV�u��T ������������^�=�ܳt�:V2��~�NP:���j$��ݨ�SM�[`,�Ξ�<bT}�XIl�D��9�'�i�DfO�>���<�浲�`���q�,�0�mӺ|��������l�e�	T�ľ�U�>k�<^�$o����#��3?�	��ӳ`���Y9�%�����s����E�m��3g�0W�_~A���/h'	��ʫ����6[{�S�ҵ��F�9uX_�8W�ۂ�p��LrY��8���]*+�~4��s�S2�G� �B��9�A�|,-	w$�@�V6��8�I/��2���?b��/��N�;w������>_�S'������H���*��W���>�$mwe����b��MdH1l�M�r+͢pEa�n���GS]�����[��'�zs�$����[tҿ�����`�l����z���V9E��ƭ
Wp��q`7.��?L4A�'�B�#sV)-��̷J�������?���}�
�Ep�Ӳ�����u�2�{#0��=�\�%?$H���:O��u��{m�d�i����⬘j�EC�t��k=���Ƹ�<�y;��%n��C�z[��`󆜑岹�zG!'�� \ �>e��j��cn�݇�Y�5����k�2���:T)�!99��|O󤗊�mV�-d��CpҴ2Ewx���&%�IeI�b��U����h�V�Q�p;О�&b��e$�t�{�l���2�lyCC� �A��?#�@��.VO�/�j���T�dw%�O%SZx�$t��p`W�C�"��<L[ML�JU�/=A�\qE��y��i� 6H���W]��Q��K����3����=ik�����>�u��;3�FE�Cʄ]`���W�����]4�{+�����y�N��E2�ս�8!6��]����F��M�k gn^�4�� Y�늋�HV?,�8}���?�#}y�:��x�~���ѥK�BjY�ٵ�7����a�z��=V�?���l�j��Bl�]�1􋬺ޛRl�1�aIPRǁ; �@�d������
m?�f	�	�:S?7t��ez��K\��死�Uvpq����4b��K/��dȈnݺM���M��&m��N§e]fW�6��t{����®Q�W����毚!�� #�ʣۨs@�d��j�6V����Ś]� `PY�)�g�gv�ڋ���YCU�fx�@H�c`ן7�����~1���C��I«��Y���-�e^�ua,@9	�	����R��N�س\�RP�|�%-;/�}����_9�3��������yD��NF�`XS�&KC�t᷄Cjyf9$m'�7�+�*���-e�7���`wn~e��1�[�1_��Y'Q_C�I"�Tʗ'�ʸűs�-4T,[��F�Z��)����Θ+��d��r޷�(�F(�� fJ��玲���tF&_�fGA����O>a�rA�y�˛���Ө�xAu󵻬�+g�T�wd#�{G��/|:��n��a�,p˂����F�˱���m�����,�{��j��[ˆ[W;�\ڐ)���R�e����� v��8kL�j�9��:�,uq�mм/��y�:n_|��Q��У��a������IJ��E������2��<�	�~��'��Ј{����,�`�a��cs�ǨcN��Sq���j'��V������}��!pC��lP"��La]h94�DH��ʚ~g�>��*}��'��k�������w�ZQi��:��^��i�m��Sc��Z�W7<�s\����9�Қ�hc�(Q��T�wa�Е�ZH�{Ϩ	y[�y�ޣ������!c-1�, ���������K(Qً`|��H��O��~4�����=B�+g�{�ۑe�_�Rz�fej�	�S���j�c��79܁�� 	�m��\t0p�a�ji7�j��e���U6��`}��K�:=�=�qS�7ʖ^oN���:!��2�
Ce��We��Ȧ:δE54�k�'l�Ҝ�z���08��&�ZHO�+�]�"����c��� ��X�L�`���F|0���������!/SLn4Ɨnq�Ø��'���0�&�ƀx�Y@��&w﮵��vƱg�F�,w�|'��*���lD5�\)�I�:��ϬæՖ�پ�X�Bb�?[g�j�	��-h^F�I��>KiI$c̬L��X�D3˪����~������S]�|��~�G~���%?c �M����|�1���Pz�zC������z� ��n�J��C�V���yeu��O��q�nS�aHf5x�^�9fs���Y�S�@��bI|��쵘z��o?�!�Q��q?�I|��f	��L�9}�Û�'	s�^M�!~�a��]:��J�\I�I�M#u����	LW?�F;I� ����0�JTJ��r1�j�_ Y�7���"sU7F.Oe��ȹ�)�$�}k��F��9U/��F�4e�g̿��M�O���β빼}���.{O�d�3�0uҴ�Mvo2�9>�V��Td�L���ٴ��В*��NBD��94Fm=}�m���.�,/�ߘ�H~D�NVk5�E�vZ#����ұunqܼu3ͽ�������0Ũ@�7NlqW�5����b-VE��s$�a�˫�^]�'?���}�	{,�d@���͊�
H�ʧt���IX����ίx���VU��8�y��K���)��Ξ�ɿ�r���X"��J8����x�\Um�<	R�����/j�^nD
��I����`9����OT*���t����݌��mRd���_N�2h委Z������T��L/Vjd�`�X5�lڃ]#�7S���3�1Ӑ�{Z�8�MZ���q;^�3�LL���.�0�1�tOC3�����h��l��Q?�c������y�O�_�}�R>[��98Nj\bs��^� w��a�DfZ��I�ۊ�/*@��X_�`~{��z��Bu�H�:i�ypz�3�4T9D��?�u�b
����`M2��=�<��V >�W�z�+��ބn߹˱�xJ���zP<nߺN7o~�\�+��Y�ئ�c�	(C2�
G�{O�sK�Sz`��9a�ytȪ&r�v���V(�Ǣ#(�����+8����=w��<��|��"G#9&*ƁP����9�O�YU�#�w�o^�v�>��#����:&�,�٬(*У�����B�$k<�V����ߞ@?��/�HO?�'��"��~�`	k�`�}�=T�2z6;��"�\��Q�f��jip0
���{��_��>��c���ݠhp�C�$K�J	*�\�	���?���2��!���M�Mw����FX�t�k�7���^��uTydEZ��3�u��׌_���M�{,|_�<?�+���������`�@��R�Yqep�;d��k��~6 ]�De��T������x�!u\��օAP=�J�G���=:��nt�sO��Ѫ
iÓ�\����C�I��8�&h�W���%��E_�,���� ݪ��Rlm���9T��EV/�������M|N|hT�}5Q�*9|SqI����v�?�<��&��@q��|����v���L\{`ˤ��Y����gs����<�ʞ�"0�k���r1���g޷w��mVP\c-�,iH>;u�43X,/�����[×�/������d���,N�O&�,��(Pqf�L�|�<��-��)���um�-�ý�[���l�`���M־F��wV�T�O�26�Wnәwd%$�*�m[s�����?���������l�e��f�6��ۏ���^;8�G`���7��-��?������k��?j��p�0r�B" �苧�~�^�u���k��w���
��F"�q�X�Xn�&6���	��ZpU	T�@�ٳg�L��q�(}�9�����ڎ�6�}�]ȌdF��=tdS����{�徉C� �]�|6ŠG��7����j���=����2E�U���=
�9�V0�g��X�Q�^'iWQ�x�r#I��In8d�.i񉐽�P�vҿ�d?�%��ے{K��.|׳�x#gv��C�J���-�@��-֔J�TI0��4[ˌ�%߹�?�5I����[|3�� ��n�.(�	��w�\g��t%۰i�ͼm#��eK;'�aM���b��>X��E[Y��s��\�V�\�!I�ׁ�=��l���c�r�1��~��`o��|t�\?�مf����������T�Ɓ�4'_�����{u�0|��V��r��Q�$7�"��E�6��iY��(���7����ˀ.�hg{G������U���,j�a�v�<̪maT�2!�<;����$�V�g�$�uJ�s�:&��p����'6Np_�mlЩJOnm�e�3�jp/�$�'{�p���/ғO>E�Ο��4>x�3X,5�D��v�S���UY;#$��8&1tP�A�q//,�k�9����$�~6��~QvT� �N�+�Wz.p�=%�&Sg�`�10˃��W%I���j���I��yP�mG��M�$r�k��������jl=6%�f.�:#e�X�O>��>��#	?k�U�A^���ɦd1���I2��w���Zig��Y�c�����(���փ�]M{���OЕ+/��|�~������}���X{�NߟN3k���d+��Re5�>��!7�{�
��l?|���մ�~��~�r_50��%��l�K5r�+u��N�<�י�+�=�-��-�-�Ej%���J/˖�ZQ����#7�����v��4F@sٛRFQK��ڐ����K1���b��~�s�ː+���7�Zs� \e���GI�L{��k'lK��Y���(τD�.�L ��n���u�a$��}O�� ��%��lʊ_W@y'kNt 5��xl�'*w��MP���D�����㺇u)@�']}��yp����-��h�@�7����l�c��v&ǵ�յ�<݄m�*$}[!�! B4s�2D�U: k�+�҉T���78����nY n�y�U��h��/�Al�qh�Y�E��H�ģ����ཹmy�v���ea���M5�믵��W9Ǹ4%V�$��G���H�e7�T2p ,��k����[1	��'��ხ�GúT)����� (���ʯ{�%�L7�
[��)���{V�c�'A̸K����B����n�u�kF|�xtB�;9�K���d�1������<��U�[�$��d��ebuW�UW�F�4Ѧ����pp_�e|�6i��S�y_�h,{_��"b���C6����<��X�-� S&X�uc[][�{ܺ}�~�ϿT�K� r� ���5�+ܿ_��3�\V��~���&�"i�����w�p?6���'�D�i��쵟��!M|���H�.t\R�x��Qp�"v��]���ϓ�s���� J���&q[�U5c����E��{)�G[O�<� �{��^���䩓�&Ia���l9��d���;�y�\�,�7�5�ly��e�X�x�������ڞ,�� �0v��o,�Y����`u�!���H^���F�bW�~ �5VYPץȱ������d��-��~�Қ@��kw
�,,�uA��3OQu��*�&iI��k��-�Ṡ}�\�>�9M�jL�ҙ�'\o-a�ڇ�	��ggt�h|���t*�.tw5dq-a���b��Z�x�����B"l��Iw�1&�����(��koq��#<?y�y�gA������A��<��'O��B"Ġ']��-u�;=��p����H���q�~���p|��� ���g���/��)��1C�Nض�R����1���{��N]Cp�q)W⏭���,�h����JPB�� aY�]ns�)W<[Y\�H��)'��o��7O��	�nn��xJ��I?�����Ȗ��Ρ���{���Ͽ���-q�遄$p�����\��K.����x. 孓[������	��9�0JYb��mLE���
f�~1��S8f4<�U̔({�o,�Y�	[I�"��V�����o���X![�ң���H�t� ��F"ָY�d�f$<�(� ��ˉ]K��6����HLjK�v$�G-[R�f^E���Q�S(��{�2���x��M���D���gt3���{�P8���'����qA�a�$�n��w����ԟ��3�Nѓ(��̳<wNln��e��l�����ź\�Q�
�W�{2��nD��;���Qe��K�Ԃ=����Ou�y��1LC׍�w�P���+5�����_<o�J�k	o�*��|���od�mS�1����\��X[g�W�r���'�����n!8E&e��/��F�/bN�&����~��!S�f��-�Z��L;B�Y�\#֖k�˦e!�V��M5 nUP�������%}X	N���������o�l8R�Ƒ=W��ϱjHjs?Z�Q�͌�u\P{��J@�g�|��yo:-���q �Gu�G������<O����A�Xk�N�)�' �9���FU�S~���C�-m��yO�N��<_�0�W���ە�y� ��XN�<���I��{��I:u�4�F��϶�k�s���w����g���ϰl�\ݘBPZB	1�u���t��-�9�}�6�I?� �V��r��Q���N�N�`�|�{'�˕�Z��������b�=-�[��.�rpO��p�/v��83~ ���;��̝t�i�z��������ŝ%g�c�d��]����J�-�ׇ�mm��0������o�]Sp��dI��V�MumN,�����S܁�\)�g��X��Z���մ��Wҩ���L �" ���:I�a@ٌ���H�0�y�Y$)k�?�|�F�3A��\��.��V����ӟ@�EP�:�V�=v6tVtv�P��d�C�	�2���X�?����Gup��x�����'���~gļ�9��(AuӺ/�j
"���)�
q(���@��<��(lH�6���%t\�`���D��
�����S���წZf��KV`����+*a��݆��M�����X;'���	]��+
��	�7.�ۮ�&9�J��|��dѪm8+�6�h\��I ��B՝b���~iDs�F��'�t��eJ@��ʟ�J�vP���#��#�����,=�hR��CE�X�Ɵ2����˯�޽���:��p��1��X��P�ʇ�����C�����\l�`؝쓬K�ĩ��a�����w�����J���5�Z��ĀE'���3���� b�Z�PbyE�"���S����@�846�3N���s���W^�
tW^x&�N�[�u|�
�S�1X�a� ^���t��u��6���.��.-�y� �A�������w �!�܆KL_rP^}V*q��{)�`�m2ѹz�mK��k��bu�e��&����20HAX�YQ`�[3�?�5� #�3 ]�//�A���VY�q9(��[b'�jV�c��\,J�Y���]�n^#�Д�fЌp?hܹn�y�b�"��k* D�E�H��i���~�
�ųؕ0'�*�ωAu�A�b�̅�a��!��G��l��yH(�w�����Q���β�� >��&ޛ;�AԶ�p-n��r:��lNs����0�\�:'�74o�Ve���]~C�����ү����ƾH��>[/}�%�-7JǢUv�=����N��L����l�5�mmUw�,���M���l�c��@lׯ&�5�����%���`��Ɨ�Et��]GàA���C���B"�6�Ԋ�)Vh� ��@31��%�#<�f Cȋ1μ;���#ξD��W�������0����X^{��̑9��Ђ������!gq"��@��%�b���[�S��R6e�w���A��O�uvIv5��v��Fj2��Y��&���	<N8�#j��:�יV,$��PD��`�k|���HD;{�mn& �,qu4���x��~Ǳ�h*,���E3��/��?�w��#}~�=xp�?�yc���}c���Ϟ9��F�6����,�# �B�e^�d����9G�Y�_�q���Oq4���i�/���J'6<��,ai�5��f��%���$AỰfw�c�������שּׁ}�~C�VW�����B��uk���IX�yT�.-�r���k;���N��Q���8����5� �vQ�5��B._���#�����8�A�p�ʠ�E�!s����1�����m\�[Q$�ĭ�}���6,�%'V�����y��(���g��%���\���N�H�7H���icy�������~��,29%�(F�����1�n�O}�@�%;�M�^�����mc�{}�
<#2�ݫ�%)+,s�p��C����TX���z7/}P,��Q�i�1賆��]��8�l:���OkS6N�oBp���T@6�(,����Y�3ǁ�ю���L��b��X#�cdnNa�*�i�*1�\��<^�I8�&�=W��9g��H3 d��ATo}�c����7��M���n5;�%��`̗��QY��l�شƣ�x�,��͎r� N{{t��-Vܘ�34�(�gÆ�X�)S��"�z������l�ZQd*�Ƣ�P$�iM���� �W^|��|�I�����[t��m�[d��1�S飍����lu�]Ĥ]�|�^|�%z���ܹsp�?�r����M� v�d��t_	��J���&�����駞���}B�|�}��Gt��M>���7KI֜�:Ͳ�݀�|��L	�a�[5ْ)!�R�8}wii)SU�^�	b�xiXλ   ��IDAT�G�JY-[s��R���`_!�E0 �p���!����{�{��Ѳ+�#��]`�w��=V�Ο?���s�Pf��Z=A��[��]�z�CF�[5(ھ&�M�R�.?Q,� ��#���}�N?�P�ₕ}Ȍ+���y�4c������~����|�����/ҥ4wA�����:����|��}ڛH<2�Gz>�p��w��a*��0�C���2���!�zO�ə͂);Q��N�
j
��os�������ư���M�����3�]����k ;��%Lq��e�u?��q���ZV�홐PU����T��%1�����5/ب	�����o$�!�@&?�p��d

�5�j"چ�[�!��~�����s�> n"/~�z�gQBPŏ=�Y[KKdN�o�,�X��jV^U��/sr�}(8rξk��И���Me�/�[9����$Ʉ��b�kKL���7�Ԧ`���r�����V��劊��ݨ@V��u�yp�% :��R%V1���F��.���
79m1����Y��uJ`G8�g_��G�~����E�l�m�6��#	ё��= @㿵��d�����#�4�a����l�I�l�����_t;��%��qP��1f�|�l�(E_� �t��:�~��6����������?�D2d��'�p�n	P�Z���K��瞧o��-�ǅ�,d��?�f�<[9{֟���II|��X�kl%~"��?��t��MI�ڗ�����֍�MZ�x�!�&ՙ%�$���Fi��焑�C�lgl�\J̕��t'"�@�u���5F����5�Qɟ�FdO1]��C�_��g�}��|�I� xgR=�ԓ�����=�ޥ�;��N�:��d��� 	����`�h$@�-�	䍵�{%{��?8ɻ��}E���� �$��%z��cU@?A!:w�,���k̽���gy�a�������C9�~�+m�ZJ{-��%]'�����N���N	�qµ(8F'��k+���o�-��h	\���N���ok�KX_�ߞ�S��Y���<C��^~��*W�v��?˞�ߎO�WL�ʣ>�C�u�1��[)����A��浨��S��9�%�C�/=@����<�4�^�(�+ʪɦڃ&c�h[��qc�[Y�(�W��rV8|��������<���ӟ�yt4�1�:���o={N���s��u���N��������7��V�����d4~��I�(Y�B���RM���-Y����g58?G�{+�g��lE��r��d�z����/�r,K�:����ln+-�d����!�������f��:_���hW5����!ł��I?���M�p�6�"�����������+���q��y���Ho��f���a��2N��/_�W_}�� ��V�BZ��g�<D��d �[��4��=yr��,�`&�er��C�!�K �w���V){�>n��b`W8��}Zf�"��e���	���h��}��ٸ
T���q<���-�S�B�9�_�bxV��~���x�ﳳw@ۻBQfe�����/����/����ֈl�vN���Ɩ9G��ot�;�~jc�C���ޤ����_�r�~��ҥ˗X)� ���BѺ|���Ϯ}���m�(9�f�Bn�f-3E�	��KV"\P�	Ϫ�le@�2��g_�JL�����j�����O���l�
��U��޲��-��"DH�1�rh,v����t�%�d��Ƭ�b���Vy�)1�W�����X�z*��&�ˏqܶ�-l4��GĀK��:�q�B�)�3��8a��J�h�d^��@L�ιƍ�=œ��:���ϸ��	o~<�x��v��Y�S_�2QhV��}rY��( �W7�.t�22���uYS�����l�� �i��YJ붢M���׵:�uI`"K��ۅ��1s�l��gY4>�(a�"��9kӂk��`�W�jEN�0v�Th��mnd�r,h�������?��?��s���O�a0t{r;aq7s��,��l��q��  ;��,h��5k�.`̊w�}���P�����N���(���l]��/��>��cv����k	䂈��^��,��5��C�s�K6$�i�VZ��U��1�l���@���Н�wx�X[[I��D�p�8�b/N�*J�e�K�(�rVԗ� ��S ht�GC-�j-����>�#���B�"�C �ӧO����D�M��݃���H��-��ܻǮx�����C��0���.�Ųu�����_s[^ku6n��R��eϲ�Jb�-|bfs�.�o�aw����"�ΝU�� ]
�x��VZ��t��Iy�T���������Uc���T���<�U�Ǜ�.2�=��0���(/)I�_^�����*g�1�'���Cԓb��%#Fw�Zikf��C�Ƭ�4o��E�#��*}+k�|�O�5ك"1k��:fb1��&sKB��J���?K~c�e{�=�T��1+EgN�b��^�*����?xp�nݾɡ2w�ޥ��{���I���v�_B�Aw0����+q�:�o7sBx��Q�$���WP�w���f4ߙ�����VH�y�j�n�(�'-�Q2*e��M�E>�؋�0f�s��Q�$���ml4�AF�ɥ��襗^`�0T����{檡չł��4�|<�1_�*J��:,�ߋ��@nf�`Q5�Lb����i����<�����U���>M���k�R��g�3�c6�F��#�r�Ta��Y�`Ĕ�Vx<�gϜ�غO>��vv�X��5��w$�!����~#��]�/����O��^�[t��9����-���8�Ymx�v"��/rmcʫ��h/,� n`�x��$p�%�%BNn��;�n�ƕeHG���mnm�3,���e8�
a��=hp���v�o-Ob�$���c�~�,���`�G�P*`������ �l3�^�{��f���X�.>�_��}����F�8I���~nepg{��h�/���ۗ�t^�z���s�A�M��`�x��wߡ�	�"�sa@X�J��b�����*5�����[	1��q<�0bU5+z{�=��FXZ[����%��vo]=��Uğ_�y�1��QS��<�m�5h 4��f�,�*S:�p	 �Tc�5��]��Y�e�is��!_��rL���!0]�dũ��ܯ$n��Z�g��c���q:ͩg�y:)���s	�^�t�����|���=��SL}������rB���O_|�y�zC�gU%�Vƀe4��>,��^�yȡM��bv}�Nq��e�+�[��$�63��X�U&z��s�Q����P߂P�����6&Nl���9n�����e�X`��<���bw�7R�v:���{Ҫg*��B@���^7��	��/hAuρ���'�\e�G=o�%��{ϻ��gH����Ÿ��po�ԲT�׌ێrav��?�|���ɛ���M���/��kx��w�K�{�9./��@�`�& |?m�H��U�����&1M���8�B,�w��a��s�k
�%C�fW�p��<X(Ο��eZa�#�7x��?��*`�xz�;o�W�𵄲�͖7�m��ݾT� ɏJ��"J�e�4�M\���ThIm�X��/���mvm���l�y�7��jGZJX�T)���3��]�:I��#)�k��� �R׾�Ia�~�K�)�~c��፮�i�\��V�S�i  �]���վ�E��Ϯr<��;w%�ay���a��� �ᙡ�ݺ}�v��@�#�*;��CK��Cf���3Ğ-B�����B�V��'Z�P��Z��}�T��(�M &j��k����� �a�G�TCſ��l�o/\��I���t"����Di���r�+U��?�)=!�S�q���róھ��~��󈆄mn[e�-
�7�	�i��_������ق(����/�̬k:��IN�}Fh�"�j�7zO�n7v4c3�Iz�X���M%���-�2O!w(���M�{n8|�(�������1�"�'	r���I�ܹ3	�^ay��3�2��2��E^D�#?w6�̓�t�{��E���5�x �0�X�D���U3PP_D��"@:�0�Tx��g՟
���f{����=����O�7�5�5}V:�ޮ7��fakZsO�7O�k��&.:>i�!	���Jz��Ez��g�駞�ӧϰ�A?4#������z���|�8�x�,vo��{��X���u�a����<�w�{�GŌ3߫�q�@��9%"���?��S���<:�d�	�Ǐ��6�U��Epl%v!��/��$쮼�=���u�TVw�~;{;�����Y���-�X�~��_ӛ��&Ǒ���aZ���5���_n��l�-O�G���:Y�b=-�$��qiX�@�K=ܾ��K��ַ�;�~#�z�ͷ�_�x�&{�\]
	l`Kx�'X�c��dX9�b��a	A��<�\�Đ�H�����9�I�	���0����x�^~�e#����_��A�`��A��I�Q���X�ǰ���G?b��+�1!C���"�=+��lڪ,�X͍)�a<�Mq���~.��r���_���{I����6}��u������f+/�9����
'!
������������9gyi���
q�%���T�CM:ٸ��i�/�Ҥ ��6�$��K�'_a�(��*���3uvXb ,p��1����
��׾`����d�b}����W^y�.\8Ǳ�/��"}��5�ʤg=���}��<VŽ�s�gU�ݕ�)i��`������R
P�P�IR�|��I��
��N�&�<cb��Q�,�����{XOX�´r����n[!)5>�B%��ۘB�2��Ɓ~��68�L	c~=�Fl��Ē��������$o;V���EQ�<�=9\+H,1��$e(�]�`���c��-XN��nR��H
UG/��]L�ccc�� �X(���Xy��\]]���~;����\��)I�e|�h�s+\�6���ٷb)��1cѠ�=|��d�+~���lT�{��a��O
���A�B<���N��s;`�Gp@���Aًa4QM4f���ƚ�r�@��'�L?O�SO=E�?w%	�g��s��lӗ_���2��Y[��=GQ
�M�p��C���,?3���aW>"8���y8���|N{��g�ZU���_���,�F�c=�7s�m��t�ڏx^J������!�1fP�8;=�����-��Y�c���/����W_�w�}���w�J|��.X�Z ���\�'+��jL�?�������{DU�'�|:���;��.��7����s����^z��`�1x+l�X4�?Sv��`xz�X�9�_���eh3����1 αu�V����<�	���Q �������� ��\�3)"��e�t�>o0��O�ϝ����?���H]���E�X-;���VoP�r�
 �p�Y5_�g-lcj� �l�gF�޵��~���o�F�s�ao$��=���_����;iLau���e1�T1r�ك�2�xF�,��!@Oy ���X�K���
��C�a�ACI�����1��Z^�,�k����>�����x%p ���7��g��HW���F!G�*ssy��thNMWx��a.�����c��n�|e�� JY�T͡�e� �ОW��f�Ky���K�%���%sv����q9(��@��Zǹ߻�k�@��a���ۺ0/�R*]�;�0;m��č2W8B�0� ��.�s�>'t��$Y
 /�����O~��o�;�Gqy>�;l�E��s�ES�����q�5�cE�Sj؜{�_�}`�8���;���5�-�P�A�;�>̩�\�po�b�x��o�s�=�,aВ�ױ�@�A��%[l��՗��wm�]tx�1���vd�M�q��n6���
rݖ� ض�p\�@	�P`�6Ũ�J�"���P�*��Ud�߸q=�=���ǡן�u�M����{��3I`w����W虤�޻�~���3�����cniG��}���1Ғ�� �:k1r�ީ���d������6=�����_�N���P�j�.JX.!�� �NXܙ�)ɭ�U�x`�Ҏ�;w���7����x�ч�7���b�5��m�n�9e1���1��͐�R�iB���b�d��������6�2����K����Ŝ�ؼ�@��z�!���{����������U�;̸��G��8���?��B
�+���Ly�ci�KA����Ǳ�!O~0��o��*���u3�Lz��A@'`L�%��߿�}���gN�ϔ���P�ǲ��9���3�K��������T���6*�|-kl���#E���w�a��Qc~E��P��B5X��莅�y4zl2P��a��%l(䤴L7�!���[��c���䳇R~�@�Cx�Uo$Udp;�䵴WQf]Y����*�m$�~��5�qF����䡅YX�5+pd��Ϡϕ��6+T����'O��:0�ov����c��y.C��m:�8J9H� ��*�?w�]�o��]z��e�H����O��_2�����D���yn>����:��q7`�w� r�^�[��? ?�Eq�ѷ���>v���j�����^q�A8�q�@�E.�=������j�5 ��� wkk�~��� �7��5[3��T�BS+ԏ��򫯈��K����u�G���t��t���g?��X��ِh0�� =��  `�0E����[ɄFGxq��j�e���g�.6�	� g��� ���̔`�vKӋq�Nɼ��y��g8�	�������Jjߚ�}���w���{�C0M���?g���xw��b6NM��}�n/�Y�)�Pq�h�0���N��qM�4#1�(�����}Ij�g���gΝ���u�"��A�P�H}�+'~���aFx�[����7�ރi)�[��
��"��XC�_J���u��	VYLB��U��Ժ۟��l���q�;i魷ߦK�.�X��y���"�n��s��^P���Ξᶈ�7d��ow˱�Ϊ�h�z�ƞ�t�=,�˔O?�j��W|4�
 }�x�!М��q���<j��6
62J8e�c^��ל�(�����<G�|OF��`"I�P���,;0ƶ�a�*pQ�_l-Yr)�$���ڢ��V��N�F���P�D+�e�]��T1w�Q��%|iʱN����K���#k�Pˮ	�҈���{���	�mp�&��~z��K3i��By�p=�����]\���G�}l(}�h��q�n[#��w;�:h�y<*Q���<{�^�������i;��`<_]b�({}Rw7'�� �-�Yx�ZO.ͪE���nrKD l��"�U6J�_���Ҁ58M@JX���hx%\��<=���C�v�*}�� Pt��5��u� ��nE�E��\��2���!��T�SVs'*5�F�D��V�!�`��w�~$��xe7}�H*���b�p-PL�� ���o�bk*�3��#�����8a�pq�%�&��J�h�ek͵[{ �^�hr�j|.6ۦ��mFX�I,(��S�����������$U��-.}Aݩ�O�f`�Xoԕ�kK�C߀>�|����������޻�s(gç����h�l�LNƲ���:�
G�O��3��[�I�m=�V>�e��� �7ml9�?�����4�81��?���P����E_�@?�Ko�L,6'���S���yt}��m�b���7�5���?�{�z���߇��<��4p�#߷���9��y7�鷥􍜃
�X/�X#_����&V��2�����Ȭ(���$�6V�v���"
� ���_�u���s&�%	�sD+&�=sxP��S�.U��������쒔�� ����E3ع��kA����e!��ehë�xz�Qζ���]&J�0��B�r�,|�2�W��B�#�k��P���'��W_y�3O�<��j��JԜd��hY2�5��A�� L�f�e���]C��W�u���.����~T�����8�A������s��,� [b��XTPR�2�Ș��V�}0�IX�l�	.X��A����u$0��0��;�#�N�=�
��9(�ս�h%����cm�XHu��Pa��3�LN`�wޡO>�������~�` ؂t�L���G׈䶒�H���3���*j�\5^�+�@�G�Ĩ�5��d�1�p�,A_4M��4~^��v�Ν;��v1����[�U�հ[w��=�u�ĳ	8��g�I�ؤ��rG<�%�D+&1�b���I?����V��Ӊ�xH�	S)��̓�b�K}�c�mX�ʀM��k�6�#^��ߑΦ�y){$b�GJ��2;�9&�!SSb�pI��!+�5���zVr���qBL�x��ٕ�E^k�/EI����H{�+�_�o\簅O���֥����Tz_�YT\K����!�ซō��׺�Tn[c������[��MŬZ6���=��c^nEv��cx�V���8�]����7Ԙ��z��Y�'߷kZ�:^�����x��5.�1�8�eW�qF��b,���'���Y���;b��CV�'	�p���Y?̂��%E����t�����S����2��f�!c���ꗽ4��P�.�R�m:�9^�>~�*�LyPX:�i�b��r�'��/��K-��e�@���F@�.�z� mOH*����<o*A�%E�1"n�4 ЧO��W^~�-�����Ӊ&Z���	a=��h5��`�����Q�ƶ-�4�h�7�Wq�X�l_O�U���,�q�>���"�}���X,*�c�{��\��(�J�����&Ѵ���J	,w�⊔��ZX9Ϟ;��8s��-�}][����^����!�zP�0�'���Urҗ�]�'�1[ia3Њ�6�o��M9�If-[�c2��3ѸOq7G��~bC�����u��n[R2Q0w��b2f��ע��eֹs��AC'��Q���B��7���]��������r���?��j|��t��=�ߐ]�(�ce�;�Kbf����c�	��Xg-S��J�v9T���8e)C�� V\�����'p��m��-��N̻�>]�n&5H������+)��}��8E�f���Xxps"_��̮��6��Q,��C�>��R�je�ʊ%�fXÈ�F2���ǰ���.�oP�׍=k�(���={`$�d)��-a���0���.~km�M��O�񂠶:<��/�{G��>��P���g��v��F�Rr#�|3���|�By��ʥ�S�����Ic�;�t�-3:�u1n����EV��J����`weu�Ä��f�W&�3tH�"��x�������C����Zĕ�>��On����{����}���"���%���)��5�J���p�C��!�]
��jp�\3���[Ius���L���sZ/ j�-I
m��}�>W��ܦ�V�YTG�r�Rs�5I�c17�RL0�;�����5m�f����iz�)�r<�� �M��� ��]se�D�ذw0��E���̆f��!7���?�U���ו�U���P0�-,|�#��wKԆF	�wx]��F�񏙸��̀�xI�j�)v�RR?��*ݾ{���J2�7���)�Ȩ)��6_[�X۰l���@zĈT��6���2?B9�Z8x���*��(����?
�qmV˭��f��x�y9ǚc�� �N�>��pPZ�*�p�W��?$� ��o%�pȿ��eN`�	r�IBA�'���8Ҭ����l��o�#L��B_l~qM�HF�x�e�"�c��+c���>��o��@���v�u�w0���P�|�v���af��<���䞷��^a	��k��b���Yt"ƪK_�y�&�l`�*�M�I��%QXr�N�g�o[����r=��à��l�����9n��u�*Vo�M��ɣ+�3w�Ef�����B�f�9����aknILR�7�lf�bLB��^��D���ޚ2T�h���&
�O^L7�1���a��q]�t������֠D;������RG�,�����eͲ+����Z�$p����B������`�t0����dHwl���ed0.;�Ė�%v���2m�
E<��s���^g� �{�1��40�pp�t>�L��&p�I	��CM�sB�G6����#fB>�4��6��i���\����f��?*D�T�q����.b$��x]G�<J� �m�߫�+��5�gc��Ĳ��䄂tG�ﾔ@"���*e�7�x�?�,;\��[gzhE#YﳷK+�l�� ��C~R����4xxwk��x~�oV�1�vjEI�s��>�[��k@2N��>X�qSv,���a�LQŲ�7�ӂ�n���V@�M`la|������^���}/�xw6�(���mX������cG�zs�Rk�$�L�Z��1������u��h�YIh4Lͼ������x==7��A�������F�*��ڨ�f�V�
Ed��>j��,Ơ����5���)^�r}`@ܾ���t��6�X�#4��C��
����<Uf+J���k�e�{�h~���Y��k��d�����n��o�_�ޫK�#;��!Rg��U�* �lrg�9|��r�av�����_����<3l��P� Kk�U�E���
3s��̪B5��dTD����ٵ�~W��Zs��Zgy\[�AZt�p��e@�Ԃ)�Z���0�y�3���^�<�ܘ��(]Z�2���0�>���E���YV��
�f�����|��F�j���dZ�����O�Q^���j�TNK�:�_�u���i'�&��IC@�a���)e����S�}<6O�3�ٯ'~X����� &�^��.ZZ�w�}�#v�:|�n޼IV�Sn��e��?��\[�
��y��z��e�����i��p���H�2J>ѝ� T4�tYPZ�!�_p��q�������ߍ���y~`��C��*�i�G���[�ִ���$:`s�c!�,l�[��o��K@�tZ�����p	���u?aa�p^�t�nߺMW�^ew�d�P �ofQ��G?�!�G��vK�8��4?.��qP���w�-N9v��I6����Ki�v!�,�0��aƦ����-H쯪�����ml��:Z|�I���!� o�j���={��U��̎J�5���ųB�����Ħnl�����ʶ8g}3cd�w����@��s5;�]��������� ح����|݈)�����_���o�V�`l̮��0���3OJ{I���H��e��O�YNY��\�I�ifX�$^p��S�}���t��i���*A�`X�{�>�ϲ����3�b��"��`]���L�����̉�z��_ă�F����UmR\@�w�N���m�y+�����<1��b�*��@dbJ]�����}�>)`?(і�N��,m�g��Y.R#k�L2\$���.��!G�رC ��g�_�A�PdwIE���6:	'�����a�ndi�8���K��������z�͆�.n�Zل�N\���L���@�_���ѣ�\>O@���՟�9����}��,�9�����_����E Pɛ�{��AFNQ��>��H�隚���%A6���		�+�ư�4@�iu_(��V�US���|��	���~�-�!ȿ�!˃�5a�<��Ede�9���1�l��b0lnJX�++��^��5��b� 0�,:}����G}Lϖl����:,bΗ�� � �L���*��t&���3��)�H�eƈ�W��s\-���K��֞o�ˁ�㜙����J.K˃i����h�������lE�.�����\1���S�X����__a���]�L�.���� Ǐ�|�o��� ���pK�X�JM�5�>?(L�Ơ9�
�fs���'��&�>f٭�E�TvD�E�	�O[�9ƃ2��!`>����Ú2�2���'{�E��&W� C��s(ha6�_�6���'�vkǀ�e%`u��d��jj���$��e#����:M$-�n�٨��x�N �)�ue¼�S�rٞ��ܷLyٖ߫����ͺ��\sI9��]�b.��|�G	J�ZGs�S�)��H��QK���R�%�Bcn�U}�nW��:���%"�94��Z���v���͆�|!Qt�@����^��WC�/Z�Ϗ�ղQF_lD0v��L�.
(Q��i>����,k��D���u`1�yX���{���kw ��3�T��.�q��>�Ag���Q��خ�����'���R��A|���a�8$��?�֒��.2�Z?��)}�5Ww���������$#����=+�)0�Z�(v�(Cr�p<2,H@���-�����f@W$T��Y,4 Z>8o��yOh����±Ӵ�T%���<�s�9����;�}Ra�|����g�Z���˧��g�i�(��;ſK!r�dV�L�眙����s�S��`���n�ڐǰ���N����*J��%V���l�}V1�]��JB�/�m@˙_�C�2�t�]�t��.�u\y�g�f9����[� ���=����ܹ�����3ɰdܳ��}��g���RJ�YVM�`F
�{Q���De*� א]��50��	���1 \e��b�ua .r�w4n�
,
�'��m���D�ӎu1�*c%��5�[8+���V�J�����j����Sz�Vjr�3@��X_[cб����1�`�c��>��#����5�ɞ%�U���Y( �T&<X�{�j�l�+CUo�8��,�ڷ��f)���A�F{�qP�N�&��P��e �S���U��|�����+%�D5W���hd��kWs�X�ݮ1G�J�XZ��>d�׉�n� Z�p��0���1*c��d����O&]��6�{UX��"��1����*Bۻ��� Ս��\+�وt��D�a��<舀b�~ aÄ���Â���b�1.3Z�g��0_`��+7�z��	�
���Lͨ��pY][	 �	-/?�JL�3��_K���i`�M�l{`�8���0�&-��6(�?��@S֍/�,XɲHq)��Og�Ֆ�����;í p�W����@˒����ɺ
v������k�]S�V]�z! %�a�����=53c�1� �|@r��[��3�L.\�ji�&� K������q��XRM�Ur綹��)�R�`b{���6R����gS�l0((��K�5�͂Er���X<��h{�����4�w��/2�s�Nx�,�ůx��z6�y0è�����ݽs;����5l��eſ�͡޹�~��^2�>��_��y̰Y����3����e�`a;�+�dޑ���bw�qϰ��&S�����ݜn���	��(����GY�T��0�ې���@�i�<I�̯����a�0 �V��I�=Bn]�1��]r�r�z-�[�I�%�U�t�� o&�`w���I9�� ����lRĿ��,�a]&���s�_�k�Gg�T{������+0	��k*)���Ǽ\��S�< ��~#{
2ҤC���=D}Ya�p��6�N�M-any�*���/3W$� �i,�5�T]�t΍�z�w�+xs����"��n�m$��<tȰ��F:���J��Ԣ�����a�:�s�AP����Ѻ�,��3$��lN���c�f���>)69��_x���åۭ�O�k`�ے�#��(t�2K��Oثm���q������f�=�d�:��+(�޹q�&��(��[�InE�u��4cv��ٱT]e���q���(��hw�aqaI��T�����r�PKJ��Dy�*�����>��%�Wd����
�,��H�ڮ����,�G�/�\�,Xq�D�ԐO[[;ъeի�oz�,� \P�n{~.�A�}�gծ�u� ,��U�����?��7����ޥ_�ه�+n'�{"�CJ��O�ݞb׳#��JA�A��$)O�k�r��RvFJ HS!���AV'i0�?��w���@�c��ZF
ۘ�9���8�3XsN�4�@4�h�v}铯t�z'�+i̡aa{��i&���:��ً*�_|-���Р,��D�m�!�h��D �2� P{)Z����￯x�s��2�6�L�����~�ݫnI�k�lt�XH��eM0"�>fCQe��\�͏��E �P^�BO�SQ���_��`k����W�6���@��*��	K�Ok���n�6�K����̼�tl��n�]c�
�@��\G#�{��n�Q�n[�I��O,�>%%ͮ8ڣ3�tЮ��ה�q3�LM��f�-5�a ��jJظ$���p�$�g�e����3����%I��*\v�j9�}7W�T9�Z?�pL���~�A�	d�YY��y_��*��[~Mm�l3��f�4C�U�a��u�&�S� ��T��!��T��ƒ������FK�z��i��gٗt��:�9s�n߹EϞi�����}��(�$ʪ%��Vo�b�R2?���O,0d�� ���f`p��I�pQ�y�9�ԐG�~�~���m�@a��8_)�7 ��F5oK�v�;\���l��\�i�[}D2��U��}������ �=�	 r$4��!W��9u��iv�][]	2y��&s�P���|�5�w��?�	���v���Ɗǹ�g9�5n޺SlE�M�K��uE�'�Lo�d"�q���I�RH�"��ܡ?
����Xk ��=�"i�R��=bf�w��Xs �;�IkA����0��Hg/\���X�����H�[P梐�7�?�*�c9�A�7Q����,�ѵ�^OˁX�}SPX
��H����!�.gU�Edw�"h;'���?�g��Ը��yGn���oTt��B���n������{�))����LCƂ@��j�o���
�� �x�q "���h��_�aKj<4��S�,>|���k� �ТTƁo L, ��?��׮s�>� 	p�<@��[v�Te����p9��T�P�_�`�n��@��F����@�s�O\���	Y#).��̒�����p��oO�@�ʍ�s��o��'S�_��g��5�x�����0��kj
Zc��4�K�g3h!~��ؑܪ��B_x�m�_ ���XI��GY�udЖ���s�XW��$>���I"cIR���Y���l.��<�����J���`r��N��?��a6��R��]J����1���o[�]Cط�,��; ]a�G+"���`۬�'o^�9�e���m�*g�,���%e4%
_�
 �}��&b��̼��`痖ӡ �WWVxs2��-/V^�S,���	\�9�5�}���e����xȵ�Tj#N�U&�d2��a�gb�
t��Z`����
v��lZ�I�R]d׽ȹ�=�X'c��� Q,p`ϐ\Q;4���&@.�e�Gl=�2���I��֜K;����q�"���oO]�9ϯ�[CF����������4�L�S'�f����U}vG�i��^qg*+��4r����#@P�|4�e>c%G���~�t���q<���>龋����jg�����mX�\�G����"�|<%� ����,t9�uk\���F�y��� Jc�e�wU��K9U���@FU��������9�W�ss�����u�������Ǭ��ݷ�g�R��VhQ��TXIaI{���M �b�F���s�p�fM�~�99���K\`�F��v�l���s�6�4i�	����Ÿ�T�[�A�5L���T+�`dڷ�&.B9	������k~-2��۶����t�u�M��@��,��0�y�.]���1f���JU�.9�\!��e�䀴a)����2V�������O(��?�7�
�b�L\MS:���O���T^s0��bW����� ��KA/�	X�  縐�+0�� �v������$��4��X��,�/�	k��@�0ƥ�݈mC�������+��^����@��rPJ�x���O>v�-����*`����GI�r��moo���j e��5�e�ZZ��ѣ�^}=��_���������2�Ǝ�!x��HRбo��}2�v�aV�E � �1�dVQ�ܠ�+H$�C�U�Y�?6��_�2M`�u4ݜT��r���o^�l�okkwY��4ТK3pi�u?�h#�Xͬ$�fQ]���1���XЌ	�/��c<��h���y� ��7*#���X%�ˈ��`���3J��jq�4��=_)&�x���ci�_]�p
ʻZ��*N���56=���.!����"�G��n��&��RJwa6�� hQ���>�kW�q0�7� |�}��,@~,��A�/3�q�n������r����0�b��UAU�r�&�@�ߢ'k�O����ڥ��6�'��oKH947+��ki�`	,����5�v6]A��8|)��R;�dY����{u��)C�?�fŕG�?	a)����Иu�  @߿���6̈́9{��qz��,X>��S:|��򗿤�7�~�b)cd7h��*ۮ�F��F���fX�~?�f���6NhfoDȊ[QܸyRcMB�Y��U;�)��r�`<�l�<_�l�7'�#\Y[��T��-Zb�0��u p៌.#ϫ��8��a����������.��>�! h���;�c9���4ˀoc��)}JM�������.P�l���#�9�Z�Nq5��]) ����1ˇ`.λ΁4i���%�I�`�����@�7ꍃ^�~���
V�ay�y?i��VP�%��!�����&`a {���R�O�m0Í`�(�1�șE������V�j�5��}(��8��{��� KE������Tmgv �����j�{���c�Μf���974B�;B�o��������}��7�h��SZs��*kƔ)�E�=Sye�����P[�����ԟ��oj-pc��(V"����Z�o:���R2l^^�'�������Ź��N"�4��I�7�r��[~p�X��r=�R��%�Y�,�
qPt��y���+}��[j�۔d^�zk[@\����E�a�bO��k"صbf����f��7��ҤJL�iq�r�7^ اa�=|���U��
7����UR&xww�7繰XT56vtnIK��ji$~� ��x��ĥ�1��s|lܜ*�#�����3��t��n^+��\K}�d(�7���K��A2�(C�ٟPȢ�k�Hok3o���������������P���*Z��N���m�V�.IZ�u\Fsg_��JG�yW;�WQ ��5�u&ǅ���&��<;K�/󓁥������7n�O����d�D��e��"��(��"Y:w��;�@=~����Y�� ��?�@�!߮�ܲ����
¬���.P_O����г�T�XL"o�+P�%恁j����:MW����~l �Ϟ=g�QՒ����K+� X~�n�NUǸ���\H)�''3�=�����C�{C�!�n�@�׀�@���>��I ���ɤ�Z�Z��R���XIu��Z��8��ֳ��{�2��"��0���U9�ZA�D�`ɮH�~�2n:�a�)���U�	M������_ЩS����0x~��[9L��6���i��ޒ��+ �ήd�  ��+�{ׂ��|�}%�E�5�������2�����b��B�cS�AV�
�eY�x&��ZV��F����5�w���&��)��>��pF�����sK	����k_s�[�ۉ�"1S�4�&8���m>�����M��k]��4[ﭫ�Υ���DЬ�������s6�N��$7"o��77�b��/�[ȍ6R��!k� ���]�7H:&�D��<g�Ll�y���F� A�Rk�{�8�rlj�gd�n[R8��ѡ�A6�&i��������قv�U���t�t�p_�5��*�!��EHq��ro����X����L��H.�<�T�C�d��d���d���7�v�6�#���r�K�xR�m�8�^Ț6�)�R �t`����r�G�g���c��%���)��Ԉ|���LP�_��ڇ����q;���t�(f�T���v��
�3�_��z�B�\������H.\�>!w.�+��P#@�1��2BLi �B ���
��!of{z�-��x�F�c����#�|En���<Ť���6���� �pgx��13�`M�5��JE[� Y�$�۲%�W*n@����L���|2qS2���Z��=����(��8^#�4�Ӓf��D����@>�	�4��2��8U&��0���5�G���m���OJ�;Q9���hm�8���R��Njc�J�l<���5���ۊ����,7�*s�XQ�<�8q ��%��Z��׀�o��T�'�q�{Ic`����䦙��W�C��x���5��M�V�&���s�l���f��;��,��i��>�B�<Ln��Y�F���n!�&Tu�`V�٘�M��Z��΄�y���K�(��]�67��dsP�7Eɬ��,��F#�@�L᜘� x����Bؑ:�}�9
��	����s��Z�V�s�YVI	�I|%{ L� *�Y@Y�
 �-�+� ���B|UA��ݸ��󾪬����)����Q���
��oLZ���z�3�<�L,���t,� ��7�hcCʮ���4��
�{Gr�b�h*��5=�!�r&���؎�F s0�ej�v�PNxnS��3�F���P�/�� r�"�ldӳ�e�y�ݻ{7�
Ƚ���I�κ�����Y~�RW��<����0���Gk��p �}V*z�f�9+�q��y�B9�י͍A�̬//?e�����.��+�c_ٛ���?�&�3�h! ཱྀ�qN-�u���"\hq�ώ����U9-�]���q�����+{ۊ J+x-�o��V�aC³E�/�
ѡE�w�m�\ Ģ�U.sT�A��|�y,[�誽���W`|[L\�+��c�J���
����[ٚj��/���̾���	�KNf�Ap;oa��Q6�	8�Շ�'&�U�[�>�V�{������_�/�DI��gW�	T_�,-/���PsB�>"x_��@�����2 �K��'�����?��Au��{��}��O�����\x��W6�̈,H ���Z2_VL��̶St��I�t��c$oS���o\����Y��X��%��-y�ipUv�g3!i�����z䙊e������q����%�:'���3[L����n��xX{H�i������/Y�%���A�_����Hvu����5�"�\�tl���E�ae�)�Ԇ�,�N�z�s�R&�`�#�V�3Պ�g������R20��*��Wc�q�N{4� ֠7���\J���-��Ȃ�9�>{\	K���\`*�8���e���ȧ�@�+W����3�<���r�Ok�.�Pay���r7ڋ�?�<�k(���2����Ǐ��Dwn���^	@�R�O�U��� �i���.�sˬ��Ԫ�8(����f�u�>��E�.��ܾ�̭�)|��2��Xj�t^sp�F?��*9�Q���^��f�K?#�&�囥%V���DJ��Yd�lO����.롙�)s_�{C߄� H-)�2�r�����좪���mm�����c�����Ȇ�i-Syqc`�X��e]�*�e*��ڸ�;	K���ȸ��;=/Y���W��rg�Y_�T�-��H�*����]S����-c:01�hꖨmR5�J��4?%_�=�j�[bo�d�Dtzf�.^�D�����λ�ҡ�%� F4���i���/9�d�& �)39Y����uQ�2C�R�k0���+u��9N�P� ����eFYR� �>���; 2��+���p(T#sv�ZWҲ��R��Ƿ&l�Zwj�7�Z�w���gMd�P�JE���S��d��f̖�ƀj�P6�W0������f̤;�K� �tCE36sii�3�:t��qN�<EG�a�����"1
�ک��T�Dos`B�"Bss;�l�^`�jc�8�֤��E��1��mS�ڛR�l,���=����@�(�R}V��r���yb볭E	:�b����Lw��4hX����P�M��/+�֖JuE�R�5���ح  �����Z��	y	3��{�u=���r?|v��u�(����?��:���P��+�s�s�|����q>�����o][Ԛ���6�ԟT\�؟�y�����>|� <�u��P� ���K�|�9\�]-�,ZV�Ԝ��@�넁]�^�s6u��]�k��ʌ����k��15U���F�x� �JY<�x��XtI�4\֛$x���jsGq�bnۜ��+9�������M$w��ϧ��ر�dr�+s^�@?Q� Rc3fp_J�}J b-0l��z&����t���1�}e�>��d��:6ύʿ�j�x�]��s��f�&�W��X��M���+h���7*��9Zo�5�d�#���C�O�ͤ{B��-��`W�ː5`y,�h�sD�1Ґ2���Q�}L�b�3|�X�.������ឦw�{�7Y|�U���0��8;7��v�'������	h�7���nk�x6*:��p���q�>u��|�2kZ6���3�M���Dݤy��r��pǰ1MM�0����D⚓����r�"Y�	�ʆ>is�i�C��%RSv��#�G�;�)��W[:7���`���^��=�m���H�1�4��	ER�t8����x�דT(�T���P*.0�����:}�$9|��>�8�T&��lK�V�Z#�u1W"�t}}��ᨅ��Uh�`��AF���#f�J71K�u��J�X�2���(Р��(>�Ǚ��}�
h�>�H-u���u�6��mpv
 	�q�0�H��RgZ��0R3��ٙY���m����-�-�8�S?>�p䤐��2ψ�yw��^Q,H���!Ap �=�'O��/����,K����[_[r�Ǳ��}T ��9�WWif~>��
�h���,��ʔ=������k�q.��[XZ��nj��
�-��m+k���\䫺Y�3�WX�o��Vt8��c׵ͭmieL�Fd��]Kx���w���ovoE���V�"K�(�H��K|K�ײT���͠��DHY�O+��1�07�u���}-�5^�FY7�kf�DW���� �`��*���w���u�_C�p�26wWhj��UX���B�8r��'�u�����z�*�<������}Z[����x��!�O��8��M 8뗼��?�������Jt]��(�ߴ��x���Mȏ�Vw�Î�-yyglnQ?Sv~Ú���/���ʑ5�LO-�gWT�}�2(H��a����zX�[��@�F)��R�Q{0-@Z����j��lQ�)x����9��4�E����gleS�q�w�KŔ�<<�����	B�*��MM��rM2\k�}ݺD1������U�S�I�)�"��SΫ�%Ӭ�n|T��ϣ��4���sU�-jЪ���U�4"��A�����Nj�5g���y̸>�V��E�U.��$�	�=SƌQ����`��E���#E�=�r2�J�R�����,(�X�}-(!���.�5r�
p<�2�[�[�=��J������k�R�l�e&�U�������{���*}��U:"DKI�}��m6�����+� `&PH"��m��Ø 
0���j���;W�5R���X����Մ���V���%�����"5�k�Y}�c�d�>��!�l��w��	:����^ ��t��E�ułe8U"U ��0G��k�3����?���{b�x���s����}z�]�K���F�Z(�U*#ɽ��J�,qb2.�1&�u�:�Mʪ�l�E,�?���@i���+�>{a����eKgc0O�ˁ�J���̴��!��c��J�� 3� �|�s��"�U5ӽ�=��j�=�=W�c<NdE,���Gy�#C8򙋌h�>��FNPu]hz^��ϕ�'�@��x�x����y�k#�Dw��fcK�X����l���w�=�ד��#���%f6�������v{f�U�{��#JO>�����6�T}Ύ	��f'��Y3C�"Q�P͞�(=(qXoi�Ѧ9X,�lf��=��[��\L.X�C{eSnZ���Ĩ��r�d�m��Ú|�#��K\�v��M y����1��P��4I9E\6=S��ƀ.oP\k�g�LBd�� �	�����n��4��^�ŵ��~��k���|n��qBVl�������1�5��T0���+0?�����c�A�W�J�U ㍳^�v,�Z�G�A�\���<���P���^3ib7�	㚙����dy����;�ӧ�ЩSg؅	@ʺb��m�hp�裏���K4@',F�\�ss����:r�&3_�v���&�\�f2V��ge��p��2����΁�P�v�}��W�&�YP�> `w#���+��������z.�~�^}W�u`8�Ϗs���*�����Wz���R�7�������>C���V�̮8�T�^ΰA�6�F��e�ý��^-v%v�9�ψ�I��$��j�����~�qJss`���YVTfX	���ie�XYU����B���D�l,0�]�Aɽt�29z���!��Ugĸ���l ����Z�R���x���u�'����1�F��ET&���}�i?�~�?��KL�.M ����ꐹ��H��F�W������z�	K�e�����J�w��=+�I�G,���D:��tF����,���fS �Z�YE�t��&Nӑ�X,���ݺ�S�}ş$[��5��3a-�F�����7�|K�����wp������J���9íN���gϜ��!��'˒d9HK���3{���$2o�D(��%Q�`e&���%�v��.ؗ9� ʤs����՚���Vh���)�p��r�����r�E�fZ�q$�?�Ѷ�nW4��u���[Z��!X!�F�灣9���z�1�y㧒V.�[���j�r���.�������cV6��8g� "��σl��\Ul~a�� �x���?|x�����/4{�P�,���
���V����I��,W�s��1v������~�����~����L.�.����5�VO�>d�2�뙳g�H+������å��%�61��*V�|3�#2#r�2s��Ç��҇�|?��<?G<[)֑Ņ�sBY�7-�Tj��n� �p���������o�f��,{T/x0��>^挲�/'���
����t��9���Ϝ�2�p9:w�<�cN�ٝb�&�2 +���A_�_W%V�Z����7�E`3�{I�R��'D^}n�}�ی��U�������kd��zg@7��6�Z��1�\�ddl�A6nv��&W\����Ar��	�t�L��Q��86�!�{N�*�̇��.!�dr�G�5d�||o���¥k��U��,e�2g~�E�_�pd�箎}��D�]��}O�c�Ƶ҃��p`r5����Ş|eB��R��L�e$��1*�����6��Q�.	W^�e�Ur�S�Qa��&`~���u0 aC�咠
� y��q�+L��V��{�(K��������F����҄|-�֖jy<U=iBt룱њ�%>��|#�����j�!����L��b�{9�9�s��%:v�(l^ k2OI|r�a�((&�y�"t��*A1��t�H ![�w
e�ܚ~("�dh�E|�e�Da�76����;�o ��׾�\�̲23=�8@�������:^`DKΌ0�.[7�-��P�sے6lcs]�q���V�Ja-�e@.'�,|�� 	�0��@��[�8p���c�:���F�i�H@�A&���{��[o1��^X�N�>%�k�"�X5,n��@�dPWUΪ��g���W���g/��܂!��Ī2�i���b��\�M�7��cS���!3q��V��Kr���g�)阵��`nX9e�n����w|Zp�itu����7[�@}ؽv�9�k�)%���+'��7[s�:
Z+cF/���H���+����_�A5�S�%H81�҃�r/_��Ż����i%�k
�����*��hL�Iu��?U���D���6J\Zv���(���2�0xۘK}`REIJ����2N���F
 Ӫ�V���.6�8��y1]E#K�R�\�1�E{  ���;,P ,�=ƹ	��L����m���;r�0�E(c�.�Աo�R�N��̈́����Ծ�q����K�#���tt��;M)Uդ3l�s{͔�R���b���ܸQIF���nN�8�@w�\�-.]��9T�RZ����� �&�ȕ�z��@'�ʅ���ޠ���>o�@�)~:T`�V�M<��[��ofq�_�����sS�D.��ŷdUa}��W������oJ�'��� fgZ���2�\��"|_��!��,��-J ���"��0(�G)}�����|=�&ܽw�>��S��/p�ǁJ��96s[�ܣG����,/q�(2q��qΫ
�م�����3���3>���$n�>�_u��(Sȕ�׶�P�0VUe>x�gt�����rA���x��8�5�g���nsRࠤ�g��^�RH�� �|�Q�����so��w��o�O�	JGI��%]���8T-����w�yZ����Bbp,M���}��Gq�SΓ�Pd�]�qqd騢���$�V������ی�����)}��H�V?���}P���t��D�\�ђ�.!VDD�S�N��e�|_�U�O������X��D݂���H�G�TJ쏭mv}�H��)m*�D�/GY��_���Tk�a�1��U�\1v��̌�@��t��O�Z8��p��������������rp"؃Q���ڬ���OH�=����$���aaKp'�և��r�����N���"�fBl��+���f�fyS����--q\���:����I�ݚ�w��e �(Z�	�A6Ox���>W}r�W�F�c������k}�� ��]�#k�<J !�=|��P��}Ѕ�"h�XAEV=so��E��9�I8?*bns	װ�� �A[�`�F��k��=�YDi��5�l��ʧEA�I�X����D~Q�T� `U/��y�GQ�w�-�	c�����[�x�~��;<>��m<�`K��1��(�ۜ�B��G�rК��M�Qg
��fvbk��R���2�}��������+�/��-g��|DQ0ɓ;��`��9��;T_n<�K/���֭[�����mvWh1��s��� x�t�l��b�Ee���"��{&7�Ў��M��מ)��l=z������>�{�""m9�,���j0� 9�e(�wy�j}��f4����M���/&'=Wߓ9���5����:4��`l��}�Ʃo���� z{�5@J��}*�G�k&l�S|����WFb*?W���dw;:u���6���Ņ��DY)�$�]PY���HG��dڹ��K}x%@�(f���Y'�d��Ʃ��*�y_�z^C(+g�����p5���s�xW�KcZ��+�=���ٳ5r(�^H�l�j�0Kݍa2��
hK�)���xM*]�F*�6��}/~�E<ػ��<�nO�v�d�ș�b�?"�w�W�Ktz궛6�0�T-������ ���c�i-�MZ ���-O�D�Y������V�{����Tf�W�r�Ž���P���l���WRL�p��QT�-�E�X�A�j��.W�jGW����5��~���P�er�j����+t��	:w��8y�?.�� ��A��,Ei�������� z�~a3@u���-Z��X�sH�������yv�T.T3�@�jk��>����'".e�v�i�/�~�}��g�� tQ,,&�ޝ<~��z�-���.��8|:�e��m����Go��&����`����Ϟ?��$#h�k���8Uz��s!����'b�䳓�0D�NV��/G?�TJΥ�}�۟l���g^@VfM�+�Wͮ���Sϥ<h��P��x['ֽz_�)Y��{={asK�4&�Q�m�?xM�`_g����a����Q���ǚ�p\F�����>�$)/	
�⿋��
�
�(�՝ꌞ�H��}[0dT�2[�?q���P?at��E�4$�r2�-+ ��7�n{U�3༨�-�Ols�:z��:�,f�<��l�!!Zis���Ps��.H���q��D���F���e?���{���C�����B����Ș5��-��<���~��;���~�QuȃJ�We��9�4A( �k����f32>l!o���
�.��6�q`1�zXڢ��N+�����.T6Z��R	�J�?�d����6����/���B �ω�\T�27�vև��te�0� �8�̫k����Ҿ¤y�n�+� �Z��;��Z]��o��Z��6W4�+֐6�6����~�]��ݹs�Yb0�gN��˗�`F�����{[J�?q��}�]��ű�����4\���Q�%v?zHk�
��FcC'l�I1�1a^���Ү���*�H��×�Ƽ�|�\�����-Tya��z��vO��� ׋+E�S������7W���M&cn��;��q��WH;���ȃ�j���ji$��z$��Ɂ�L@^n����_�A�1��g<w� vv���,�@ �>k�5�8��2�g�~��D�F�_��9g�1eyɟ��u�ߓ�������žk� ξ�>P�l<��S���v�1AD�^�4��=ۡY(͍�Z��.^�ğAX#(��ҥK���������䳇[E��s�f��}�1@���&�u	 ۵�/y�v%(���N�����ד��d�*�v��U�U��E6��D�}3�&,�������z_/�2m�!C9
v%�s=�8/�Sђ ;��&����p>��6�>,���+[�[8�k�p>�|��y#�+�۴�l��`�`����|�on0�0���i�lm��`���O:�޸��8y�+>"@l�<���՝���1`daM*�$(\�q\��fУ�r��w%��d�������3������>��c�����|���ϝc?ܷ޼�i����g�ѷ�~��a�=��,.���<7n��9 �j�`p����++�ic}�vC�����J�=:c[)Y}���~��^��N���e�̾�>�|@.�?]C�q�e}����9U�m����5��4p�:.%��Li��F5	�`����F�����C��FA�A���}#x��0VT9�9��Z֥b�y����9R�@�)O�<��H��8s�0�����o��� 2�lP(��p��������st�Nq܃�`]��r:G'D@~-)�]����V�+���/����T����{fc �Xe�ŝSez��Zk��{�/�|��y�ۿ�[f]��iZ\\��Oh�iɾhP�.b�3�P��X}�^-��t�/�.i�09�*��ɱ� 9���.6���Y��ϳ�L�p����a��Y=4S�+ܟ۟t�k����Y��29��x�N]1K��\��/b�z}Ϡ�MTa�nl�x��C����W��n�\� c*u3������}��QRO�����E:z��?�?~D���iz�q?���Ł=�Ϟ�w࣋�[(Iܖ\�+�(ǻ)��%)���im0�An ��9�@r�6׷i'l[�$�jvE�� �%����w�pv������W�Z�ﭫWi�f�3G�� r���=/\'$��3z��	g[x��9}����
���o��ՕU�x񢤩������Q��"�ug�8F��A�$ł�g�j�ufvRgt~U��\�����ǨPO�S>>p2f���8�n����Z�}�ɐ�i�=>Y_�Yj}����"� v�;IC;���Z����8ׁ���Ǣ�`�b������kܿO��#���� ��QX�:�����Ju��b�!]&�˒�5�#�M|���=���~oMߙҶ�u���x$J�r��&&=?0�f>��`8��^}���:�8��;L��}ya?q�G�XxC���?s���|�x8r��Rv��J���B�D���+)+8ں6��F�w����=~JG���#asǃ���Sku����eԨh�붸+Ҝ��կQR�`�̗�r
{M�'�:a;WӖ�G����O?�?�V�qr�K�l��_d����R}���fw��t�ԯdB�<���먃��
kv�(��a픬"x�.XI�^�N,�޹w��>}ʾ�Yg)���M��T"�Mا�3DI�(�`��C?y�f8��y�6=|���N�YY�OG�c7&��J��=]��x �mz���p�'a��A�/���i)Ȑ��-�"�x ��}���n?�[8��`+,�M�nFq
�̍�mz����|�]��
ݿ��V��hc}���z���3g��ߧ��{�A,d��{�Y�;�*|��=w�Y]���OϦGKK��*��4���h ԃ��t���a��������uSWk! ����`8�X;��ܶ!Z�����ͦQo%L�T�����D�n9�7�JJAW%�F�bn�Y�W"��1�1Fł�kn	��Oz[��ʱ��M���J�*al>�֗��B�1�z����'��(�@� �ǌ�ǟV�����s��(Y���s�l$��j�����ϓB�-��YҪ�+�(p)d�v՞�hS1��y��,8]?s��c�qWU���+��r�������;]'��r�I,M,�M��
e�g����&^G��`~�f_`��t��]d�AB��
�d�I2ϑ0d�ǴSv�"�����%� �%\�+Ȳ��pB\hvV��Z�N���	�I��ie#�_���uX_��%Ap�A$����ì)�����q�`K�҅N#��6&��,���1 �|mD:�?�6�<�lR�bm}�3\&�g�� ��V6������R�eҬ�U)�Q�H��i��$��P��4s��s��$��ɹ;�t�i�O��5���ЍɥM��G�����b��2a�_\8���b�S%�6T��A?6��lk{���x�V:� �=~L��ܡ� �`�w��ζúJG��:�HǏo�1/^a��w���z��Bo^~3����x�z�e����,=�a�l�e���+�� �z(TA��n;��� [f�ɓg����v�ر�0&���E`���A���N��k��b:���� #66w���J7nܢ/��� ��J}{Z҉]�|��엿���D!E����$����8����I��=y����w�5�N�l�W���`�B~ޛ7o��X����d��U&3bӞ`���Q(����Y\.���k���%a]F-�>��2��&��4���
� �5s��4�������i��o@~�F~gn �H��@���,5��+���.�YO�uo�Hcj��0�B�qnq$@��/�X��X��6�XA�uy���Y�4��W�������Ƀt]#_{v��4|Wa�]铋��
���ݲ.�qQ�S�LL1x_�5q鬮�I�o";�_��:�1�{+���g�ל�� @p��M�/8���|�?��*���!�DIr���%1+X�9���w������[q���@�Y����K�=�]��D��(�Y�1����|%we+7��c�8�R�q��x]��EC�ġ`�����-�g)2Zq�qb�N;N��n������w�q��>|����vha~�7�'O����?z�7�cǎ���i3�
�2�&w�3S��1��JZ�,j�,/�Tn?7��M׬���T��(�ollѣ���Ν{�J#ܭ�]�����}Ӝ�3��n+�@�ig@�mm���&ڻ����	L �����z /Q��2��%������[t� ���<����NH5�� `��k8홵�+@R�ma?7�b��΄{�r7�t����]��Y8�2��AZ2.[�.b�bqI�(Q���3�H7655��eFݒ��1�x���{�_f].�����w����:�K�sC�����{�GO��rቯ���N�<��I�>��+��nz��p��5�m�`���e�v@QŤC��fI�L�3�<��,׺�G3ӷ���)��s$�8�Q&I"��7&gs(��M`��FM/k�ZE��h2�uǗD���9���.+����쭂�f�ߕ�+9��╚�~w��q+펓�F��ۧ�� ~x�"�J�Ա�Ǵ_��miX#g���rF5W��}i�-&�hd�ۧ��?0�Ⱦ�*~����9�M�g����p���\P�giiQ2U!G7�D��p��Cf}!���R�
��,ծ�}Z�t��M�dܭ��]��D�[�Z�-M�V(�	���g�30Ӏ$��v�4���R4AMZ8o�kO�4�v��-�8Z}��2�X��o�
��go��3#��l���q��=f|vz[ȕω�᫇���ɐp}~~��=��fh#� }mu�.���oD�f�Q�`��Ea��i	�B.�n�MWA���tY���u8��m��_���sYF?Y�u7;;OsA{�*^�@Rda)��X�"	R�k[|�z}ɍ������U�s�.�~V�ۊmQ���o�$�n����6�
���\��ׯ���mι{ፋa�?�#P0&��h�{)VVi{�"��M�sG�}8��h�_�� 6�97��0����x����p0`��~ ���2^����
�M:y����S���%M�,��b�I'��ો�F��ǟ|B���e���S���k�F���׃� <W�ԝ��ਜ�һl�j��|��m��������ƀ��w�k7��c���3�H��p��Yq&��1U��]0yc�"�Rd���X@*�S/�[,��뀧&=����S#�+1����2��;s�N��q\l��kl���eS�]�:Զ�
�G�.�(1��|��H�'>�=v��{,6�*�IH����ʙe������>0C�5ݦ��ôhH8�x|�JQ��1�x�2[DW~TS��\�|
�r�{��r2�uٵl�[�ߦ�5�T��E/`e:s�,mm���n
V|��gvf��I�h�rg3�1�y�?��;�ly�֥0�t�Q�q�Z�)mF�֕������?c�n���3�����6am�-S�UZb�t()+����B�B��&�1-��|��I�`�o#����U�.'B�I Xw'샰�>f��2��:7�Ug�>k���}:~�$�2b���ag��AhH쾹�ž)�������ɱ��1�.��N�+�{˘�$���5�T������Z=���ތ��c��'=�4�-K絰r� ���nW�mн{����;4q/�jjz��f�9���,g�7��m����=���<�X�X`���
]`���26J�KH��O]��7?�q(���W2)��փ�{�6]�z��x�:y��=w�3�Pv�U����-�E�Q�Z �`W�r�C�s�_���w�������g�!�;�����\ߢC�0�P��L��e�K.����<���1��q��}��0N�5�� ;��愪�x𸷻c��5
`���t�ر�����w�}K_]�2��9����<i�`0��m�/j����Kl��9.e��RYS�r]��.�	<Y��Xi�4@H��'��T��?9�5���'�}V`3�
�zή�S2pg,��k�/�&��7��u~^��x���b�6%@@dդOH���l��������$y�/������c.�4uC�~(�nuoȀ�����]&��oLl�uhe�ϴ��c�h�:>�Y��#gw�x��/r�8����p�Ue�(����L2���uՒg,�x˚�9P�����DJ1(�K�1�w�#�ߒʙd���� U�c����6Hw��w%.��K��)V2�et���-+[��O)�p�Df7.{-QkT7*��	i5$�Z~��a�D`K��6k�0��3ϬA�R�<@�_~I�k�o;В������s"��f�J���B�y9)�]�RwؙL$ǂ���$�n��߻���+A)��V��߳�D����:Gpon�р���1�	�2�qfCʇ�id��d�~�H�cl�����[�;G�L�b��`G�� �jgg��f K3\H�!pk�𜇶\��u;=5��,������R�}C	�����ÚC���7npN�{�n�g�2����FU�J�n��u \��o�|����q������>}��l�?}�4�������3�_�0�,EgZ�A��x��P8�d&9tO�I:U��G�q;|�rh�" mw&��N����g�Avl�uk}m��ߦg�8ġ�ô�xH|��"�աC�,������ ���<g� ?���/>�<<#�{��	�A��}=����~~/ ��e���F�iLGc⒴�3W�<u�Ξ9+}}a�(l�Vfz�sO��\֗K����ct����[(�����Jx�i�*\f�9�m���i�jl�]�J!��G�XJf�&9e ���|2�~������� ��P�c� @⿵ۢ������
v����<�U��s%�Y�6���VU�꾳��M����dv�3�Q�J�bo�*_�B�E���R�~�����}�܋A��}i� ;�|�G1�L�t�R�.��G�U�r�E
n ��a`�%��g<�H+����5E	.T7nޠ'aNY�]�.�֦ͱDp���>�p[:磕_��vK_V'�>&��LLTv#0�����҉S'x�w��q}c����,y�̑��n@�����鳰��7h�����9��W�'��.���ee�)ت ��W׸(L�^�d�Y��_eӑ�ʲ�����쳏�4x���Q��Š���D�c������e)5
�&�{6L��n��9ѓ�l��J��\�eeܫcK���+��p�*��o�K�5�?��Ɋ����P�v%+��G��!6=>k���s�ztm|�0��s{7����#�̶�:!����MO4{Yc�`E�^�J_�5-?}�%v�p4�5n��E�S5�۾r��:�?ۈK�';q�g�U�/�ix��<�Ǐp�|aO;β�:7;� ���oQ��]f�������J�2����������Z�혿�)y��bC@��uF�~�˖����>�;�os.Kl6�'~���HE��� }¹.�?O.��1 *ج�,:$w�:���[oq)� ?�9����������t��M�PA�1��E��n���4�ߎd���a�9?�@��]~�2�q���s�X��mKK�2	�̢�6>Ŗ�ק��],��D_+���7	+�
"���>�-2\���${���E�6k`7]2$�d�f� 9=��E �t#
�(�q���	��)�E��A�x�`7�ca�����l}��f,y�N�T���lb�^�W�r���
o��3�Q�n�~��A�?�?{�zZ��
`^��1%͏ܧw?n��%��*E�u~�u�xҼ
�_�*󎻆��Y�񬷐Aj0d����B�sR����.����,�=\:����p��BLHL�B��D+X�$�%5n
�㘂2����9}"��7+?[���j1���vW�)�C>�v�OVD�~��Wt#O�����e?A�f�;�sP(o�<�=v���5���qkwZz�=	B�Z�fx�}������ՇI�Р� �$׮}��m����`�����-��;���lГ'ˬ���В�łl�n�&d��ˮk��Q�͝L���43��*D���Mڟ�HD�!J]��X��hS�3�K�z�n���87���DV٢��aVb�Qf�]��.Gk�_v��b߾}���VY�30��Rg)!�Qf�d�A��b&���g׬C��7(�A^=
��u�|�(��B�@X�����\2˸�
򰄙�Û�k����	��� �,� �ww��': �)�Dpݹ b������2�Bw�˩�?_� 3�/d����Y�j�;�Տv�`d�� �A9G`ٽ{w��9�fEo r/^�Ȭ.����%���O?���%GJ^a�ʨ`�B+m�aE�Oܹ�V`�z�i�Ν�^�P�twJ�P���ԍ��V�,^C�{�x�$R�\����M�ĬZ�GҾ"ѐ�K�C�kƹ�(E��� K�U����ێ���x��+e{p��b�Wۣ��G��ݰ�w>^B,f2��#�������(F2<�&gi����$l}�����C��C�Pv�>�_��u��p���u|����*�d�$�����]}�y�M�I�:�JArv���\��(�'碻)�	Y@��/\�X���D�r��i��P�0O���~��'a/��2n��<���a-��'�wt�s�(:y,���շ��&Mj�!�D��z3ߤ����8��|t���4U��8%#�{{��ϻ¢h�`Ba� ���bj+��al[�t9�[��3!6�۱����Pp�˗�b��>�;[�j���g��������TЋ�`>���_�)k��M@g&����Z��J#�3%���o��VWD���_0���\g0�~YA`	�8LV`�������D!� 'i9NK��B�D�=b`x��Ml`/�ǵ��f��?��ˍ�`�!�%/��ͣ� z���o\�������,��\$�8iz+��A0�ƺ" V���{��Np�M��.�i�v  � �ag��}(��6[� �a��wp]�[��62��/n��
?Kl@ �ȳ�r�KK���P!L�9r��{�=:{�o\�S]~>O����}��7�[K>|�唍9���e���xh��Z��Q�p'�)?O!��E�3sf�w��n�[�.����A�>S��m�E���Y3������4T��*���h���s�'I�="sA��8�|�6� ��i^���Q�Tf �T�7�����zQbQ\|����c�٥���ۥV�u�u�2�Ϫ���O��k�n����Gq���5�L�b?K%���>�5%����[�4L��9�#�એAN@֠:#�R�d9�Az�
����1��+W�����7��'���d����eZ/ލ�%Y�Ǒ��+i)y�I1ٍA����EYB���M�$����L���)�Q�	��t���}���N��� ��l�7ҋ7��������+18���7hnv�������"z�]�"�]���v�2�>���D�'���j5�ݽ�V?/���#4�e?��I6����S���چ
!5�k�o��@;<@]u�_���������X�YD?@��gO�Н;`sor9I@`���	<_Q�h� �㟨��}�<�ZQ �.P�����������b�-��L
�k�7��4O#:9 ��� Pri{�0 �ۻ��m������ �;�#�X�)���P�{�`��N��K2�����ЈbǏg��7oq���B�,..r?��b�z? �?�����3����[����~J+�Or�&��I3��݁
���:�UL����0���r�P,��,5;�3Ӽ��˲9Z�'s\�	�W�|� ��m����l|:�pNvQl�\K�SRu��1�Ǩ�U>5�C�k����"CΟ:����]��E��%�g%~�B6aΕ^�兙��e6��Mj��漼P�=b?�*�4}c���v��}9l�F.�<�	�Hw.�WO-��z�5��d���
�M���~/��|�!#76����k�z����1PV�����#�萑����SAs�s���è�¾��j�U�MW)m�j1h��*�MQ:YKx�]f3$�-��-�z���8ɹF�B�@�&�%_�d�<96��R�R7���K����X��x�Ͱq��Ç���#v�3��խ�0�B�>�:%/�na�7}3桺h*sD�c��&b\h���kI����DA�l#|�x��qK����P���6�߾ӡk�9�\v���/�p�M({ݩ�Vܥ��u6!cm��'
���,���w^
{#�(��.g��{�KPZ|�����r��(0Z�߅�6�յfe9�yK<�3�A�7���M�;���X	ra�f�u~���Ő�z��`�����w�|��kRX_�JV,:ʦ�.,,2� ��ݿ���Mf����⾹���]�t�_8������ܾ}��\�Bw��7�h7�����m�8&=��u t1�Z�0N�(�̉�2���iW�VQ�eN�\����^r-(��N?�ed��~5�u�$�M���t���"��6��[izJs~`([���A�Y��]�ӤY����M������I=�o�s�1�٣h����|�5����UC�#-ۃ|���x]��Ә��cv]�G�_�IO��{$ �嫧�lia���@�:��(Ȟ�����n/\&��<Ŷ�|�3���yi�o�P�f�b�����v�*7��$�G��+�hn��|s-����/~A���Cz뭷�F��]���F�X��M	��Fa"st���lR���༒\z�yI~Y�-}�j}���L��?6��s#X�<m�w��}:�"]
�wa�p��f��
�4r0�Z~ӗY��Wuʏ��Q�myd����F��*��A4�I͏ٔ�>?�h��ؿ�U���h62a#Ұ{��@@!���aA���ӧ��#�t����3(��^+���C6U!��b�+���:�Ձ�e�NnOуݙ���itS���q1�ed�&)-���R�)�5���+5��.,.�,�u�;{�V½C�&�pm�e�Yd�@)M���s�\vQ��.�6K^�▵��8���=�6�]��Fg��d&��~.�k��$ȦǏ$h�|�� �����t��Y-x�XaY��-�]<�n��2`�A�.=��d��k���dϑM�qm~u^
@�c!�Z�%qE�K�x�<*mh��!b��U��Iy2�[�N��
���MW�SYf2F��\�[i�"�&���z�s��z��@�Yݢ��;�A�H,��Ϫ+ց���R@J�s��;9���k���<�wU?_!�j�B�L���p���t���s���Zf1V�'����}.��Jӽ�嵓s=��d����x�=%���� ;�\��ݨ��Z*D���a�P�׵4��T�.á��i,�^`W~$鶶�/� Dڐ���1����X�Xc����ޠ��_������@�ns./��dK��,�p����k��}p�������>�'Hw�./80-��P&��I�"Rs��l�d����"�F\ �Z�X	����@osd3��D�g����t��9�NwY0�vi$sw���XK�k^��.�P��h�Z�/����FF��(;.
���J����H.��mnK���"������ZM.�����ν��:;?ϑ�(M{��Yz��	WC�������(Q�;\����{�,��g�-�$ԕ߶*��~�Ln�f���92VƮ��$@��A��|��G��ᇿdfTr�v������g(Hǆ�>��(:���>��+Oi3�c(�Rc��/6�[��R@���f�k�U�D�
d�9�7?;�.��޽�)��|9�Dx��%��O��_�7��� ��g�}��p�8��(�Q�XlE� _ir�l�Ԇ@a{�����(��q�̌9T֩`�z��ؼ|�"M���	ﳏ}��v����}�U�]�^됥q����>Fv�xL�Pe�k����yʸ�c��H}�X��\��Ccx��|6AN�� �H���U�"S�}H�� u�Z�L���%w4���}��))����z�݁(m����'�s��K��U�	j��\	���AJ��e>��A��/��T�S�(����O��(��270��<�İ���Vɉ��2V�d,���
����	�J�#�|(�%zl�X��XfW�K}���򳽏r�v�)^���Y��#���6�� �y�]�������~�M��侅��<��(�8��'*v�s �ױ#�8��v�߻�������qm]�g�DE�o7{�4���r\ieu��֟ ���9[[��w����꫘&Zu���*��V�=�@�i޸��7�*4&�-�Ƞ��ۦvP�?͵t��߫����e2o
y]M��d̐�T�FT�Rj֔B��cC����
R[����ۦ{n�ʳ�B
8q�
}�w�_*}�$)幛	�>���:k�6'I�ۮ���������r�p8D��4�~��d��~�Ԃ���VA�2���)�R4�����1
h�8�z�S�,.ٶ(AVfvg�B�[j	ԕ��$�S��|�H˅�a�~Hϖ��Q ���+���#q�����c�vU�$�l��.>Cz/�/���a�/����eK�$g�"	Qy#�5]���@��T�&)��~|H��ģ3m��	�m�gI>O���\��{Vo�{�7h����xK�_Q(�a2f�0SJ�1���~�JGC�R]Y����j�~��5�^�����J����7�h�Y�%�F�e3�����.�/��
p�����y���㱞�
�aH�J՘�xެSdX{���O�%�!��=Ζ�XI�٘I�-\����H"5���ZV\��刟�a6�f�y�z@�;K9&�Հ���G���.w���`W7���<D��S�3�^��&����+���7\��!�����6�+nL�1X`���N�A=�D��կx�u�=��q�s糲��TϤ����̈��A�"������ѹ�y!VDӋ�I�[烶���:����3���p�o^[�}��9\�%��Y~,c��M,-U�$	d{��� �� ,�<d`�O'�[=~H�c �)uCf>�%��FXڙ36�ʗ��>��x�Y��Z���@�����2$��Ԕ0W��X��w�1�����3p�� �up���o���3N�Z�k˙�a�]R� ������YC�1�,�i����V6����nn�Ed�]O�� ������@/ҋ���3�?<O0�_~�}��G��W_K�(DCT����8��FkOwL���q_���&Ro1������
Y��cY}�us�d0;�y�ߕ���9��~n��U�]9W����Z5�g�r�ףʿm�Xź��d����+�p�3���
�_E�x��#�ū��}�}�wzf��{\f��9ؽV��>��~��>��m�t�&
��L់����/d�!ד��Λ���vNWZ_J�B&�����~�+ޭߏ�n!WFnLc�������������@�e�|9�-?�4>�A�0�k����6N0�����1K.��1�YH)�Q�>oI��>����_Bsi�R�4W�)�ä���Ì��󌶚���:��^06��!�D1.4��Œ�&M8��U�g���qo>�����EZp�)��z���Qż����8��+�� �ۜ��Iy�r�����U�B�S�&����s�� �Q��Yy�:�E#����R��5'�~Ie�sV���Θ)X��_�.�µ8Y!�n&�����{�69��\t��2@� 	̔� Q6�s�}ε�G����p��8=�dK"%Y��I �f��]�ֻ��kWU�t���dc:Tص�Z���6Y�
w�5���q���1X咸H����@��i�8����M�dh�gw���� ��(�͡�0"��j�.����(��@�����RE)f���?����G|@�nߦ#(*QKʞE��������@9�8����^���*�%C1�^�(w0Ϛr�J��ô^���:�g��,��,p�7�s�}i��ܵ'�n�o��Uw!~��jv����$@���}���"O�D��b��ۯ�~$�~m�����c2�4���[g0����?�V��X�=�l}i����NdmK�477�zrV,�'���u��1i��@P�s�\�����/��1�6��X37����x�,��z��� ���J���w8 bk{��C}����_�sg����`>��3����?����w�7H�H��$m�� R̬�O��M9�ڋ��M�5��ʊ�ok�a���6	��~��n����&��{x��%�=H�Y�A�j�t��~��Z?��uf��Q﹟Y!�,`	��<�ź���b��L��(����, ���r*�m~�v�r��p	�l�6 .΃O�~�ͯ�|E�~�1�F�K�9���a�J94�%���l��c}��M-��宓�e�h_���p,~kގAeR����Њ�=w�Ӯk@��F�5�8!�#Aa�9�k-� ,.""/����jQ��3๹���&��ؚ����)7�X���$�H�P��D0���]`�_��+W�~Go��}��g��<4ǂ��fw� �Z}vm�Sz��޴�����%�fW55��3��X��N���U�r�s��u��,�Vɻ��lJjJ��1�ٚʽ���:�-�~��BN�������c/,��C#YΈ]MD�6������vL�M����{��~��$�\�;��c�fL�!l͈���/:�p�E��'���=0�l�T�8H�k���|�����
�K4�U��wT|��Z}��B=��K/��E��w��4�<�-�/5<�Қ�U��K�cd1Mn���������:������?�3���S�O3�ER�'�x��͕7�����;�o���L/<��t�ݕ
D���� �Z	������Z��w5��/C�0.#�7������8~��/��X�<=u촶���|�']ރ	�F��+�.���-�q�qwZ'�u/-�e�7�iqy��D�� �kl�b��e�Z�������<�d?S&|U������>�n`�o�o\��L��Q���}��΁#Q�ǖ&Ø�N��AV�K$�<L�F�Ch#9x�S>�z����(����x�"���
�-h�6�o����hg,�w���}��L�۲w�H��Ǵ�r8Y0�)��/Y[�n�О-�~h�B`���s8|gi�Ο��7���i}mꀵ��jV�o�NC׶�d[ k����r�?�@\�+�:s���v�"����V�mh�yz��L#O?AK(�>��X?�s�� ��������?� <�w�;0�iZǳ���)���$����0m 3�:�W2�W��u��P`��ݲ��4zہƖ~Ɓ���>:0�����Z�|�i���6�8��3j�1�y�윚�)t�G�`�3��˪t��Ly߷�TL�d�/��B�	�SM����7;��4��6=)iU������N+U,�XL^�T�1eA�S��)��C�)l)^��y��R	�� a������p+n�
����fLW�l[WS+��Fea(�9P~ȼ�cJ;RGKQAʼ�D��-�2�$�o���]��Ez�O>��yX1խ��Ӆ�.����|�d� k7�ߠ���}�{;�����lKض ���jd��)��.��S-�4�iBt�ưGz��2�ǫU��3��:4�g.^�g.]��g���`AA�^Y�KF�bj+���)�@�t܀Ɲ��� �X�Cq�X�E�i/��L��$Z~��<�����������l�ed�}��>�����5��h���J�v� a���N��I�D�&��v:��}@c��[��=Na�Ȁ��ni���\t@A(��XS�\|��c*\(�ҩ�5J�%��a2�UCf�ޚ�mPI���q�вـ:�	����/��i�~�ӟHj"�jc,m	^F��A�~�*9Ǿ��I���h��Բ`�xy���t�/�޹@Xc�jֱL6�'��������u���N��|���:}��@x��*kx��acC�c3^C�[���î�H4����1��ϝ=� ���Q$b��=Z�w���up��/�`�{�9���E�A����!z�5�[t����{�}.ݎ��E��
A���<:=�K9��ݣ^��&Qf���r$�L���|�y-u'��GG1Н�b�C����		�9P&,�	*�Gg�c��O�����z�g�:��&��Z9L�k9�q��!�D�bL��}2��7�adx���!���~���W�\L$_�)�
��w�L��-��霕�Vmd�7:f�W��2��/Ʉ@i�I��IeA��l�H.�v�#q1c7R])ۆ��\ӵ�N6�%�#+�D�S�@�}��u�������"L,xy,��[�l3�M ���}�bw��Y�JЁ4c�+�K�kA|��&B\`̘M�f
K���`Ѵ:��H�fG�t'Mn�bU5�'O����࿷�s�3`�݈���ݢ�+�L?( be6��?V-�/�:KÂBJ$�>ؕJQ���95M+�V����jn�k�ى��Ʃ��uS�Z�0֡�����+1l��V�y]fa�^�ǀ���A�C�V���'�˴�eA*� ��#"ah����[[ � �9�V3^��x>t�����;����i��D:I�J�����2˲��a�qpi��F�O?M'O5��ٟ�M[8��cu��1:q섀�f<�s�fb��=ϾҠ0[�Z��;�y:� \��>���1n���D*1WHC�]˧� ڊ��x �/������Z�HS�R¦�<L����7qٺf+��z	�2����;O)�ܷƲ6����`���)-�%�u,�X�$�qLZF�})�|�Oo�_y�����z��4�N�icf%��ەDb)		m����;�	��s���y��H�����/w�s}���`;�#/ ȝ�jg8ў=)�h7��@�oA��
R~0������YN��&S���D�pj9�V��^��D(�ܙ L��C��Q���o�>����T.��4&�+)���x0yQ���'N��L�r��j��xDT%�d,�h��p�ë�}�`40c����������y	9V����%Uϝc?4T��INX\��jR������M����~�4�����b���\g�L����C��`(f�����\�i�t���_I�%�2 ��'�B��E���F��N�C���DνK�4<�0?*�\��(���|y1g�8�sȀs�k||aQ8�z$�� �����S���Z�ϻ��B�xT���kip��5��w��3gc����Ǐca�R�n�\ �%��
F��]���ْ,R�RfOjr��<M��X���u���[5�d��{��Ml}�/��H�nv�Ő�}'i����G�NL��z�&�P`�������	�Y�{ �3f���<�����	83�b�g���#�A�5��VUp`�We���XJ��2��c��������n�t��e\�~�,h�v�-������������k�t������N��'�/���	z#�!�{���3q��UH�褖��o���}�
t}ť�9=9��g`�l��f���ηM���h�2�����h��+v^YB�N�Y�7 ����L�8��u�DYR�0���{7�7�c��>q�� C����A�E����ͩ�Z�Df�D�f�·V����'h����+T��晈A%@q	M}��g�fa`�
�v�F�p3��Ϝ�����.�\�lew�Z �@5�mfc̼}}31%���0��)ǫ���M�g�2�4�U%A1WW�����|%�e*�ş�j}�F3������"�죍�̦��������Jrw��fp��dgΜ�}�u����#)�nrH���=ހ��*�����@+�VXp���ʊh�a91��e��V�Zs 4�H�x��-��~�	�, <,�H��,��X��� ��|�Ѥ�we�2�����|���60�~��(���r	%��w?�b�����.ʬ��MA��ܬ���.�U�,)�*���ޯ��$�M�Ic�Z��g��"J�q�$kܽ��u"�Ř�킧���g��iZ]��ʁz�O���i]0������(���{�K f9��|/�e��A�D��mp�7Ф��| �vT���9�G�=ʗ�Fr8+TE���+ ����2��in�q,��r�%����}�&�Mc*�-�.IW;ry��1$��ڒ<m𝄶��?�¨
�&�+ܜ���4�Y�����쭻X��<rCs���"�'&[�6�U!��� �<����qMS/�������l��+J�6���<�_�xK�8g�w���i��&s7l����� 0n1��}��b�~�\��q3�,G�8�`!p	�zvc8~���.�B��.��\�q��A�X5HU�,�@_f"�6p{{���,(�i��
�q'A��������g�Wi���L��S(�w��cF0���f=_�~����͛t�ԍ��i�!<ŕ��8^ag��	��#�ch`b_[ԙRp�6WӔd�m�+i僸� �#4�W�\���~E��p�6��~�l��|�4)�� ܢ��%l�5���q���Fl��5<|���L�d�0�co������o��
Q4Sl��^����JP���L�(���%����sZJ*�=�{0#�_�6���1LGأP�����q�$ݵ1\/�=���ms״{��R,�௭���l��F,����vFF�+�5�b�ͣ�[�A�9�C�	 (��*�T�����!� �� ~3�L��~A��Ґ�^��kwg���K��r�` ��vG��]�_2P��M[r�F�A'��IF
���@3�Ԡ�S77W��ĵ�\?&��i���4��\!,k�k�e`��c��˘I�'�Ĝ�S4�#�
�sp��\��.����R������F& ���`�&���%��g�ժ\_ξ���!k��2��m֦�=����i@8�,l��[�������KB7����ѰR�(Q�5f%g������ ]��Z�Gh-�Gz�zM�c��pw�d_���]���)W����k]�U��kzZ�#�3�#�����V7����qv��)��"@S<�P@���f��N�X@VA�uE5���ݕ@ԁf�@*�!+�~�߸ή
wn�b�{��unQ5�q��	��>�؍_�Kyawe����*��:�%&��Y唔��� o��2ƲX�D��� A1"�����Y�FIC��6�[��aY��.��W������.�`���}�~��d~R��LE�:(�����J`�U��S�1v��Y������ZZf�}�z����dо�P�YH�]z�,�z��j.�.E�U~S-0�C�	�1�w�Jc��,�����^T�O��gk�p!ez���Ep�����Њ��*�� 6=1�:j�Ҡ.����+�x�=�m-��/(�{҄�^���P%��}GL�����#&�V��R��`J~�(�+��%gC�1wf�v�.�#L�}�&]{	��>�D�E��1�����["�=� K~2���T�D]w��m�<�[�,�m�LkM�d������%�7���HO�6k�i��d곷�m�os�u�-J��a�s�'7��EV����w�W�o���hD Vq�}W�KN/h�' ���@�*��!�Ae��H(h�"cԾo���<�!�C �ë��cO`]9z���"羭���=�)M=�<&}k�V_q�/<�1A��sc<�� KG�J�`�r�_/�L�� G��Jw`��j/!b�8��=��B��v��{�M�E�� ��p�,N���y�[�;�ݽs�n\���kL���":���{.:��������7f���~�67ﳀ��wd�`M�W������nh�����#5��4��Q�˟M����H�0�3�1�6��1��>��p-<��t
\?�1Pº��1�t�:y�qº��s�$֥��=߷yR@']�ߊ����W���2�#�+����*��%Е�X�x(��B��X�S��o�f�+D�Be0��D�����������9�ͫ�A�2xM�s@�m9-�p9V\��].�C��R�Cf4�⑵����;Y�T�A�w%���*>������-n��f�\�D)�3-�j��Wk���6�>�a*���I�Q�	h�Wb�:	ډv��h�ʹT�fu�Ӎ!/�\�8����%/(p�~k��)>̹;A䁼a6�� ��冀#����?��nܼլ�%�m� �l�`y+���t3c��#�nt������*s���ٷ�ew�e!���ˠ��''�-�g`w.3ڌo\$q�0�w)�����f�n��B�
��J��r��olK�E��=�f�zh��(n�y�.���I�B@,�� ͌��4���B����,��z�̜5��\��ݮH7i󺎚l;��_���yA�+�%&>[+[�O�,0m��m���ڮG;�34߁y��
\�q����$��9@n�9m��	n*H�u��5�P�L�B1�eZ^9�'Z��;w�� �,�����\�)�^��n~s�����a�A~7X��n3��g{l���ɴh����{��ϵ�[����o<w�> �6��nU�40�:�5l����#is����~����\d7�<��{�\���۶��n&�������ZW#���ඤ�̥�D;�@+��Y3����s]΃���>����>�"�x�d��E�L �v}��5vv�?7����`0���`��>`A3�Tɧ��;�w��k_�`}}�o֒_��V�������ү����G~D�6  ���`���0����w��#����3���T�1��o��C%ls�#��2㑾T��D�o�7�-��J��>���{��	��Z2`x��q }0)�����|�fwQ�r�;�#΂0K��X��U�IP?ՠ�n.�p�[+��6M� (�Sqv����KI��搅��+����}��¡�UY/�-��M�*����@5�e� #��}�����gF(���}���ځZMj*,�F%kF���¦?���]���iq�"[�:�K�%����9�&����}�7�ٛqm�襜xU�k��oеk�����64'�B܎�5�scc��:ł3�h��GZ�δy^�55��i�&�	-�`e����gUC���}�Rl�5bم�4OB�dT�%]<k�~X����	�P���X~�2N{�	�\,߫���A����A�=[��?����8��&����7H=��]��	�_�o���^{$�;�T�i�jP�H�!�k��w��"s'b�X�-!L�_�t�����Iѩ�.~PQ��WJnh�7S׾�*d�K���B$��r.J�~������W��o���x�?S�ali�Z	�ec���M�rCqYqi` @�|�y*� <����[����f��;���7�n���N�:IW�^��?���8Y:}��,ג:�ٞ/dE���ge��0%�!�,?��eV*�Ț"�����o8jJX\\L����aE����Z?�����_l�V�n+�ZmeA|~������ڤޱ�O?ٷT��ѱtw�H�j�&�E�կT�Zi:.��%��}Re�$:��i���,./Ie�e))�B"��(���U��z���?Tp�Ҋ�?������$)9\*L�5}��bS�N�7�I���<hb�f����54;�+d��?���V �]�4ab�J_ȗ��.�1aWh!�M��!�6��&�ݬ��jR4�d&�����ޣ'~�'��W���!��u2H0�h`�.�[�l�)�LkTћ
�x���֯X�hF�����]��s˱��y��y�1	e�B�s���S�Bk��^o����O��߼�����kw��4��b}`� �}'��r�mKr�8A1պT���V�W���|�]�{97W���>wk����Hz���$wF���t�46�q\�v��v�j+�5a�'oE�[��ɼ�I�h��X(T��]8C��d�n �3X_��}��.n�q�l�4	��2L)+����������f��&�6~�D��cJ.#7B��}}�
]��Sz��'9A;R�%����g��q�g����x.$�_Y9L�[��@5,��-I�s���i*�Ab�S���5��}5���d�l��V�l��Bۥ�����K,DR7��IV[;U�� t���y�\k&��.f�`���e#K� �R�٧�1 QP\a��	��^��l����`B_=zD	��VQ�B�ӓ��?X��E{��}+u\&�.3���.`�QQ�&�M����H����)�9�u�l��rLb"��0I嬝��J&�Zy����k\U��ړ'6ֺ�4�W�y�IOP��	8��f���k�a��9q%m�~K*�f�&U������a�A��<�"Y_@�`��J>��l����7�M����yJ�!��Y�E���>�zAyCǶbB1�*Μ���5��~u��-��tҿ6O��y�ȟ�`�n`����(@�5җJ)��
)��j6��R�A|<�d��$ɋ5O$�vG�T�|M���b?A-\�T��r�ҡyL�H:�����=c���G��~nmn�hg��J6��Ds��F���t;��,�Ī�I4#�J�!�j�9l�_�<(¡A�_�܍�A态-�ջBz��g�;�z��'h�㖺4@Q�o��u8��Eu�I��v�q[Pak�$�Y�B"=��^��ʇ��ԋ�//��:����[Mp$���g˯�I��~�ɟ�s��N��=�+���ἰ� �g�.?�~�C�>��AI�R�A���Q�w���-,Ƭ��W3 +�[iW��)���Hh�k2��>�i%Xb�[���e���##ָϮ���v�5pl*x�E���i��Ǭi�A���Bk��oZ�b<�a�Yw���|�	?e� -@ҿ����+qG3��.�u&���$��݂���������u'~��4v`�փ&��*Ru�*SBH�n�4d/K#ש���d�I�u��?�^����)�.�ǜ�"��z�h	�f(�#��I���T{��+�)�Xym���r|�����m>/0
�M�Fv�I�j��(�$ic#\�ԩaFR2�U7��c3?.��7��ÚP�Sւ2�@�v��Jz��O���g�9�.BV.XH���KX_k��R���� ڱ	D����W~�ؘ� �W�����)2:��=�}1�)49�,����i��-J��Z��3�)6�����#��]��L�v�$�v-�B�&~�bJ� 1�TL�
&,&=X�n�r��v}�y��~#��0��L3ј�������ܦ9�ɓk�1M1;���I>Sf�F��'I%�{[�1�}���~|t��L&-�D`5H���+)b �Z5." Y����x�{�f��my㾦vrpZe��+�g�B���3�g��4�) �l����p�N���i�B��ֽ��"��7�>r�L���:�S*�����',��6�-|�'g�8ۘOk�7�M�PF�p;��fc�mPh�_^��'�[��~U��H)#��o.���Pl��r�5�ʦ)]�(\�:�_��t���L7�����3ݻ_s��P�z G�Sl���s�*��ƞв����H��R� P�2�]�?�.PU]Q*�lE�ƚ�֨{Qn$����g��dZ�II���"�A��+�c�;4n�^��l�y���V^X�쟘�5������`������3��_Ө�?N�<l���wΙpU�9-4�Yi+ӻm�����;M�?���R�����#믲%�X����WG���q��<�}\����M/`{I2qX�I�Rɺ�3B��Sb�u�f����8a��7e�TZ��+m����X��Hcp1%��&k��M���XJ1��1���?v���8.����#��3�%���l;�6�C##�>���{kw�0�WB��T�T0��Y����L3(0P_P���l�>�Շ��{3&|��<���Q5m�=ds����Br+��\;Z.�v�0�.���r&���u̍Q�{v��5��A�*�=�fLc�1�t4��H:Pf� KI�j1���>Jk�`G���?�抵���i%�웏�D�7����H��[PƂ4yxn��]ݬ�3�Y��`.�0���Z&R���[h��L�z_>��`�瞼R�h�;���f��k��ݢ* o�
]g�1�9^�+�j)iP�8�䓆�o�5s��*.Y�C��7�jrԻ�ܦ���P�?�e̽Rp&�e��B���4�\��6YX��[��~�ј�>�/&	��ϥ~#^�$�|�n@��m>�S|J{�>�1y�{�b�.���ե�؁S*��\�T�~�a3�->�u�(	h�qb͐��c�IY���hĶ�̟���&��.34��=Қ��q�Aj��B�C%} ��`�VF��6aq���K/�D?������;�2|�ťeH��\�&�[�V1���/~�P-�O���0���9O�3NZ��Y���[Z��|a��|.�ޣ�x�����\I�m�8hI�D�2�y��y�L����av4[ޛ��Q5�"�"��r��� �<���m`hV�O��{t=	X�vf'�o�J}�+��+<����x�Б܆F9e�Y7�A�ZT�
�V�.�:��G8X��������3rJ�(uA#85-FKKE4!��n������� �����eN�;W������>WI�,8*�*2�ԙA����W3`Q%.?��JJ�-fv�Z��gϱu��MOМw��=�H���9&�ͨCۇ45-T�9
d�P����G�,=x�Aǎ��R�(J"���*����oܸ���|���n��"�8�B��݌��u�o��j+Z޾�m��` ���ڄ��o�d��O|5m�~�����Nм�\�b%�I������n\[��⥩d�h�=m���Y�>��=A��c9M�Ɛ�1'1�p��#���Oӛo�I��J�.^�#G�rZ2��M���{��)���j �����[o��I��+����Zf�����m��mL�gUҶٿf���0=�
q�������)�b2�M:��[��E����ң����a�Gv���i%��P��晵�(�0���Bb����QYY?!�@�]s��$����o��ʚ��)�N��J9(`����lsp�n.�/�\�I�����D�Ƣ7k��ҞR#C]!��9��F���;Dś	��cmeLľ��ĳE=Əa����0�7�;�������|e�����Ϣ�pڛ@���4�9��������ftQ,Z��ǎ����rU���O艦Y��2_|�}����vk�P��Q�M<K�.Y�T2G�*#�XG'P�\�9�{��JO,/q�h��}7�d�Yb%у���,jҷ	k$ۍ;�m��vo?��fn��̛�
@S�(�gn��@������P�{�%��?_�6ܙ���V����,��z*J��bUAG��%� �>so��O�^��f�m��yr�)�y/��b��;�X�/�~B�1��pᩧ��f�B���/��WK���`�cq����vMK�� (h�N�8I��G�� 2�I��Vl�7�	�7��*�;=�(�WΕ�؍a��*~�&xҘ���
�S�e�����k�9~?Ji���od�4v:W�?Ps���F��\�kP�E-�vQF�͎���`|U- @ܤT��,�n���\J���A���:j���6qOZ�us �մ�����9T5�Hö���|̣8+Ü�;P����������45���ܜ�T�&s����#���\��ZT���Ḯ��`Ye����=O�s~_ί�l�E��1%�9��sJ����O͘{�`�+*`!P-��I�m��9�+OE-,����t��������D��?�@��CJ��x��� �?�ןЍ7��y��:dw����X����ÂhD�UCǚ�Ԗ�0�f�e��ɓ�ēO�/� Wb���pޣ����b{�t�ޝ�1鳥��s�u���'��ElI������řbqNўHr�4����E%XS����wc��t#�5���r
�	���P���w�_���c�����
`*
��2�4c��.�5�A��V�yŲ#��\A�KS'Sb��`׃���9�^绂
� 1��˿�+��?����>�AC��7`�|*��q_lm����VkV�
�`kk����9�R�*3�h�J~3�g��Z�V�j)�|ޘ�mN�Z�r����+��t<V��h��RR�QM������ό�f` C��#��������4Z �(+
'�y���	�̀HI�\��h>��4��D
K5��B��ƖJ�g�N��\ �V�������@���R�)�BM�˴]m�n�e��}d�y�G���tD�%z���57���5H�Ae��ج	Q�����D��֜Jlcs�N�'E0���`�Ҁ����%~?�B���A�r�YP���%PԬ�A�4WkKր�:����d����u��f� �f��^����o���B}>ϙ!HiߘS�������Z�`h%R������%�BAA��(�{z�4���r9KE[\hi����n���k�͵����r�rGȅ,����ex���bB9��hko6 ���>�`h�߇+����;�:�������6(�'Q?ߖ5/ds5~��M�@#���!W$��E�,w,�W^{6I82ǚ�V��cmu���E���9=B�kgɳ�.�����i�(��=��Pq�Lf0ۧ�r��U�����C���M7��\��|�s@o�c��[:����w/+	��z,|�C�����J�:��?�d��+�U��L����qK�Y=��x�h�����0�(��y�+�޹}�+M~��t��uZ�āq�����=`�`R��R�F�B7��@l�fӛi�.\x��y�.��M|��MZ_[��� ���3�y��K��l@�
M@���Ïd�ܺВ����&)�(d�-����{������Z�.k��IcO�3]�4ܦ�3��	����I����6q&f~B��)b���ߐ�ZT� ��A}��>λ�- ��x��:QǬ	"m��5ir�%�	Q)���JG�%J�ùm�T�����;&�B���NA�)�=~ L�Z�V�9=H�\�|�hs'�SCԁ{�N����`�>g�1	��i|n=�}[w��-���𴑺[���L�@A���H�W�K?�����1�[���B��{~���%S�<l��������ֵ�%�e��!ADj��9؛NS�W/áw� �Yc�"��
x�y���� ��抩u������ˊ�cڶ�q`Y#S��տ|�R�k�w����h���]�~*ω����}�������>����o��vkl^v�ʝI�ƃ�X=rOoB�m���ٺ��3ݣo9�T�nEk�c���p� [A��7�RL�����^��{�Ξ=���T:���RQ���Ziι��F����7�������4�c��sM�I���=�]Tb��t?
df	I��O>�~�ml<`�v��<�_����v1�J��V��*h-Q\Q���+�����Q�Z�}{p�F+�  �2?]���3����ݻo�'��
�� ���7��]H�l�`���a�u�Y{Ԝ� ��$��b��t3���-wH��4�Wq[XH��r�
���M{�ڴ�Qb�|?D�o�ֺ�����B�)VA
�
.�/k��ܻ'	$�K����>?���ì�X�OD$3��q��ch���߾�fn-҃vJ��0�%`=���d���3=.�c��i~��[�jd��@`J,�8��T|r��O�.���;}��Q���|����7I��v�P��b����@�@R9��	h���T�)��tAS��sB�?}K�y}&��c��{�P�(]���*F���Ce�L��G�BƤ��N��o���fw�9Z�����c����������H?�����.-/J�� y�"p�x����
+�.]���]����6�[�E��k��	�M/*�Df�ґU�R2)\�r�~����?��?4�G��5���MK��8kJ�5I�@��F��H�F�����E�w<�����n(>\�{.�<�\���`&��=g�h��=2��D�bÜ�x C�ʹ}9U�8���Y>��W�z'l�G�l�얜3���f����A�XaS/��n��`6��wG��3�]��d)W�����5�iq$H`�M�[��i�9�O���$�-�k��Wȳ5��6�l֜�u��Ƿ܌I&�Է�ی�4��f;Cf�O�/�n��������Dh���`��[M4X����&k��9�4�YP�g���?�џ���/�������������x�д���vM ��Si�8�p���f�:cM�7���s��cA��[��-�S�Y�@�K͈�ߖ��?��=6��*�����4��4@�ya��1�F��)�X���6� �47�*���6�_���7SZ��߭��{���q:q�mkk�hcc��ܹ��Y�k���c��|s,1;{��}�Y:�<�5<�&���S�=��������+ݖ���$� H�,	#�?���c�X�T*��ppLʻ����uo���?	��c�B!I�S�q�MF!�g��x\���GR�dMH^Kb�n��o�st���-i�*�"?=;��h�5�T�˴��IƂ��"QMo`*Ø�g�Y`Z2m9&%�Az�T}Ak����-+�m�/b��,�q��M�'%`fK���XA�?08mO��+0 ��8kU�3Th����Ԣi�$@�����I�P#m������~!+ʣ����q�{��X�1�)+����{O{�B˲��D�'��X,�Y�3�����Ǵ/����cP+�êDe��z�n
��2�
IAbA�$��R�Tr2�� ��>�k�.]�ľ�, r��]�gΜf��\����>�
�Vi�݆�g�jp-�m��"~��!�83}�V��y��J8��N��
K�M���[�����Fi�t��6�ir-��
�{K��R��L{,+T��D��9I8��-��GJ��L�o�<���(2+��s�����/E?������������������]��P�dD�/���l����4�v�t�;��M�&���w��RM/�h���|#��	ZVH�L�b��g���.����[�u�� Zh��ӧN7�5��3~C���iާ +7`���*��A	�H�O|�e�o~<D�z�ե�����fd��.Kc3ݧ�4�$i��+3�HE���v�}�*��ˊ��m�$D����[}���� �c�̒�R%b�d�����vׄu���A�]�$�
`�(E���7'����3�^���R���A3!Y0��1���]���9UJ)�* �F����^��o1��Ɨ�Dۥ�3�]��͆�<��=a-���Z���'�v-)�a�Ǚ��v�{��[UO 7�����uL����K3��YKz}Γ˕8%3�	�L��� ��/0����F�����>̱(&����t��5����`A�h��l:r[#�R�!���� � �f���UN[g|��y:3C^��<�o�z-���I�R��
&5/�$�0?Ԯ5�ݗ8���k�QIQ�= ؀S��W�� ��_�t�	���+{��@])��8jR�K�����R��������@<�ٍ�s�2)�n��{��ɿ���~�-�h�n�sRi�[O>��^X:k�&��!�l��?�{{,b���8�gW5>���FI�C]H�� `�=r��s���26�!f��M�?ض�3�!/���OjL�DмGMf4���|�2;M_x�������醘�� �_~y��}���OJ����].�
�.�P�|�̽N1K�0�M2(��2�ٳ�/�jpmh��i����%1pщja��̪{7�"m%���#/!�d�"�ޡ��5f�ѾGGk�g�_e߲���PЯ�`��
�����6#����$�}�$tEݴeBq�=����:A&���(9��ʩ���"�`������[D0�/��U���`���~��w��HS�-,"����ᦹR��ϸ��.>d�@3/��ǽ���߃]3za}r`LIm}ɹ�@�t6?�8x!~?�3�i��r����ń�i�*Q�hԴ|9a��5�;t�F�HK��$��2ׂ�nh���ݽ}�S;r��C���cj����t�"�ښ8��5P�P��9��z��5�vc��r���$x�.x���JRm
E?@��-��1�ެ�����KոI��z����Nu�/���:C:��0E��,��~>��Uw�g�L���Tq��a��Y&�W
��v_ɀ��4c����Z�U�L��<c��R��Y�xt�I�8�mϋ�<��p�f�{rݦ$.���i��@!�`�S�����կ~M��}��U^�m�p��,�{�׸h�G�@���,��c�fu�yȥ��tc ��s5c:��#'e��׺���kJ��t��GO��[�C>k/��b#9���B�\<��ct��ma��.���N?�	 �.�{���i��m�-���;1����gm����^sО��;�����4{�Rk�%���T|���.4�Հ�qN��I����o}�γ�;G�KYMhuk������(*O)hd���#G���?��k��z���I�3a=�{'� X���r�*n$�V.(��M�m�[������4i�zu�;/����אt5\2���c�zSU���/t����~�@�>��u���//��S�EԢ y��r�h٢��o�@��V4_+�p�m[�Y�c�ji>5ݢ���
g�{�����7n�d�������p��z�@BC���h����9�x���]�,����M�)���в�x�A�_��TW��@%����!�ˋ�pB1�Q��ͱ\B��ךNC
E�>��dH��q��@7�*s`{Ѐ�ioc��}�̡'�ÎV�}�UyeO{ 
z�:�+
e)���Є���RQ��֦�ա��G`���u��+:�=�y�ٲ���
��x>{�溏O��.�	�W�S�4�DbiUҪ�j���mb��ػ�-v��oՂ� �w��].t)@מ�Rs$��׾�[@��&Īa�z�m.&����^�ot�4*ű��2`5��	xEA��`O2��@�]����86�*����2�y(z�x�#��SA.Gjk�z�AHy�JQ	��q"|ޅa�}��h���9m�N����P��`?`f��
.��^ҷլ_�W)�Q�2�Qsp0��*VP�t����3�Qư��%��q�8��2-M����^L����\�˓T�$��M��.������Ӟ�ڒ৿�8���Ϝ�n�t����V!�`=#P�'�7�'���c����9���-�ݰ�7�5�:3�^m��P�\�p�d���Ǹ-E��̶��&�@T�n����q5p���Mh�_\����tKɰ�S�s�l6~�jEǩ5�۔����sN���~�,��o�~��RA�l�¯%�Dp�9����@�Z�yH}
>��y��W�g�y�]?�c7�W�u�}��|���w�f������p�yvo]zL歓�TZ��
������L�x8�����յ&!����g�l�g��Ѷ���j&��~���O��+W9ڽ����������n�����]���_{-���86��_Kc���|t���z�d9��R���+�:���g�n�Iu���ڈ.���ـ�a�A�B�Y��H�9͎4�e���4DS��n�x��vMs�Z��-=S�1����z�5��e9�����GHph@D�Z�".��-��s2σX�}coϠ�7B�D��шs�63���Ѓ�8$�@���є�Fh5�S���y�'d�V)��V�f���ed������gj}��?G����M��S�Tz��_oyI�����x\)��fw!0���=z��?� �E�)�_��քa�@-��jr%��g&���u�bc�`�pۿ^pFK�I��-5��}}�kճMf{�gt�A��M������]U8 JM�'s�(9t�-8�1+��|4����|/(f�O��Ѻ��|nr�Ht۔�0ab=��+VI�A�6�g�Bi�4Z��f�u�>K��ڮݻG�O��?��?f_��ׯs�	��v�}����IX��6���'U����6Ĳ� �gw?-ڱ�#v]Pj /@��`�������5��|��{��=r�KH~������o~��/X1��͛L(a��v�J�v��
I�R��*�a�_�u�8R��������fl=�4,�IZ���[��/S��(�V�UK:/�Z�nH��5�7��+�!�On��\Y��c�5������6p�^�$+�B�hZ<ɎR;�۷�[��I
��]�"��-���k�<����b�9��w�4+��F#	ޓ >��Q[�����js5�~�NS�y.:>{����]�kv�3j'�9w4Ebmy�5�A|���e�ѵ�1�>p��N����̧P��M��q'���f@9�z�Ӆ����u,M��4�h@3A㷴�� �0� ���c��t����~ڬ@���,�@���y�<����Z��0�5!<T~M���V�SE>�,2�Hj���D�,����Wcz�����K��Oq!�W_}�i���D��,�F��[o�M������F�U��Z�ٍG;�f����@	.���_2��F���W��̞|�EVۃH�iqi�UR��c�tE>B��K�v9���r���⫈�6*��r�a��R_�L0�"�@�b�H�f≙X��Z@�;<��z���p�MKZ j��7-�U]�O��)T���Yʛ�G�p&����]���n���1��{��ݿ8�R3"�nc.<�Ք���J��W��`� ���cc�1qܩ�6{6g��֓�I���V}O�+���c۝���Z����Ie���W�a��Z�S��V�`�~� �9т�U�:pL`�%̖Z��4J�}��E�ʅV���iX�:n_W�Y�,��Q�9J����ś��z����˥_s�eok�,��$�lխ�T��Z�����\��T`"rn�zl^���_B�c�?}V����`��-7퓝�]���(�'�"?�q����aBOTx��JW��F]'m"���I��<hfIH�HA�)y���r�@Ϻ������v;,`�{5�i�I��z����R��k�_A�
��m�`�Xl�n}��/��������w�jw���3-��WD�׊5��XZ<˰�}�i����3�.*��q���e����w|V��}��cdfm����0@�Q�,<b���������g������!���
JkF���U�����g?�)���_����l9)a6B1f!�Yġ4���hv�Ҋh���_��6�����}��}�V����䍙!�9���Q���(G���> �R�J��vΘ���v�$)��N!M��K�ɧ�䜉7n��A:�H#��j!�,PiaJ�7eAX����ж��[bg��;~��!H
r]�wL�i��i�a�GBZ�<�.�c�Zf����fΕ���.���b�Q���V��l�TN�@�}P`L	����K6�O�b�G��8Q�n������`�h�!c�Xk��3_�]2>��:O����\��5�}7,�%5g 5-hP��eɰ���z�}���J�)�9��L��l��������lB��cJ�Z�-V�ET'p�ϔx�#*'D�7ɭ*~�\�ʽ�����h��T��Z����{R*RB�O.�k���lك�K�g��>�^�
mjou�B���'L��+'�=j��`�ʰ�~������g�ｒr][ys"J����+g��� ��J��P����=@Hh�1浥,(�_�^[[�*�;�X'U�͞b��|�B�"ꋙI�:�KFgc�F�/���.tA����tҺ�}a��X���tְ�n�H�S1G?��e����2ƭֵ�S������P08�V���/��)4^��J�O�m��^-�1I�@�SR)poa�?S�p�u��z�w���B���w���4<�c�њ��9i��=V����[��{����_���"Aj)�6	-�~Ӭ�>�n�7���6u=90f��#b�bگ~�k_����d_ξ��a!)�2:<�R�������Ո�3��@ ❻w�=����_�5����;kx� <�ӠՅfhcc��K����̄�:U���j�R� �W8���O���!�fY���V$B�Eq�6�A���IO:�fs���BJ�R�쏔��5�ζ�݈���i&:!5��qR�`�X�[�F�(�>a�{�q��	C�Ba/c"���=;TK3]gQ1m�6��myX���>���������OUv��4MJ���Bp�b3�
Y�$�bA��o�q�`��b`�\�&��d�h�*i������`,c���{*�� ��F��3�:kUW0^h���EO���x�I��t��i��)���6H�^m��Gz3 ��~h�0���okY	��<ڄy���?g�[ͬ��o{���3��p(Y	�+4m���z͠�e�R`;u`�d>�������̶���r�q��������/>�[��i����J��Q�}�+Ժ}���wS�������)'a��ݤx�;w)�Z�O3��/,,���E0�MQ��oo�M�f��/���KgϞ��^|�^y�N��.�KL��;���7oޢ+�������|�z������W���W���!Z��9��p��]�eR��ˠ]_hJ�V����6�dX$����x~���x��l�T��MX���^Q�f C�+�L�A+Ob��=B]�K���i�Da8�g��I d0ጴ�	`�s�~�;��ٴ �A%A�6�iZ_4 ��H7��jG>�AΥ�G��z�7u.�Q��Y�^49���뷿��4j�"�{G���1Y��D�@�]��AkN�:�i- ����e�3Pܹ}[��7������w��~o-	�I���(&�ޜ��d\��������u�d�v�cf���?9�ꉢc�ȳ���/������W��Ho��&W���y[��</����/Ԕ�C@FL��NO^���(i�uQ����Y쓸��A�B(c�����Gϵ)���*�j�����{hf��+�:6��2�k�]�6U��ZU<���G�}4ݺH#�om��y�O��)c@�S��'ւ�}Cߡ�D�?��?��}�{�=[�-��	<�n�����@�/��e`����pZ]������<)&�Ӎ!m7x�0���.v�_��>�<u���������q{�G�qT�x�� x�TC�����oci���� �^v�䷷�9���������{�!(_0���Ϛ~lѽ�uֺ�҆�a|������wU��H�3fߝ�x�4������ �=���7�m:��B
Zk K�bj��(c<lsTa������-RZGx��C�~�%���L�򊱢��y���jMИ��GJ=/i�P����e�>�{�f~�h��&�Zy��y��Z/�_�m���ME5�Q�ʺ%2ב��M֦������B�{״��I�y��]�4�m��n���8��=���ɓ��#<��^�B�x���F�~���b�`:�<�  KӸ����W�˗��寸�@0��X]z�@�*�[;�"��f;��'3}�o!��ʹ$��?m��v_���s�[˘5�0#J�b<������}�,Y����ϛg<e�i��5���H�C� ����L���[O�В�>]�����%`�X�_�˯��3��Х�������UNd�9�530m�e7������j�E/,�{���R9�m7['m�������旜���T������ܹ�S�h��1���@0$�t7����>����&f�Av���'�L���s>t0����Y�F!D�Y&kI{��	�_�px~����_3т�^����n�0[Y]�����߼r�������5�\� & �H�������}3�|�1���7�xSo���5Pkձ�)Hs.��L����y�2��Q��M��9�KH�J���52#���r� r�f��
���6��L9G�8�1<|��O,Uif{x|�e�th��5W��"�h���
k̍�Ǧopc`F �*d}=֨\��T���G�2S�Z�3�1_�o�?�+�o��q��z������^堨#���˄d\j��&2b���]Xآ`����;� ���sG�;����H����_q��7��dZ���&��h�hx��2YPث�x=�$j�3���Ƅ�b�	I{�~JfQ���=k�}c���E����!�eēl���`��gw�;�6������b4\�SQ��I������(��H���X3^+9������se��UJ����W�|�ge>;2�a���������\A�>�����\��}\���-�k��ƩZ�z��\���Uϴ�r�/8u�Ds�b��{��onq\�ixg�{��:�5Y����4Qd�T�1��=�E��z��� Q��C.,.ѹ�g��_��_�+Ѕ� 4�OV/`320P��q�M�O_�Լ.�����1��ظ���j���(U>�7�:å���5�)ܽ��H;�]9�L@�Q��G�\~'6.��%�&J��Z��'�� 2���5�A}�௒���]��uu'�ӵ�?3���F "���Dp�I��Hgom�nL�}�h�k��)���f1����'�����,z�(��e;�	`�R|�Y͛�y�G�q��Й~�7��9|�5���<���ޫ�s�%N��|��K���ޭ���F���Wm�Sdm+�!��۷n1��pW��gL2�A�&�6�v��d����J
�`~Μ9���-���Mkk�c˚{"�A���Ʃ��@�U���Ut_����(d���I<qZY?���E�n=Zm��@�@�O�<Հ��n�˃o�PC9�ht�cpe�*�\'�i��[6i���<&�O�F��_�3��{w����u��׬��ꫯ���ZA�Js�J
1��V�S����!u��b|:c�]X��~T��v��i��-k�c�#��%�a�~�Nk�J��XW�>�ڇ��J��lI�؈�|݌5�4�����:��:mS��R���J-W��m�:�|�,=�	�d��$M���VH�mȲ�HTS�6S��#��i����3@>C��u��]o�쒙ƹ���^Z�<��vtʥ�:攐y��/.��^�%���0��5[��Ђ���>f�9,��]j�a\�sU-t�ͅ-�:����3�G�b|cS��\�[�F�u��,8�L�/]����n	(���q�������t�"�������y��^{�u������VU& �M���Ri��#1Ȧi��"*1��y��Ƣ�q4���!��<П�����x�kt�	J�i�؜�����Y0� ����%�2���JֵcR��h�$8iaIrO�wgk�vw�h��Jè�2��q�:}�������-yt�9a��A`�Ff�0�^�hB�8n	��&���ҥ!R��fF_s��a+S�Ύ%�l-xV�h�BP4P�K����Tw��*�8���zK	�I�����Ԃ���P@���<��"����Қi`�oҼ�5����%�"��� OA��'D>��g��Ґ��;�(�"����$h3�RF6״�1�K��63����ޓK\^�/����=�����J
J5c�����{Wsc��z�B�9kuҘj��c�̧�_���"���O�/�H���}�@_n߹�3��q,t3cЁq`O��ޓ���{kt�[4j���[��qYc�X#<��U<���{x|����Tn}s��R���:_�t31�yr��^��^;g�i��d��FL������Ԥ���o�̦�N2�Z�h����|�I߂5|�a%D�k�h�}�@�)�����u�az��Z�҅C4�&��&����|�����z��c�P��h���iCD�������9�-�����-{����vµ�N�Q��ze4�ֲW����2� ��.� ��#����5ퟬ �-�T��)r��
Mq埳�C�!	��J��z#�v�M�g��2�*�����~��J}�a�s7]��?��g�<�г����u��W|���<w�*��X�s�И��O�V��]���^�L���8��G?������?z�M2�i�,���u�	�� �l����������E�ح[�R�(�f7��eP��L[�Cz⩧�����}���o���y�>�2w	�LHo�{V
t�>'"`�\�N�t]��Y�m�Z:��  �PIDAT��˴���ni����+o&�KZÚ��B�I��
B�g�>��G�L�[���:F��\��%'�Tz��\�xv���n�΃I��'��umÇ�H����;I0����M�Jv��!���A����Za��Ul8i��.˾�r/������񆐋R��Z���0=�����tm�)/�[
F,0��F����D�xإ��������PV��^9LG��?x���?�#��uom�n~��!@i!6{�PCoV�����{��^4�cHP���}�&]��5�l�>��>��S�կC�������t��'/a�Jo~ހ޷�z�~�����5�]��6��^�=�a��o}~�yo����'+{cAg�f���2�����V��]Ο���*����hռ�H�
��-5��`�O�wnD1`U#��0-m����[�ڼe�:���=�6�K��< �<��Nꓟs�'ň
�b��uʢ����3!��Y�;�~A#�|��@$+��RmӬ^9c���p�!,�}�o�O�����oV���C:y��Ez1��Q�2Ll߻��%S|ve���4m������fH�f�Ti�y�D^]=L/��2k#$}�.�VQW	���c@0�/_f_]h-�;J�N�a��s�����0�o8/.��c��|�\�Q�5vR�	�C+������
� @����k WG�g�"�u��צ�UEB��>��L����#�����|0ͬ`�\C�Z�	�3U��2�wX��6���`��@��8���9�J� |Tn�{�0I�4�\���P���4�����̖�:k����		P�G|y����"liqiB_f'��W&l�A�0�5��-P\^��G�6{�4WVҾLh��: ����`7�EC�b Y�_k���ӧ�䉓�u��%�GV5-T�<����Ȼl�ٿw�ܣO>�������x�~�fF��6�.ȟ�+�\`����SO_����*���7�bC�N�<A6w���~��t��S��?r�:v�B�~� �a3ޣ��q]Ͷ�b�Ih�6�{��9� N᫯.��/?��}�{.���3��`ܖ����/��#�Ĺ'�FH��ttl�G��Uq>�W��&҃`�<�����F���$t�n
�W3���u��{?÷!��D���;w6)���[��O���.s�i��M��(#����R��ѐf�[Ҁ���05,5����Lg�ɓ��|���qRp�V��@��?%��T)2�tZSz�>�k��%s�*��~��K�R�D2�:�k��ϽÞ4M�sn��`Y�Wm���h�Y�Y8h�c`��$��/��n�b�W��zAE[4�7�vW9��Dø M}�}���Ӈ}���E$2��s�>� W���O9�իW����}�U6���.�� W[ۛ��=�%Ƨ�f�Ӛ#uF0���'���^�+_]e���U�:Jց�NtD3����]�O���o��߾G��rI1`�ā{y/R����3�1%�m`$-���q���Rа����5�v�Gw��l��נr]�5뀁�rf��j>�M!�m7�@�
l�"���ש���)�ҸX��Z-"jf�6�Ȧ��ӛ����Ͳ2x�3���G�� y�E6��	�F�V�J���I�	pZ��6����gK��z���&b!�iB#p���,�:��>��,o�₸���5gK�����o~��"�%@ܪ&�-Y��?�6uT��Ћ��^�����l �+��.qD1�ݠ(���}��*��8ڀ�eZ5`�I��n����E�!�`��I07\i��0��F y♋t��Q�,r&��7���4��Gt�YW�Я4���O��̑��?q�>��3�v�ʐ\<$j[G4�em�A���ݦ5��B�D�P^��X�� ��r�N�Z����.c߻u���k�E�I���G��d�#���M�^��ʐl,Ic5<�z'�I���H�����sg�N?}�O潅`䎁 �p$��j����������j���k嵾�u� ��5�|��2	.v=�ޕY3�vOB�s��]�ܽI,���pI@F+v'X� �2�N��g��Dǎ��/;B�-��Z�ȍw�6�FK�ӳ1�� ��l��:	��%L�-���Tmj$<�'�|B��p�	i@:hn~��J��y�}7���ӟ�+��<��%�\����B�D���9��͜����~�XЋ-$�+�c5�74��y����?���{��f}}����{\2���Ǣe�POd�軌�s�л�c�_Ĕ.�I�[���!<{��n�7����{,�&W
~�X"5J�fAN9ʹˠUK��| �@z���0�0 �O�����&�$"�.lU	Ч{M,dZn�g�{���W�:&F����~`����KK��3��� ��4��F��
���ܑL;P\�v�N��E�$�n�:�$��&�7���饗_�A��� ��f��[1�k�M��wD �?��%ޫ�-��u����`�Le�_�9�tC��?�3z���FO]z����6�����t����ޥ�O�3/>G+G�h���}������[t��=�������nCs*0F�d׼?��B玝��z�i��'�ѓ�_����%������P�Ǐ��C��� ���Bӷ�t��:��C��/���:�@��A�+��Z�G�|>���)�L����n2Vv���H3�m���ʅ+J����A[�b�=^�9�ӑ��ᴓ jWW�����ǳ���c�mB��P����@�G;�L8�h!���z�V�!��4��\�@��~.A��_�c����uN$`$^Y���^峕��rօ��pɪ�5/���G=��r�TRR@���8z�p�믿����]�Z32��d�߿������c��A���4�\���d�>��O��)������ES5�)Hϕ*g�*���l�L�V$^e_R�Jf�f���o�ܺu����Za��	&����ݪ|�T��\�#Z���F#�M)!�k�|�)��w���#8F�p���a�P�n����#¡}����k�hw�M )�궦�US�b.4�Q,�κ6��1���ڊ H��\Z��C���wY;����}��BI]�VL�Ib����A�4Q4%�>� sE#������/�X���0/cg�Rd��!�0K���e������
}�6@�p"�ch�:�d�R�� ����1�6��?u./��Lv�n��6�������`�omn3�j��i�Z@��{J+��h#ht���A4�CH͛�0 �m@��6ƚX>�B�:�5�r![Z�Rf��`�|���A�W����G|�"�%H�'O���ë�a��%4E�*��d>*)�
��9���bkM;��7����6����B�pqH]�x�"���k�?|�N6 %��H�Ź��Ws�s/�H�Ο�㏟��jD�ܻE�m|C޺J��o��x���o�j�YO�Z�ט_��cڼ7���>��F�a�ܙ�t��s�}����;t�;t��a:s��?u�N9F��83R*�mo��ƃ�;k6�z�)	]�^��WS���!�Y��@���O�3�>֒�"P�o�W�@���R>���g`�+��D^?m��~��&5͎�>K0<����ixg<R+����.LZ;}��Qh�	�����L�H�B�d��d>��U!I�N�ҷ�Z���%�s�m����C6fXG�?�`Kc���N`��@�fz���Z��	�d�բ�P;�Þ�汷gϖ�:+'�^N�	YCt~�l�����4bM���O��=���'�Gt����������0�N(������9� V�?��~�����պV��:2|ۊT���<D~v�X�GQ	�"�_����i���c�U��5�1P�aa�i �pa�U��ێ�Z0�-\U�2����R%�,�S�`�j�\�e�_o���^��O0�������1��#5�M@rC���օ�6ѷ�jwk��g����тK��B���C7��$�
�h����ȰF�0�3���ML���VUg	����ya�RF�S���sqQ$�"�S������D��I���Y�F�k��$oZΊ����ӃE�عϚM �u6�âfp 8�|�gY�Ij6�iN���mi�[���y��qe,�QB+#�_�ݢ�?�>��o.�s��9p?�8`�Hs�ETk�?�Vm6kdgw7i��ڒ�ǔ�&��;�B١<��m�To�-�Wtk�\�x]�h)��.F�1f{�.4P�N�������l\�X�6�����(,���b���~�;/�������)�i��	���A#��
4n.r��c�p�0�h@����W苛���f_6��Π�a	��٠�k	��RAm~�n���;�tkt��lܢ3wN���ݯj�Y���ߺ�FwlpYa��3G��j�8��Xpx�W�6�����R�Ց�k葃�t�@E�#G{WD�!����k
P����|=���,�%��ws�~̟s�������UvY�7c��Y��f�Mip�v,m�6�F��B*�c��(i��ƙ/9kbp���g�˚­-��,�Ol�f՚���I1e|��sm�|Uμؚ�n�*Ī6Ep�w��S�+��tm�=��� �r )��|,���m�uB��fEJCW��}z�'�ȱ#�J��ԩ�v�wv%H�ȑU����o��3�������w=-����+��ٍ�d��K>'�A]�Gim;�CwL��y����H�E~!'��0�̈�&��$��n��ZI�~.�`C�b��p�@�#h��06��X���؀߆���s< �ɫ@/�鹍��ų')�P�<V�k�c?p�e>d7��0b�>�����g�=�亮{�}��9 ���(?�ٞY�������ff-�lI��H�$�S+�3��	�nu7@H~�P�U7���o�F*`Yƀ��2��� �Y9W�?:�0�}Q���m��;s��h�3��<�O�yJ����	�<�6��8�8�s�`n�� � ��Is�����ߧ�Xq0�g�����M�3u��	��l�ݻ��죩��q��3�c45�M�����y�̥�� ��S>G,�Y�kT�(|ZE����)�n�3GH��o}'`��l���^ �˴�<`W����ـ�C0�c��h�/6���V'�m�gt����8�~̖��K/�K��J.�H�p���V ��:���ʑU-=�ѕ{����W���������i������r��v���ϳ �����M�s�1�;�P?�{+¸L� ���o��nn�f؛��g����	:�axޫA��	����L����@и�$�Y|��Z�|=��3�g���5�mf�5ʗ�d)>�}��l�+������*2�'���E��k�tG��렃�n~��=��g�}�G]9Q�'�����X����npU�ns���^E.=�(�����������4�/�]ۿK?��W~�\���u��.��ߪ��+W�.�>Y�Ds��_k��Ɗ��˴��u7�6�r�f���d��~/�.TP$�����7.��l�X�0�g�}ʱ�Ν?h�+�`��y��	Z����cd������르�{]g;n�,�[���⤙�N�
ғ���8TI���c���Qkl�EM���@!uҍY��b�'�U�p{�V%�Z0qbpQ=�8�	9u�9:s�,;��Bʟ0%9�@�#~��Y�ɹ���19究r��81��w��K	�kڏ|��^�ϩ qّ��Ș��{��'��r�&pT�s�m�>Jc�H����l�q�[}n�:�Խpm��8Op�uJ�"J�n��%چ�*�kN��@]�� t���:�W�S,��k��/��R�R����15����������i�l�������fn������Ssұ,f��1�wj� #~�R��3-}]���gkQ� �6p
� �^�v�� ��ϟ��/r���gϰ���y�}�.}~�2}��5�ï��:[b���+*6��i��mH�2��RQ"��6��h������g?������AX�y�axݧ;��yx? ⊎OЗ��L7���Cz0ۦ�r�����L��p��U����5d�6nI�-/1]�"5#�)�}{:
��i�7`�7S�( �;_|��uzx���O9N��x`����t 0��'��/��]#����S��������.iMSc����F:d�&:[�X��)����>�geׁ邷@@����wwy��I@�"!��rI_�Jd���L&C(&�;T�f7�m@�}z�M^ŁE�,0�c��Z5��_~mގh����:�N>�ƾ��Ε�R���<7}~�OK:6�=��E]�τG�S��iS�K�������A�/rv�r�J /�ib�>d���h@�r��q�3�_l ;X�5�hwq�N���ѧ�}F7��`�����b己��#z�>���)���Wsy�w�4D���N�IͲ��$e�5�Q��e�D�*-x@$��;�����sB��bm�	~30WL���!?�ׯߤk׾b��8L�V8�I`�����`R�S6	�!���������V�p�b/$�d&����	5����L�x1��f*�M��{b.i|	�M��3�&Ƹ ��` �H�`��2[��f���Q��Q꩎�ۺB���Y^������ᐶkd ���]޿A�.]� ��h4f��L��5���fB�j~�Yb��*�nf��V�����@Ԅs1�T�h�\ITK+�b�7
�N)�qN�i2@R�}�>Űb@�+)��Y�G�}tS���tL����:0&,8���,,�|���#�?��Іop��-zL���r�3/|����"?�O>����X;j�a	?MkbQ�rč�xq�G�m�Sp]����sz5��8H[���N�n|MWѾڷ�j? �	�?ޡ��q ��K}6�r�g/��U/�}�
:�f�iTj��)t�p�����t�U�-AX
�����} ���l4�u��K�Ћ�/��'�s稿:d�q�3��W)���J4�sl��~�t>���Զf�fİHbL����[/��\�d%3ߔ7͵O��H���O�͎���t����X��X����%�*A[9�,��?��,�,~�\�6�����f���iL1>-ޛ}���q�K�ۡ-�zi4Ja��ZQy�i��T��q���c�wMѶd�}�jM�b�賧�c_e���&W^��%X��+���}��]f����o>dp� ���{�+J���/~��l��B��U��ׂ`��q6����S��ִs"��~/ͮ,l��+~��e�\h���U�k�yH�r�j)Us�#�M2�0�I@�m��ś�'-?��['y< ��߼y�*4KG�g扳0p]�{�6O�����]�1�u�˨�ѥĘ�X�<u������)@���J��2� hu l�bb8�z66�A���i?�/:jc�y�	�����;z�磅Ϥ���)+���w7&�n�}�=�j'�_O+��9��jh��U���aM��H�3�\��L���]  ��I�[L�X��D�3�RE9j�䲐^�~�撲���-��x�X��Z�{�ڬ���ZJxoboඍ�^�4*��W��i��]9#m� ���Hµh������*����� ���ʕ��ɧ��?�#2�����=��s�����|���9 ]'����p �W3/Ay ��N��7�y�~�?���K���Ck��77oЗ�\������:Շ������`0��A��43ߛɘ�^�"i��Ă�1Ϭ���g�/a�� ,�S�u�s��)��܌�q�m�l�v�Uk�p���=F��YS~��y�{x����5(P���6�V6�]�$��L`Z����'��r8wm.���9ؓ������M���^bB�>��=�2��p��_��]4<����qjF��&��v7��;+-�K��sc(ک@ǂn�7�b�&9������%��/����-՛�e��
x9rK���IK�IҾx�O���3���G.<�/W���{8�kwszh~��ᰪ�1J泱f��$��\0��-���i���;ߛ�O�ŬQ}�k̥��Va�E��Y��V����b&5W~��Y�,EZ��H��\�:����<�GVx��?��b��v��7��?����=�6�&,Iؚ�b��46T�9�'��	�Z5
�~��W�2M�ҫ��&:������H`����Z2$���yƉ��<!��i��q�,/�2�Ea�a��x@i\�k���Tr�[}̀�w�K/����?��?�J��g?���������=�q��o~�k.,���C�"��c�"�/>7�d�J��S�B�Wη��+S��� :s���D�FyI����c�?6��X�g�CFc��H��������@ j/^��xD'���/P��`�'�l|����Yz�'K��D{��͚襡�i'	��G`̾�k���|? �{w�;�4�^�?9��zc G���&�ƹ���ؽĄm`���b?����<qy��>�H �[>��
v5E $��9|8��.�q���ьU�]N�[��#����g~i��\E� ƀA/�Q|6Z�(_}��ڡ��{Ի-�őAei���� ���,2M���4M7γ<���������_�x1z�h4���6���+�ӵ t�?�u���r��td��#?��0�cfB��2�h�a�-����C$����tH�66h��͐O|6�p|��OP� x�O�0(A狭����?g��ŋ/���D�y湳t�����+���Q���'�t�%h(!ŷ>4��UF_�q��ڐ��C��!�r��C����,��98�Qh6kT r�qX�s��}�k���1xk>Tk*ĸxn~4m��]�Pr��0
��b��2rPb�V�_NUٔ��h��Bk��G�|u���%ӋA%�OJ���>h���q�$Xp��:]�y��}�� ������U�6��S{�#gֹY�m~��x]�	 gBG�k"Ҭ
��˶��1ߍO��
��}ZF5HX�!����N�]~��T]"��}��):~�x�;\�7doB�����֌)��
ײ��R�4Q0��"K\K���5�k���ݲZ���� @x��Q ��  �ؼ�<j��BE@L���� ��0P� ��浫���@��`�a-"��"w.�H�G�7��=���ko����}ί{-�A,vh��v$ ]H(;ʕ��A����fGK;��'$��c'�UJW�b6����n��['��&t^��c)���ZC��q�u�6kk�r*���T5�DI�����(�ww�ݥSa�Ng�K7iR9Y�*�Ď:���:J�]j�`���b ڬ� T1H ��f�%B���7n��0~f�M�/�^�<��[��Sm<I�p4�/��j��t�@Vb�k��+@14���Μ�&\�-�����A���_���< �۴[�G�D1�� ��0ְ�`�<x�0?�0ܿw_b	0��@��7��$����W����~��V�F����`��Wf�(� Ĺ ���w��X�;��{x����=XH��mWAX�6-�W ��~�G?�d[���>T�{�G+�%:�r�����|�@w�V�1\F¹��brZﰆk��o$����f~`vxf��+C��z��N�z`i�^�޷��>
B��\ ������^V�1���"uOw$�(���.Z�q�2����i*�����s�#_�E�+/���L��{��;���pt{ѽ��l,skK��l�3��Es�k�$�(V&�F��ҩ
k=M���z��H�|S�+~�����\m��)�]�+�<;��՜*�A��i�S��'�BZe�����켿qN-�[k�͵є��X!�&
��`�����&
�2ĺ��D�]�bϬ8*�8�	]O��Zb�PS���P^Ȱ�� ��R��������N��9��I���S�Su��f&�֐�I��(�����G0����3`rz ��S$��?��C�8�Ν�a�L8!�~�A`U��}y�Kfҹ���%�"���?��L ��o�a�ekkG�ah@�~�{|y����!�lQ��IԢ)G��Fv�C�Lr��L0�V.�/�ejV�U osʊ��4�17��b�E�L~$�8�����Jn& �~�t���͵`[(�>���p�`�Q�Z��2�X��/���-�o�i󢹗Lʧ,s �	�_'S��4��b��swN��-�=F#�G�7��	~F��&�$���/7r���6j�oʧ����?u_�o�sg�p���A�4�t+S�j<fRE�	�K��/�~�{8�y�G�������QMLE��B
�XB��BT�o����� tsg��.��hg6�f._
{p�GͲ��Y �;�*��B3�Џa5���
 ���:���.���)� �9	��F��pu3�J)�ix����1$&Ghu� ��|E+K+�uw���v�f2�a�f+��S'x����4׾�J��E���RP��O��������)���Ͻ�
�켜YFK��g�s=٢FE�Ze��	=
=������%:�K���?��Xd�Ӓ���i�	$�t��;gy
�ʈ iw���ZecFq���9��H'�qו�)�r �3�����Z&L��>?�*��e�ۈ���[j�����30OV%��(�j��4t\Sq/Q$IA�U�]�:
P�ڗe��T�?�v�>�7Ө�;����f�I��������%
@,>�9X����޽����� p���tnݾI�� �?��ooo����=��n_�������:���K'O���?���_ �#[���	�AD7�	��#��;�N�X��������4�Ԛ�<��b�?3�i�X�;�TUlf�@>�ZϠ�80 ���t��-z���{���I��"��`�j5"+�;n����1H)�0IB���j&�X� 
	��-�,щ��%�=�>Ϣk�7|J�����<#����T���3	*���r�S��&�=��͝��.{r_�EH��tT �X/�5lϯ5��{�P������vW��n�D�Ï�����p��	vG���~�с�h�4�[co1�V�7���5{%�aWA��Ճ�l=�ip&ܒ��7��B{eb\x`��t����;����L�=Z���}���Z��0 O�i�s`H~�ǅ8/yT��y���T�`��Kt8� v�w;�
`�F�Y�B�Ʋ���r� �y@�6�-�(��3��S ���	@y�O;�^��:�y:��):z��U����x!|����p��bsYd%Ӆ�O�ǮN<ғ�L]��{*�՞l@S����z�s&Af+��K�w��s�Zuʚ�cw��l�d67��p�~9�@e�J�{���n&i�����j^�z�a��]���y��ոN}+՚������<��j�fy�d�۞
:�|^CA��M��f��ᔥ#��.�����jvr7\|r��sv�&��%��R��)�&�����W�K���\ $ jF���g))3m�iă��F�qv�=%b�+c��lY{h�#J
Hť�	��	p�6"�n�>�cf� ��e��O��  ����4%��J,��G��T�;[h-���K�ɜ!U�?��*Ӂ�`����9o�`�~6��g�whɖ�,��'B��)
�)  ��A@@:��~�x#2��[ �^g���I0�9��fn�JQ��T�U��]��[�];�Ѽ�"88^L��J�;.�G��)��\��]��V)8<+ "�;z����Dt�`E?�2�g&�Q�]I�3"!�	��HK4�nU[l2����riތ���N�G��_Z_ʣ��ܬ���[�B���mz�ko���9����p�B�T|�5+ 1�b,�ހ���4�v�(�	�A�a �0�#���i�G����
Q�wh4��JX7�"���]��\��ju�XO9�E=T���?`w���
gm@m����X4��U���{�͋��0�,:|p��\������믆{�ؗ%��?kك@�<�`5�B��@�%Z��q��-��F17�Ҿ�-r��<�̞�k�̗2�T傥�%�����CW6����f��V0�k��{�L�w�����¨�C1O�6���rV>~���5�撐����ݦu�r��o��U��k�k�$)=��2_~�&Z=�_��n=}�=�&d� I�"���a�I��q�u(֖	bF_;�)����������_�ϓ`t�VO��2��@)�.�p|�pM��	��)�+X_�p˘�)�_�����]��vMe����@��Fjz"�?M�Q�3�ܷP�K5)`���8x�(-���V��yx͏Lj�Ob�Z߹ʙ/۔���� j�p,�2�����108ԙ���2�e�49��5�n�����&��|Pc5�g�w0k�Z�>h�O�5��'���/�K/�LK�<�a��UR�O/>��M�Q����=D[��ۘ�=J��8؃A���Wu8����)�e �@,���a�h��y�Vx��R�h�yϜyN���A�8�e΢���oj
��f}��v:����OJ:�����jf��}�]���7iE��j�\q�5��Ei��$�-�#�ď�-j*s!�R����D4��s�̙{�ڣ5���uz���n,L�>�S��6\��l�����E����n#i	k�dm���ʬ�u_k�f{�3���t�����!y���{�+t;�,ܡ8D��l�w)��A�',��E͘���i`�9���G�&C��.�� (L5�aE9�����W�þ��/�gl9�Uc����!�Rh�+i�z�� ����;t=�σ�w���CA�Z�^�/]���ӽ�d�͌�Z?2�����t-+�r�:���c�K��w2a:e1�gF�R��C�E�(h�jtq���}O�i\��5olN��K��2���8�_�ѩ�2�MnޯQ�Y���a�xT	���b�sw5��r�e3���a<�l2�j��o�P�e�i0a�o�q�ACf��������w�#h�Ԋ�@q{�F���2@���a��R�UU���Y~+�l�+���JG�96��jXk5����Y�z�=�9�	��?�/igY`A���h�����m�
0c�޳��i,�Z^�u����w|�2.�K�tb*ǡ�`}X�>`���C$�����o���OK=��׻�τ�FGH���j8�ڡE7.�/++��N�^�}=��ɣ�0�"�͙3gX[�NB� ���`�]
�dk��Yc�a<���F�U
��_ܲ�Ġ�AH'�����g������vj�ԧ��'^�����I�[�?im�~��p�q�c���5�x��\�U�Xj�YD��(�Ł�A���DMgΞ���y�^{�uJ�UV+���^K���J��>? ړf!p"�y�*��	4�ͭ�˲ 8-��5\�oB���f�.H�3�@�F1� g;P?NT�Ki�D�r��az�����.����B�H>D>���Lk�ći0X��X��Ǐ�(�.E=L�akķ_��d?c�$�	�I��`wЇ����¢#ȳ�.�C@	2�li��J�A< �7�72mPzwJU\�\,��.M!��@�Ͱ��<�ˉ�� �����Z
)�ڃV@
�Z�$;;[Lx�;o�Ye����>M�y!>L#��Gf�/>���=�ǥ~] ��A��w��^�*�7�.w��ta�N����4 ʍ&M��p}M�UC+>�a�`���^�k��R�Ac��p���B�C�k�W�n&�'ẙ��:�,���&����'���º"�^���7^���n��п;ʰU3 �x�,�ly�+��/k�j�4��3!Z?�g�g��w�[�kҞr����-���6��|�5��hq	���>W٘t��?q�@%������׼�l-}��Mȫ�˫�{��us��%AÔ-���V/�;䚗t�>�S*����hyi��i�M�Z
�51�겖'�k�|Y������Z�Ul��W�XR?$n�h��炇�>�t�	�	��$�'U�l�&��8�fs�{�'npq~���\�,e�r��؋�-�D����Z)�br��z�z:k��Iq%�\����J���sKvo����4{�
α�nS�6H�QfI�K�!��7�u:���d��b�VU+�e�%�o��E`�e4"9�Y.pK�&Pco�]�L���q�����E��i�g�] \�4~�{ߣ����\�`E��Z$52�� �H,� �/����߸�>������J�j��t��/Dg/K�:	}��g�v�w�	L��7h�����/�/#/��g�o��m�|�a�m2OD�*=�4�_蒎�rW�E����L1�.g`W%s�,-�����C�.W��Ba��3`
�hcM��f��,g��%��~F`�t�;� ���lڰfZ��P�MU�B�Y"�)EѰ���#|/q\�7+�a�J�-G��O�=�`/3s�}��w�$pv�5�frmP�9����T��t��"O�L�KI��3�ܰp3 �v�̥�6�yM;f�կ��.E*�ao�Eg:c������2E�V*�%ׇY�r؞\��+���
��Z��Mzx��=ő���sa�m�]�JhR�*1��.0�����5�c}�E~�h+ �>��{a�p?D���_��cp���@����Ӊ��|��(˷zzv��zt���]{���y�`PD� �v���3;|��*FiM0�������
����x�%��{�d��Jy^)���;;dSv[�n�e�;���@6���8�8&�ս��f��3��	(6>+e;eA�����z�n\�L�� �~?
�uVL��T�'E�{����̘<�{\ܳIJf���4�x({`��4��7,ra�"�gc��mI�gY�P��Ճ���<����-���ۥ��Z>8�*P�[��i��h�[/ fӂs��L��I�C�	����O�M�G���\��D@��.j��]Tj�d�۴�U"�_]D�IJ/;��a�\�Ϊ�9�9��)�9D_h<A���t?��,f��Q	�"۫T�I��;֞�_�����>k�.^������f�Ń�U� B\u��u���5��/~A_�5���?�hnm����E`Z�ۂ��� � ר�L�'���7P.���(>SjaWV�36�
"�����I%��WE��Ib�C
r8�F�kh�Q,��:P�-'��&����L@C���EC�@����Z���O����<��S�x�)��8`n!�#ŝhGDSm�j���Ji�8`�=������cR��� dN1�R�ڱ����*4MY�d�>l��6cH~��:��K����X��EX�U��&DE�Ke�
vg �U�M�tqD�wNF��[O�������Qs4IP���^�Rs��L	�Ĳm�x�(j�����E����铜w r@�$�����r�0�ʩ���#���ن�K�����R*U�~ W���� �my���Q�0�	��Н��h�p51�Z|$w�u���������kw��X�lB0�n��Q��$)�k���@�g�9?��A�#����l� ��Tk�Ś�)aZ�z�B�	��Ulb/_'��\��z�h5��nؽ�L�j�{�ϣQT�� hn��4؍���m�|��k��)E�?Xȸ M�\��ǞO��r2��X��^���G>��\�|�D�Ҟ����֥*ݍ����2�r��'L�`^���S�3��?[�Y��MO�i���.���U���`?|ﳊvN��$z��q�1p_)�� L8��%!�h��JH��h+����
U%�t&:�Uհ��E��+=q /�����g|Ǌ��*u613�� {��o�x[|zb�2�.�`��,xf�(u���i�dv��iz���������`�,eh�R���A4l}:s�t ɇ�7_眧 � ؏=���v����,
�$\�r��
w	h�j���~���s^_�	���ϙ�޿�7��K�Q�b6�QI�:v��>8u�ۋ��L��ْ�q 塟Ќ����a�]��Y�,�V�qY�ZR��H��Qy��.���ct��3t8���|@5,�*`E%R`Zz5M�r�͟�H�8�
s�de�����"J+��F��/�\.R�cL�!��yq����//����8q�N�:͟s��v�I�֯��'���.��m��8Q���TIJ���$7�2�9���Y�? ��/�x=Ćè-A^ƃ��YAV��7�L4�Z/�L��ց�2*a�#ai�q>�u�N�ӧN������=x�k�H� D��
�8��W�>�y�V�Z�N)��ς Wh٧�I�װ?e߹��th��ӱ��k\ܘ F5y�TWcW���4���@G��<�`M��ڌF:������R�|�:Ӳ�q8J�i���|YShr���)
�QP3��5+
ڪ=j����ȩ/�Y�����qR�^��o�C�-Hs���k16�M�rqL|�,z�ڇ98����k��&��I�����i<�@�]87Uρ��sP��s��~#碻����돋[E�SeB����M��ե^���{&ڍ�r�x� V�s�O���3?l���XMhURե���W�Br�ϪV����98����t�x�iU��5_�J�o��X��D�����~�k����1`�;�kř�y�Q���o�͠���_�E-5ל|�rQ��bF�y��[x*
o������z�.`���įL,�� l���_��_��.����A�X��'S�����3�ѫ��B_|q�5�y$5��w�� ��) $@ۿ����Z�3L�A#�6���,��������	�ɤ�'9�k�̙���������Z]]�r�X� �w�ܥ;��������ȀZ�F0I0�CPY��ٳt�����+��
! �Ǚ����:�۵v���YX5�Q%$ҽ0��)�GC?[��!�aKC�u����w�R�YZ&�	����{���P��^��D��`Kb�߃�D��Ž`�y ��Ɋhv[�ǒ�
6M*��Δmz����Xr�ܰ���F.^����_������͛ao~C_}�����L�����m�ۄR!�RQ�kvQ��|����TР��6�qta��)�~؞4
�/��G������s7��W#�ɀ��Ýz��)�[��cI�PJ�=.���C�"��`|���DM~���\W��dΉ��H��R���]lW�d�� zb�&�Y�.��֕�G�G��1TU�gZ���컮�.�B@���!UX�Ə'�-<k���[����A���G]=1a6
3ڧ&���U`3�e�V<T>�8��Y�D���T���*�+�e�}*��\��Zi�{Pj$�/'��n>hߙfsF;���)SG1o�e.�5mS�Bki4C�Ղǜ�J�D�o�ߘg�9�9([>d_[�`yy�gb�}ދ��L[8�A�*�`IG��t�o��F���$<j��-�E���k�i��݋Jx��	�=�	7C����0X��ş�����K�y�� 6��" �JhR�H �H���7�I2�|�M�{��u�z�2;�@��Ϭ0��w�9ޠ��mg���+/�L����X�Ë@�$OzxG۠Ey;�s��/ S3L�HYe������d��$��4c��^�X L�?>����U���Xr�2�g��%�g|���V�CO%�:]MZ���/)�z4	����Z���P֙3��̥P���4��kp���q�|]�)N7R�m4F�U/_&"}	��&�r`�5  BY/6��Z�[�p���5<_�@�;x��;xp��(XY�Z�0"�rgQ+9�g��}��*DJ���<��k0U�	�r�l4�\]x����6i{kK��-PG}Ƹ ��k���N���7f�~�'!��Ahڑ֊_@p����!�Bk�-�ѧ(���B�=���?A�֥a
>A<E>�PxVj�������L����z�%*�F�9[�/�6FR�")���o|5�S�O���(�ǒV�������Y������h�A�`<Gm~��9������e��������� ��j����
M$�57�H#іs[�X�c�ٵ��x��e�˂^��{ꜚ�x�-�#��ꌖ�)6�� fm,���+2�h� �G͵�9s���[{&e,���>{����WA��4����=e�f��� ^l��b/P��N�����&h��tтH�$k�HZԴS��SP�����/3 *�3���q�2�M�!�>%)ݸ��j���rŁ��5�5���h��!7ʋL���5�Y8la4�Lh��L�	����Y�m\�2k,�,�[�9����ժu�b��<��Ο�����0oޫ��������p�"}�;��k��B�|s�>��#VdN4��s�@Sj��ݏ�E���L�����Ћ��6y^%��V,��`� ��Ņ��~�}~�<~��m�"�76�x|c��/�CH0Y�� S�˯�>e0����ͷޢk׮����p;���@O&)Ϡ���ĉ��_Ǖ��{�=��ƀF]��R��S);��������7N�cۓm-@�Ȼ���Z���Sӿ'�NZ5�Yo��!��i�fV��Ŋ�2�G?�ty���YWL����ɂˑ0�U݋�@J��)�}V�Ģ於�s󚄧9�9]t�BӾX������\��=���17�9��j��]aK6�i�)Ɯ9��h�;�ju� �>uZ����M�d����� d~��3���l,����Y� ��2�E�B%ZL�I&n0�� <���90�\c�McB�BG�{�P���)��i<�s����Z�貳�MA0`P&�}����Kz���>�\�O�A΂��")�֫ZRQ����������2dE֐����0��U�7ƻ���9�k�Vy��%�|a��j6��H�j�EO*!���9�w�ܾ�NG�Hi\�X��v��h����,04��u?;�1�6��'�6�t~�L������wo�[Y�"�C/�и�)�}�az�l�g#��,#�'�޼h��g�3�U*����c5�Ax�]���w_��c`O$�2���+�Iv�q��`�M,�	�X`��Y�L��`�˙<<��� �Uk >ï��d�������S*Ƒ�n�v�-�C
��(��+Xr~�<�Hc��{��s�OR��1�zm\�C�9��|��;gV�x��n�)��XZ���R'R?A�f�bN�g󾩻�.F�'ch�6�K^q�<J2NX���T�"��k����w��vUw�>łf�� �9�1����{?���z3`�+�9}��_�rF��l�w�]���ϲ�w��r�֏}�1��W��Ck#jl񓰇���#P��u��"�п�˿p���7��=���K���C�ѥK����� p�P{��E���?��?��q�w��4���f�>��>������7����o�I8�=F	b5��# ��!i�k����GY&8��J~9�9[��ef��a��^7iU��H3��<���h��[�\��x�ݝ$��K0L].	3�lkэ���wX�_)�N�+/ʎz��s�2�>��_1'N^%�!�=�<���M;���`��V�;t�0�!���X�JsJ6h|]͂�H8#�E�F�g6�5�6��ݒ���l�e~~�7M�x?#�FH��J��1��R�e�8!�ZܼM{�f0·�{q/����z��;,�޻w��/� �n��6T��j��i���Q�L���;�id�yK
2o�'Y�+�B��("�D��y~5`���wu��ǐs�Z��	�Td������Y_5*h���*=��b@h� ��q��,467��u@�v���W�V?�̬/���;+	^g��, �8���9��`�tG�� Ac�70� xf�4�Q�/�v��*��2Sqz�dZ�X>hi���o�2�4�Ѡ����\�mE�eE������L6�����"�i����jq�D��@�P1�ݏ|�rz����I����%Y��}i��m����e$�e٨w��j�8��9M���ct}����/�p����$ �/̇�<����?��������(��i�Wb[3 �n;�=�n�ʥ<�Q�NO�8a���k�Vb�&���T���pB�����
8��6��DZ@�w��?��Dk	\���P>�i4y�Q.o�i� ������0L�<h@���E[ �=J�.^��ϟ�sa�`�{��a H�ٶ -i�KmV�0����O#�Y�ń#��k���f�@��M<� �	K7��5%���0WѪ/�6am��"��Q�sbۤ��R 0�rX����Ҩ8v!Ҏ\���0~�y�:C0%��%U�$n>�Z���ROsՂ9Ls�caass;jRqཱ(zno"&��J�&벓+D3h��#�;���y�+��hyr��A�F������E-�!��AZ��Ge[J�����#��1��RRd?q�S��Wߪ�!�
	�9#�k��:
��ٰpu3X����z1?v��m[LZ���U�bS�xk �dQH�$�q�lA�P�B�g��+}�iv�V��l�I�XL[8c�����ʋ�tY�lDvh(*��n\:?��h��Y�X��;�Ǐ���U���]ܻ��+�C�tO\��I�*�����A�ǣG�ٷ������S��P�[��7�ͪVe��p�TC��~�p�u�;�]�9�Jc��G�y�T�`��t��݊Wd�/3�d��nSO���`�݂ҝ-ɂ��W��teQ��n5rƓ�Y��Rj��پ�����ݹ=�.|5�Ǘ��G�6/��X�	� YK
3�?��n�a��9R��t����Q�=ܘ����Ds`�GJZ`1�W�#5҂�v��/ï{��ra*��TiV]�l�y�$�B�O_�O�t�}���O����k���5x��H�Vh�f��>��Ο?�~�8��B���!7ϲd��x^vKZB�M-@/\����g����u>��8齻���:�wl	zss�5.�Z���(8T2��6�y�F�n��+�/Q�yy%j]Ɩ�`�d���%����<� �����J 4���*�}n�$�����ޥɘ'Z�nOq�1��}�*:�o�"6ek��8�%R�����_qZ�J�w�X8g�I���f833�h��Ŧd��8��a��`�&
sK�[��mr�Jr�\ǜ�\�!��wE����e��bL��k��Bb�$��4�)ڎ2�H	�T·���eQ�g��˗B��Y[uaz�텶��A6+9뿳�Q3���Fi���`��B���0w�����u&��+���w�vG1Z��ָ���R)��)��<��k��W1Iφ��vRxF
6ʕŢ���r[�1i���*}WY7�h�7�F�����2\���E�Ka��ܙP��N�ƅ�츏�>�� �}�R-����������ϥ�F������x�Rs�w��3��1-��N���X�,���]��i�s��l��j�D^�A'�C�M�Wio�|�o�^���M-6\�;��m"��l��o��\ަ�E��.�ޘ"QҙY�T�Ÿ���Y5@w  ����x��d[؞(��L)m��-s�p1V�
�����8��gw1q[�H>�҂�����R��eȱ]�#Bxe� $af�8X!��(\240lh�Ξ9C� K�VQJZ��-'ο'��Ǉ��N�	���f��6�f���.0墲�R`�U!���ok4Շ8��[צ�m���ӳ��=7����p5%����o���&����M�y'��.�_Jrnh�Y�6�G�c�]ڐ�V[��$�Ρ����%�����F,	�W�T�����چ��H@^�&uhl��nI���啥�ގ�o��{��6�����{�m���R&��� N���Α��#�ٍA*�-1�9�K�&��wk�~Z��MSK�����{��0baX�[�o�g�:OЧA�@w=��_�q�s���j������B�h**5�i%2��e��٢4Ы��?KYr
Ae2���h��NCM��cz��.#�kV����F��tl�}F�k�'�֍����e��Ȩp�I(��k��J`�����:�7c�۞���XmH�����IF�>��
0�VwF[�	ċ�C��W�E�&9+�
�.|����'>��#�J
s��$�_�ܚ�Y6�2��c|��{Y��<��,�zP��J܍��o����;����\�(�ZOIs��s��]��e�G_�VK�`�P�t�k	{�ֆ�~���C<eᑻ����8����a�?PV�i�����y��_����p=�%�Vg�p�`o��Cy�8���ԏ�G�ԺH8������Ӎ�DԔ�����W�J*�����ɇ�E�-���{��+���s縒�� ������ا�t10\�,t�ח�B�5>2D�6�k��f6�y��E��=LG��*j�(��u�O���Ǥ-Z� =#I��`�\�,)��EZ/�l-0LgH��[ �N�$؜rGƦc���ה�x�H�Ϲj|���>z4<�>3;h��#c�9/_fN�0�����h���=|D� �,U�ȜO��Y��^���,t�,�*��܌m��t����0�-�+r�,�1����A�n����ށ�)`��E���5st<�q��+��{��s>���Z[]-���we\�4!�	t|���Q
t1s�ܪ�0��,.�@���y���_Ϧ$�9 ���R�8j�-
������N��:ZS��usyʆ9�}��L/��kvQemQݐ�k��To.�d_[�}|�b����h!��͎���_�!B�ƁUڞla��� kaP�Y��"Cf���M�Ո+C<�(k�gpA��G�`]3�o�2ˊǋ}�Q*7����<B�h�(X�\�<|'������(sdȗLא�~��<8W;�3;ǿ�$/qkL,��T��E�]��=�P��I��Iu�G �R]���N�6þ �=�?���a0�v�l;���=�$��?�4ӎ�zCh����+"Wtxqmʇr<kի-�,>�5	:d|�(��Y�R��E��u��&����.���J��LNՅ�2!�"-I'��OԲ�g�*v�_���˖�5�r�8�Z�����޾�Մ�r�"#����M��
�F�=�s����0+F�������<�����,�@���E�3a1|�j9�BGN���u���V������1W����7�zg�/��ށ����p�M�^e�H�Ckk�e��Y
�2ޙEdw��G�F��JN.&;��f��X�1�s���'��ī��J?��O8�����o��\�"�y:���������
����G���j��ļ�A�����Zb���{���sg���Έ'`�T �?x�]��!��D+��چ|�$��[2�)��IU��$�p᧾T:�����zƀ�F�I&͞����T�QrI��7� I'�VW<� �[��pe��m&��gOs��M%A"b�p:)+F2ki���R��H�;���?�}\��v%��#Qb��y!��ڀu���}^oKvd(��ڴz�~ߘ�y�R�{������}w����V�����P� ��Ĺ&�S���\b�?I�Y�"ak�\1����3���}+�9kl�U�沫ͮEt+�\ǵ2�G?Ț��bK���Ǐ��ܷ.d�^r�[��Ʉ=�
=R��f?l�G�yC�*�p����1(<�Q�H�ޗ��ڙ�&�PR�)���g��d�e6��UK�{_�p�f2�z�a���O��\��7��O��u�k#�a�r�*��O�,��t�e�js鳿w3/����V�^�No���q�=�ߦ|�N��r54g	�k~�Pg}�u0��#ޣ��FW���9�8�ܺ�L{j��F�C���7h̀�i��pR(V�6����:n�@G `!�E?�=�O?�������&~��K���&��{� >ۻsn	N����~:���7&�Dͺ�x~��V��0��f���r��[��xO}��)G����֦/>w6�0��d]/�+6b�}q���1vڀܭ�@��Hx�X�lm�-�t�
�\LB�p�����_����O���EY�S�����֜�\��������*��k�v�4O]Tb��6���;;"�97f� ����e�R�!������ǉ?(��41����W_�.�������<�|��-&b�ސ�������u��C����{����ʐ�AHV��ؼ���"��S&�OωDԧE�h�a�Z���ܮ2y�׬_3ez�s��,I(����
`wn�b!�fxY�
�[��z��¯����Q�#~'�\@ӝ�l�*.l�m�{��T�w�Ls���f-HC����`����e tŴ�����
P�1sT29��	��Ɲ�FG�����x�=3�x(0�_:�~��QZ7s�!�u�R=���;֩�%�Q�!�ˢr��]&�'9r��v��MV�~A8�Z^r���7or-�G�'xi�&(�j�g'��>��a>PJ��1�x���{�aP[!�n�Ӎm���l�i?�����,y�&�����h����.)���dp2�7�tf��
�!f������^ N��>F���6oz�iz,y���H�Q#��ǜ9٧5� .���3��fز��a����i���`;�j�7�����)T�a����J.j1�K~^�drl�\�$�����!��rL�'����-O�p���˗9��&�$׍�R�s��u�����N�W]eQ;mP���Do��`�Esl��M��-(V�S�+�޵5��X�J��=�ʬVI�R�Y'JYx2�(�	y���_��>�ӧ,�!�]@�R�d!u�[f|z�l&�kT��K��|h���Ͽ���vc��Rۗ���bU{#ɶm#Y�4��������3g�pd7����X_̚l����Ƃ�i������/J&��{��ӕ+_0p�D�&����ZH�x�.�����
o��]b��$d�F�l���i�wL��2����Ő�V�d$A-¨�dOzL��V��Tsl�`��Vji���Z�?�9�L� �;;[Ȋ9�� ���&.-N��iǺƝ}�4�i��y��������P��hqQV���N�M1M(6�� ����,v#���؟�3SrU���T�Af��|e(&�w1Jx�m�,�q� ����<�5���g�0K]��=��y����ȹE��=�\Z��X�'����c� ��A��|@p@�&�����@7���l�>���a�&�Z�E
��>_���f`8���㶾E4�aO!.tZ"B�6�ӌi�i�Nh�ff '^�� -�m9Ϋ9A�d��K����v팩7m��Ct4�SokJw�Ocל�ǂ�@0�csv���g$�F-m*/+�C]��4a��L��Ch�>�sB���*ʞ���_���D�l&(7����8c`Ņp#��ê��*����%�Z3~��r#�u�����Ŏ���9��F�3�U#�����+WY�sB.��{L�"��V%za�J�&t$m��_
�Q�뒕�Z@���:��R׳]���1k�� ��7�o>�ge�yʕ�r̩t�_G�<�}�[�S^b�@O�Rh���=
%�7��ǎ�xI���M�L]��k�]�X�NORHqj�K�K��@ c��}�������B�Ξ9�)&���f�����ݽ�⋜�%�a�?t� �Y��s�6�����R��,��X*w�
D��?g-ۍ��$�<L��&nP��~s�kf�\��f�%r_���2��5��o��k��׶'ń�Ꚗ���fR(�F�NL�#��;��!$h �r�lZ���_�U{W�9`�l��RU#����U2�b�I�QC��� c��2g���OR�	�X�����29|��[�����"f��/���pE}{{1��{E�;S����/����K��;D"��9��D�����D�ڋڳ莒�nF0�.�*�FX��PR[���4�u��i�V��&���)H���:7���3�v�Q>�+��~7��� O?N�}��hv� ��>�Ym�����V�{) �fK��R⬭r�����R��[h�U��V�mڰ���i�q�y#��ܤ�~����*A��6���1���ʔ�H�N�qP>@cnLj�=C�����#�\���x��nEE;�x���jvm�u*�
��X�$u��N�{��ΡLR���Z����0=�3�Ed��`8�JF {���wu���r���Y�%�����Qw1�Fr��*x*�G�eewv$�G�\�k����&	������a�6@�����;`����1OgZz��怟}��}w� �eji�9���(2�]B��\�q�GZ�'��-��ft)3dbϜ:u�����xP^U���ܣ�aMg+�+�f�n/���c��z�L����%Mh�a��(��Ue�>�+˴�ӑ�G�շX{��6tMB� �E`��#�آq Z_}�5�@��la�.�(*t��x���}���O���05���.L�������ՔO���� ���Q�/ZI�Oߵ���a���%)�n�migl ���K_S5w2Qof�2iD�*Y���.�`Z +��E����N��$�/���N�3U�o��|C�{��[�0���ȑ��E�]��=z<kc��2���O���lݔ�fP������qۻ���uv��%�3���|	���E��MM�̽��[�C����_.5H����
�!�n�v�,0���b�c \�x�g ��"��9�O��i��`�}��j��..s��!�W��	�
����	���
r���R�a�y�<��-G㓯,k��psP�����
�q�@�
 �&a�L0{�@��ȶ2`C��~��A��Y�݋�ހ��`7F^�$����C�T�	T6��SK�-b�.
�ba�O��2�Jg5 ��m�d��Ca>�h��~����c�{���Rm��\%����=��5Š�;F�%-���e�\�=j��Q3'O�8�
�K�k��GoG�w) ��۟�j�V��Y�ɂcn)8�îb�Pts��ŧx��a��������s�ե��(���"R'����@�ֆ��tPL�7�rŖ���C�Z��e�U*�r�X���:�XB�L�A[���FX�����-��s�S��eRZ�6�|�f��Ս�B�k��`��}&Zo��#�����k�1x��s0i�Ұ���4<c�x�=r����8����~6����bɼc�Ok��V��������3g9X���������Ga2'���ݸ�x�9E`Mc��>G
{���1-�ȳ�!ۂ٘"w�n�ł]+
7.J�:��rfxnZ2mA�VN��TeU*A!��5�xJ�R;Mc��]X��M�6hN,�Ȣ��:)o�~��10wsj�0�h�L��&�{��QBgI
���"����WL�����@�Zk�.����sf09e&���c1���\a6E@�T)�����C��)�h�T���&'N��/Z�^%�_������]�0n�A�C�h4�MM$~�Ut���v&Y�"��i篸��}���d�� ���at��޽�s	�<�-�"��6�SBۅh�p? Vv#��L�X��w	ƃ�Z4Ҁ_+���`Ma �;�p?���2��<!�p�p�v X�a�N�z�G#R�8�H��ϪJ�rÀ֙v���|�,cП0�%f"`�PD��截�@��5�߻�oң[wh����A�a�[a��B��7o�v�4P����cv�MyZh�u=Vzm�iBc�i0>�x�	����''F�Hj�!������[ߡ��/1���s��B#�Y3���)�M�o�����H[�*����q��gAkM+Z�|�2�^�󷺲������\cX��,�p2��g"�H�E�mXs^�kKPl.Z�R۶C�S;�%������N���[�4��{�~a��Z�E�E�+@��ìy�´?����J�X}�,c�*�����-ڹ`�)�w��p@ ���������ϱPt�ҹd9�ں0!J���省$�~�[9u#�� o�s����0[Ʈ`��b2E���:�Z�E4�0"�����>\,b4֍G�O���������{����o����?�?~�G�|�ָ��u/�������x����5��i�p.�s�^�ӧ�c�T��/._�ˠ�����HS&U�~�q-�@�=v�)���x��`�F�,�D?���>�c��:����V�|#+oA�v��ZN�=Uqv1&i5)�-�61�Ƨ��y[�|]*�D�*T��rͮ�Y�cք~_	�sYт�X�+�3�d��{�f�6u�qs�&ZG�}w	7I؉�����mZ[�K5�qv�E#��3���kEi�k�S�Lߞ�uQ'u8}J n/O=v��{�4]�t�/�H�,�+���d��e�L��/��T�D�渎��Шm����~�� 3� &��l<�a�`����o�д�R��Q���z��b.>W�g۷���0��`�Ť��v���������[A{�tm��F ڣ��!�����&m>Zgw�E��}:��b�q������hګ�i�Jn5p6N{ղ�:Gi�������6��G�]]�3�&T\�ĵ�jc�n�<�;Za.I�[����BW>��S�4�ˊb�4+ST走���A����]$#L�L�J�U�1$�2�lmp��M:��^w��MH����b�����=�����7*��ee���3�/MyAi���ba抛��!���u�5�05Řh�+Ͳ�\�V����(aD���+W��>���;.����A�:v�8�r�p`OB����cU�$��My�OA�]c`���6��鳛�M��w'sR�e2�h\��4�Z�DŭR+�y���\<|��'�CD�|w�~����իW�捛<�ެ���w��s��qZ	ʙ�m^]Y�ܿh�T@76�9���f���$��i��0Ӧ]"�"@��8���7�,�:���1V&���#o�n~e0)7mw}���f:�&�RC��e�>��f2���[�%�_L��!F�g�h�,{�s��sQ��'�'��0�,�rU�4%I���q�#��l�ܡa؁0�8�KҍY�$�l�ŗ�d��!6�쉿s��F���l�2� ����w����L,��*W0��V���6XD��o�vss������Am�Yj#4��Ep^{(�>�(��8|w%rxD��2��TG��x"%�Ҁf[;���y0{����tԀ�3� #>Rk�k�Qtk��ht׷h �t- ڵ0�#=BS����M�7igc���0 ��'Nҫ��B�A8�����L��O���h�Mx}����|���Ŗ8R����
P�k�^�7�������1�7m���ekm]�7r���#�'����`W��6L&��~00����w˭��@�bkKMyf�'9��7�W��n��/�+W0�vg�����rv��os�瞦hz�6��}��Â�rpi*Ue�����v�\3��P�e���7A��*����^��6)p�<��7���?�뾼r�3A0C�a��pq���_���\j;�Kv��J}P�T�&}� �d�n�`!�ˍA"�SbyD�m��y����$�!��_��G�c32�ZSV�`���Axn޺�Y������W�����k���	ϲ�.`��[A��C�D|���c�m�f�>�@~��)��~ċ�W��E��g�=����.}��%�f�ӧ?8u��5Y��rJ��kь�U2��f�d�m�R��&˨��qj���q�׸xLH�}�žhI�]�����h��\w=�'�6�ֻ���f�Z}m���%���y���fښ�EݯV7=;� �!2
�m�l��.��b?1�Tb�R{� y=S�^������w9i�nT��8�  qH�b}��h·~}c�-D ��y�8 ]�YI�kv��I��:?��CѾ�ׯ�r�+�+�u��%�}�ݽs�9�����@��ք�X^���٤��ôt�(�]n�=z���(�\�T��$���bZ5��� �����v���;4 w�p�( ]�ئ@|��5`W�� �'�6�8�Ai �o��&9v�����ܢ{�#��W�f�Tֶ��|�[�<ёӁ�	�ʈy���>"���S�T�E2��`9�4�H3e�di���X#���ͧw��)
��Z�Կ�ݫ[,�W��~��ș!z$��{�f����VAn�9���V���[֗��4w�as�i�1�(nRq�&h�,j#��A`�}��ό��'H�"�]��)?�\[�Xv���!�f��eA�LW���-�o?�ۤ�Ss	�ݍ����eH9k�ļ��Y��y�K77 ������������' �by�魷ޢ���g�F���V��<��Z5ħl����g��EK,m�ls���������s��?���K�}�̌P��R�
U+|-	�H�mf5��BK�A��d�Y��
jji�H�+�zZ���'���Ya E�$���'�D�^��Y��y4s��}6�PZ�-FO��q_�S,*��F���6�%i����m&��<���E��/j��\�A�mܥ��h�Pl��Zծ>.Zx�]1�ujK��e�&cv�������x8ďw��3���{״}�s���U��e)�G�4��.Z;L���D����e�(8Kg�G���'_B�����5EmyZ���o�oA*��`�ṛ�;��B/�PX&�]� H-2�� SQsA��aZ:�	�6,L��0s�� �_z�Ev�@.���6�[et���v����i�δ
 �^�˻�n���fu���ރ��@4�1����'Lȝ�o�GP\ pL�oCdO	�n��M(�E��Zv.�]h��&4��qF0�Y���	%]k������?:��Q7���]�UN�8��b��*gP��u��a� `�ʧ�e�6>��򠺤Wc������fB%z�5��V`~��+x�$�OtE0�����H�ք���}�����}�@;$�jM���њϵ��[FO|筺���߷�Y�9�{7��e��k�K����&x�����qӵ�s�k�Fe���.6�yI�! �i|��(~{��?�}�P���.����s���Ȓ���>�U���>ot�?ɕr�l���q8[�:��V�
7��ڢO?�����
��9��=�.�yQD��Fc��7b����9�4?�] m�4��e�a� ���;��1>�t%����Kt�ԉX!�B�W_}�n����a�k�dO���%��
! w��D�Χ�;���s��*MY1��Ǭ_��&�5�ٙ+D\�.�"䫋�&Nu�}�6�Io��9��o�_wj��_�l�_`s����ר���[�]�8�k�V�4i$V4D�nf��F�,W� ����(�� ��(�Iqm���� ��l"ኾ�Jp�$�t�B	���WӭhjkZZY.�򠽕�qf��b�M�"�U ��e�.=��Z=ە��ƞ����o0k��=�����A��f��L�Ʀl4�YamAH�x3?AP�4�,�����[� ��C;p_��Ajn AD/\��N��O��[; ہh��J���2q��{������R����
�����`��	p���1��0�z��@K;a�o�5��?�F����ｙ�Փ0�)�Q�BP�=���u[Z:{#��\�Ε��G�����h�4|���ڧ��/�>��N_�����پ'2�~Q�Hf���4w%r鞑�X��gHW�*�Y�G�|�Kv�TB����.Zx�Jk�0ٚIZ�4��/�`��<��`������RV9Դ�Axp�7V`�I���i����>#׼>�3��n��{wg��|�>���Poه]�`�}�~��i) �T]�4j���U� 0+i!wX��A���T�Y����/�^���)s�\�Z�a�hT0j��gQ�\���a|��K0Y���Kt̈b������&o���smrw�3�����ѡV�.�F��_�B�����$|Uq"�d�3�:{TE���~F��C/��3TI��@&I��@[��Ͽ@���}y�2=~�Fa�8��=+# Q���K�g˱�q�*�l%7�ԯ	GsnHՔ�	�h[M�Yj����YP���J�r����N��iו@�3}�%E�$�6�}b��X�.Ɇ�i�3��F|�v��i�0 hݰ��ل)m�ߥ���ɂ�T�".=r�D�j��7:&�˴&����	t ��qSM���_:}Xh���4�܎F4, 0(�{LKr���:F�od@�5:w3�c+[�)�uTZɫ�q�Tq�lƼ�@��~�����,�"㧟�����r`�����aѶ"�74pq���K����۬F*��4���v�&����b�=x@_~�=���ľp�y:�?���������\�U�� ��-W�	�\«O�01y�I��ǡCP.�h� �C�����)kVA߸�2��gN�)�p[�L�?EJ��F�}@0 .�.�� ��o2�e��$|��<%�/İ�t�|y% �[v�r�+��|F�Cdp��?Ds]�����S�e�[��3��ˁĿ��l����O��ԍȢ媴���� 4Y����K�K�}^�v;��q\Rץ�*̻��4�.Za��>��	�����v)�g���3���?`~4ݟ�B�86@�/���Y�5vQk�m�\1����n�_ �������{Z���s��K�9v������x�m�(���*�^g�fԴ�Ҿ���b���p�x�\p.b&A(��d�	�LG�v��sKQY4��=����K��YF��MŒX��t�gy��X���L���?� 5@ʿF1��8/
K���+t��@�3��pͽ;w�굫��W_Ӎo��k̒ �4�Z�h���/h�N����BS$��裏Y��ر���3L��
>{7x��޽CW�^ᠹI`���m�G����}
�i�J��
�r+��Հ���e�FS=Q$P�&��&R�����R��Y& �׷I�7xk�V���`JrG1g�x�p<��\�g�sȘ�W(�L���ܹrqN���2+�U
�Zp���S"V�&��qlo��\܃��i��\������iZ0{)r�תnu�
"B�v�d�Tx���:3tҤ�3Χ9Ľi�+|�Q��]8a�R3�f��=+t��_�ʇ���������h��Ї~�h4�8P��{������I[��A�ϙ��"�����k�ҙ8��,�� P�@ܧ��}��.�놶H�lo��L�G�C ��N�n���3-��)�Ma$�s!h��Pu��)z��w����pe�A	*t��즱��f~��g�z"��]֨'9��=�%���WM�L����A��Jn���*W|m5���@3��fL=�J�s�����pyI�W�$<��鷭4r��o�Ɂ��h�kbOҬg>��ψ��6���k��hw����Ez�:�U�Ùw�\�� &'�l�R�=��y����8���V���^{=���������μ��{r(�Yْ���+�����O�s,�l��)JL I �ar�W[�U�^��@�,��G6����n�:+%��n޺ɱ��� ��E�㐂�EՏ���S\Y+���F/�Z{�`�>�Ϳ�@���&�p�"WG����W_�H�s�α��ȑ�<��>�=TJ���� �B1	�Mg�4��D{�������S�2��0m~��u6�� >����^z��t��k��O��lmmpB{�zI�b����9�`�ع��O|�[�s� �3Q�IE��EL�\��]Z��t��u�Zk��Z�L����{���+�V�$����1s�w���=<m�äe�3�
R8"[d]s��%q�hgT\;�,��3��V��J�k����ZTu��/+�$�Ƥ�;��Mb�VW%�u�k�[bv�h�  �s^�ԭ��V!%���+�2a�2�D7�s'�"�V��^�_�\�H��}:�ӎX�ބ+ B3h�!�60�>�]p�H��>������}��\���_��߯~��y"ԟ�L�.�v����K��is9
��/��鋝��P���i�n�}�B6�5��W��ړ�s��m|0m��Sӎ�Q �
��?y�Dj�E9�<[ʰ� 0�� �"�31�"?�L���vn����[�NO~T�g?F���cb�mA=ˊ�7�p^��_��*�ż��+vq�y��Fֈ�߸�]�nj�ʂ��������&:lq{K]a��R�#���4��3��M��_�9��(ݘ7Ĩ>���ت���ku�l��A�h�k�M���ǭ��X.�ϳӅ�^s��w�`�%������#��/��>w��<�6��i|�&�� �����W��-UhwY9k�3Ϝg�*�^"=�{|��[������Yi��K��T��}�J�d�Ӡ�6��$��P�S�0�>s�~���_}���˯��e�`V��igg�7� ���St!��/�D��\�7�|�>��*���w�����ڽ�q�b�D�h�/-�xÍ'�t��m�}�svW��Ѕ�ҍ7�K�߼Kwo��9j}�K1��Fw�(�:O���E9�R&�����QL#����N�R��H%�"��W��۳vܕ&�G��.�d�3�Q6��f�鄁Ƙ5�^ZM�S������~C�-kf�B|
�	��9����eӌ�$Agf��dﶙv���Md~���j=�j�@��ȉ��! �C"w��DQ��%^��C����� �a��؜�y;�aƿc��)�݀?���dS�(G�Ms���\5���A�S3���% S���Y��q�5�ѣ�9ͬ� �����ᚗ^�B/]�������S��*Od���/��ޒr���H�H�v���7�|k��~��HW�r8pʝ-��1�(`w�;�^�S�.�F�4ٞ�xgƮ�t7�����*#��L4��� �)�/���"��=dƳ�>�/}�%�|�2�>�>�د7oޤk�>f�k�պ1ִ�f�)�?N��z��l��:6Si�&���Y��T�
�H�����#ۣ�eK�����N;�+m������y0m�Q��4�Ҍn� }�M�L��A�W�l��г��e7�L~NpAON �>ZU� �`1K%{�ar[+&hT`Q��$'�z.ێk[�����]������Z�r�U��w�=w?W�.�}�ϡ҇
D۔��J_:�kȁe����f!�mo�9B	�K����ͷ��$p��0M|h�������=��'?������ }F��!��OT��H�B��^�YƫLy�۴gO;Z?B}ھ��Ǿ�ƛ����#.�{.1��Ą��FP&�Q���.�Hu(=�9�/]�"W.�Ě��������t��=l򖸪R�蠅�3X��5�!q�o�	�� ��+�VCe���`��0}xPl�9�C�T�o<����߷��ZX7?�XJ�s��@�UD����.�0�Nf��������o��������ǗY�+�,  +�����O:����5��vg7�]���7���j�m<�Z���� |���p�o��.�|u���b0`L#!lR��옐;� �kN�/ۓ̹D��b�=\���ž��O���q��Z�d��	�@������|�]6��:��I�ԭ��Dv#d�8s�,[�N'a+
~���G������~|��>\�q�KI��>�~���c�]�j4�>o��$�<�`�9��`ʃx9��7L�i�F
z#k�cv[�@�DHK�R����%�����h�իWi}}C�v�5|�����S���u��i�(Fz�D�i!�wo0D����5[�V4Z�-����ya![�
���3G�'��nZ�|��xm�s�~2^�<��n��v�R�s������
�Y��r��U���)ݻ{��H�]Ii�R웬����,a�ߧs�f�h8�֡�L����*��un��Ei>p����QY��{�%�b��o���}��ߣ���w�BB�.-����'\�r:���cǹ�=�c�U���v#з��m�u�&}�٧���:�P�3	 �ҧgcb^x�EN�����OR��v��yz���g���]���?�J���J72hH�@y�>sVQ�5������G6�K�Xs�E,�fmԸ��&���'`�#�3������ۜ9tF� ���/���k���7���P��|}�YK��Ǐ�9��t&7jXQ�
=)�i��µ��6�)$��t�c�UAsm�Bl�2�͛���f� ���bŨ��.��z3i��^�]� ��X��}pa�:ĳ�; ���p�!p�99����a�3���Ta��������$h�4 Ahx��O�(C�^a_���s$q��0)n��M2����D�s�yA��.���Y��������]���J#��S	��?xpA��'N�����*k��8��n6+���=N{��ߧ_�����@�8�<}�_�`��Ϧt��=�Zߤ&��A��	t�RL�Df�v"K%�n�L+�l5����m�<+�ȧ�sw�^H)ఛ���M7��J�>W���I�AN��ez5�^�\��`l��>���û��gׯsP+�p+�Yc<���� �A�+^�ؽup��W�	��2�4??��=�T~�(B�_ۨO�
G�tm�q�B����T�Q>T�+e\���C�-hK�b�`ل\*��6u���R�������g�K��[b���_�dA>�S��t-kɷ'����� zF���EB`O<��_o��^<j'{����	�vҽ���}ߵ|�5����Z�o |�H��5�p��w�VK��H��w�}�h�������$E��T\p��	N�"\�dc�Ҏ�W%u��~��O���� ���׾N���w���3��z���A_x�u&��	|���:&&X8>��ʗ�����Z$Q:�7��x��y(����ko��	�K� � n����w�G?�!���ÿ�ۿ�����6�6y(�ڜFm{��S�.�o�U�083��Q$�dUWH�l��1Nh�$ ��5�r~����K�)�*7��s���I� �8v�_��L����j'�fH>�~�h�
���
�ΪMUh�hX�(^)'ƅA��!�̓�T];�(��q�hH������f�0�8�얒� n<: ���7�(k���cܐm��*�kE3i�FՒ���T���[F#Zl�{s{+k��	��t^�d1P�l�w[kQ�f�e��&j�hs�.`)k�k�̃h���16<�p#���e)Ћ6�K�_H!��%����g�=��^1^�*.����9�)�[�0n�u����x!�~)Ѥ�y� Om���tc�.�?X�To��S[�9{Bb4Q����Y����Ƽ!hvI+�c+�ͼE���i�A�m�$	�HM����!:wF4���ַ�}��X �'��i�(��`1��8[䙶�Xd��c���&8k J��H�rrf����d�R�f�U���E}n�����,+[%��_��f�eat��ʮ34p�J�V�n�"-���<S��Np{ЁO�]���� n~W-��YlL(���d<��Ѝ�v��/(t#��|G��~�M������J�y�X|W�moͬw��{~��6t$��׻yu��}��W�O�n����&�8m�>���<���.�N</kbl�X�I =p�	C��J��θ�7Vȩ2i!�͠g�����?`�P�8��0E~�o%��2��on0�CC��{｟^�q��G���?���	��|�z��hz�3lx������_�۷��ҹ�=��{�36m��x�������|�KLL4��� `�N��W�df�����Ȇ���QR�`�#V��dqv���2P��m;��"�EJ�|�e�,R����˼��d� y*9�m8l�K֨Z�շ�XK�3���k� ��å��F;�/	����cC�]��R$�ί!F�}�D��`�=���H}Ӱ�F%� � $�+�:b�d"9EE�M�E��/�}C���c�Ǣ҂;����io`lp 4�a-c �,��`a@�--�� 3�b6��s<Fu�H���kk�Hc^�E��z/��nk��̘bߴ1iZ-B� X!�b.<���+�+iަl!A�0��Ej5����M��~.���+�
��U��_&�a�`����~˥�/���1?r�(��֛t��Y:������k���g����6�Z'���:s�W�hC�@B���56浹�sr*�eD)'���c�-u�7�]K�^��F-\]಄`�t�K�M�����7�w1�j�u������#�bf��R'.��Ҫ�Zۿ���2��2�)ƅ?��r/��Fr���3x@a���j?� ��CD}6�E��W�Y?Ř�5�=��	f��ӦB��iR�\�^����[����c�t���g2(`̩���'k��`��;u֏G���C�[$'���3y����"a�	 �ȴp��	�KnQ�>d�ڿ��_9�rj�=�^���E[��ǟ���>˩*^�5z������_�;o�#�s7gn�a�'p죛�� 3�~�.�� �>����8���6rUnm�ǟ|B��}�+oqPʱ���B��	u�-4��7~A�0Z�5��$���\�Q|]�"]�I�nD�3 � ,��@t��Y�!�@�l�9*ߢ�[��+�X�2h�'�Ji�����:��8^O��3\-�Q<N'8��և-,��t��oE�+@C�Z��.I��j��ni��ϴc��)Wx"���.p!<�;����M��d�fY��5uUm�̘}��`v� ���$�S���O?岸�q)������� ���j��4�V�q�1ǆ*,��c蚕��R�X��<�N��%-� �r���I��YX�f� >�0�Y:��	��^}�C8�e 3�'$cŀ��>I������j�@�W?��;۴y�>m��H"��O���M
S��q�^�ѯ�ճ ��FZI�ZI��H����5�>ڤ�q�I��@�ċϿH��Z�����n:�Xಀv_�z�]��(&ks&v��>n�f<���
D���Ʂm3����ϳi���=���<#��W�w휉;7�I���YGӽ��s'���3-va����ŗ&��۬�����:�����ѫ��Q/t%�����b�44�����'�˝0���l�S�����$R��]#�������a�`՚ ��qa��|���1�/���~3�;�a_7����ݜkD�v��eM;`93K��	k�nܼA��������Y���2W��+|+>?��:�L� �|�"��;}�k4z���X+��

8@�4� BH?m$���^y����>��} �/�Ȁ	��ѣH�=�l�xv#)pP�]��9�6�ywws�Dq�P�m�`�P0��Gs[��ƠaM �^`�H# ��E<�$�vdmM7[`�k�խ�eߡ^w���,��-Ym��iC'S����@3gJ���W�{?���`�}�8J| C ��t`�c��:� �@����g�e�5�	��u�m�߭��'"p�
"��ML��KA��" ��	��'���ܼ��歍Yˋ�S���7�A~to���r�+Œ����ըn�����*�Շ����V�g��gdD�$	�	���Z����A�,'O��ʏ_~�j���^E�?�:z$�Uv?@���/��[�<nii{J�1��쒒 {���܁NÊ� ��Q�Qn~N����O���t��K���|5���~�J|�������o�G}��3�=*cS��q��{�P����=�;_�Q���ڪ��nv�l�����=<( ���w)X��m!����ӟ��s&��� ��n�g�x�R�J1�E��X�_��t��Ϧ�+���y�Ds-t�o�9��Z�����J�{H:�C�=�\)L��q%�:� �<'сe*���a��r�\5�@`w���L��\�m������`�|���?�ӏY�M �[��H�)�bB��v�����	�r^�W^�`�S	�^�t�.\8�fE+��"*PP�� ���&$��3�'Ѝ�?�я���[�������f�Tp C-��=��|�g����9�IM��\>�j��Ϥ=r�sd?�r�G��0�<���e>)��dR�Bs�@���ϓ,0S|���\�� ���'�!W�1�/CP�{�3	�G��?aS@�Jb�o��&�css�6��+������>���pxuY��׸��1�5��=�p��;��S3Ɨk��Ѡ�݉��B��'ِ�S�.�ًT�	VK�*��� fX4������=���F�MvY���~����޲��13�2��
I,L���� �6\�P�B'��B�{X� ������x\ 0b��Gk0�L#��� �����@/�/~�r�kﯾ�*�:s�W,,6'0�o��WX[Jk�׿�5=��m�]K@�v:�,k���5y$��̍ |�y������mml2�|�������_�c'���K��믳�י��si��h,��p���?�e���˹�����ǠOt����G�O@�V�O{BD�#���u8��,k�_�o�"�ܿ{���6�ᶰ��z��i�{���&�{xw;��Sk��dɇZ��\�$������9�}M��g��@����w����1#8.?-��H�c��g��߅�����D)��g��M��n��?̓����׮�'_cs�����%6
��1� Xe����уG�ߡѲD��@��D����% a��L�"�?��SvM@�x�3�̼�@4R�@�M�ݻ��ʗ��	��U�4d�]�K��ޟ&`��6ַ$���!r͐��8e<�-�+D`�"@-4; s &�F"/14�0��>s��`��_t�K��$@�\)��p Q>T�6�i�0_���_��	 +�b��cj�h���vTJ{P����m$��vjs����~��v_d����]B�t���p��j�%A��f��8�<L�i�2Fќd���nJ��ͻ�����6Dpc��I(C�Z0L�f�S��'��4oǓ`m%��G�Mk�R9k���:��(c��mN��&}�	G�?�� !��p����圯�	�;{VRƥv>��ԩ3t?�Y=p>|R�3?H��.�ь���X�y�P�r?�`�����c�+��=F��{��g�--%�%�����ox. ��C�*�����6y�X`KR�v���0�6�L��h�Z&6f�8�����[��h\����t��W��
�-�����3>��}��<��T��eV�d�XYmm'��ۑ�ux���a���ԍ��_�g�\�3�Osy��t>4����ɾ� �  �����j�f���6K����y���E�Ҳ-i�	�ϰ�<'����s�Rpό��6d[-�Ky��S��m��>�Zx��ȶo�^�kaZy]��U���Mi�
c���=_��l)dy��
u���jp�/���|��W���`��!h�`߯��J�� Y�P����4�?q�<R�˙S���i�e��s�c��]����6tn]�ˏ\���y%�"�ؙ�J�C歾��7���͵�3��{��w���j��Qi�c����s--�\�w�3.��e���n6�,`4��7�G7�TS<�����2dm��^��M4��>Aj=�)>�0�h�B�+Ș;m��y��q�0�A͙��0���#5E�0[��\�
!���F?9hv�A!x���ƶZ\=�"k>� &�������n��o��s�^��R.]��o|3��S�2$b����Vp�զ"3^h��������C:���
�!�m*n1� ",��Φ{@����t�	���,K�W�3f������uE��g��©�f5���Q�U�"uE�� e�p�B	��3g!��ӲP�8�p�������o�!k�%�'��q:SG�@Wơ�r3TzDjj�G�G�zkt\jI/e U��V�G@qS�Wֈ9l�<�%�
��mqc0??�_��馶`�9�,�.Ϧ-aAȂ��qYٔ �-	����7���St�ȱr>����!�2 �!��H\&���יx 1q@ R�E��Lm�,�������KTR٩�n9;��;\7 ����Z��ogs���N�I�5�tyF&by>e�d�@y�&U����҅c[�9�k#	#���}��۳��P�r`Z��fW�^c?⍇�iws�� �5�p*`74��d��*�(2����p�.����}����+��q�x ��е�?��9����p�b�ۛ�j���7Gs� �
��+����}�4�T�>zu�z���*�0��"B��"ܪ�`Gkk�b��5�S�׏�K#S���L-3<�8W�b�#�~z_����>��un-�^�Ɛ����̯CS�&�w�����Fо��}h��1�v�z��7n�s��ɢ.�*D������.8�X-�����u��;S�۸�
ϊՊz��+��8���O�F��F��Z.��N�լQL�s�tM����:?5g�͙e���G�ִ�ͣ�J#��ܞn�%O`-�p��$�i2w���F�6z������_g����wl�D�ZZ�� MZ�9*npB|$&N� � �k�rşEGS�E�< 0|d`@ڱ�^�����N#�G��	��AWp]@$3�� l�}1� �Cgh#���X0�=��G�'���AS��%[�_S��֞l�>$u�M*k�7�⇹;ڥ�]�;Q�0I������j��`8h������h�s����1�H`[l�[t݀��>&X�,9� �X��S4C	t�/K[ײ���|�v���Ok;�\f����բQ��{qu�%ˊ�3��U^�kP,eLZe���'���&��R�ҷWR�a��.��*3�0I](���$�M�Ya�	��� :�߸?��@������s�>��u7 s�l��p�d��&P|��װYo&'*�.�G�i�P����d5߅�cdMa%�v��U��}�+��\k�ݻq��As�f7Ov]tM͚�ym�3�4�������w��&��{��[o��Ͽ��9}�4Nc~2����s��/I�?���7����\3v'RmU��rƝ�P&:��5���|���W��r�>�@�o~�θ���j�:k�����P�j�k�}���zP�\@�&LS�v4P��ܵO�@��h }c��2 @-�}��E${\�� �,0VR�-�]^��I���pb[�4��O
!�>�B��3�A�
Ҕ �:����4{�������%���in�ܜd-�i ��D���v<ݼ>��M��M���S���Ɖ����gղ-=��2��_cJ
iB!��5~��T&�Q]Ԉ-�{_k?����?)R�S94RcdL��w(��?�H@��^`�^#�k�=�)����oѕ����8����Ec�-�Z̒�� ���������j`���}F���g`�̳����H�����~�^?g��$b� 7�S�_-� ���u�&�ML�N�'kq���l����e�6�R8c��hK�/)����U4�Mɻ�y,� <
�4͗���l8��`�r�b��3k�\x�i���4"�B.`w�yk[M�&ύ��=R>�N4A�����V�E+J!��͵�]���4���SȲ�xl%�]̌�Y:9ߺ
Ȑ_2�������ʸj~\�!e�����p ��~-ݜ�D[��8V�	+5T�����S:���F�1�1\a~���fpa@`(:T�_04��gW._a�0��H�ξ�e����i�>׸�~Jfc�W �z����>�lT�V�9�V`Q�=Kc��1�l���*=����2�u�'���&}���Cq�J�D��p���8��'�s6��;��y�ŋ���	 hp�gd\�N&9��gZ�M-���>zI�ߐG{(c�+�e��p`��� ������8Ʌ�Y��>1�t���T��L����Ӱ�c���|s�C�ܳ�Xܐ^�P"������}hr�׷�&�`�ׇ��mBE��0�����)�x۳��Gn~��r}�/u<�.7t?�������B�;�i{�k�B��ֲ�Iyjٻl=��g�dt�>����v��g�C���vi���1Kq `�2A�zt��"� � `���P�`�iK�B� $����ͷ��k�Zi���̀�ݿ'�X���Uٖ�3\3[��u ���կ���E�Q�����K��E34� N�|:1}�1�Eby-!ff����k�2s<�y.g����8��pF*=sj����Z�4�vI�/�e�jR�͵<��w��i1��@+ $4��g�dT&������E_�������"� |��#2�1��Y�e�h�\CP��̼��S(nY�U�Rn	':o��W*�(��&)���n;���� +�-Mz�P)p�59�>�L��ک�mZ,2��pC�aY�.)�1f� �*�h�g�!�kk
���>����\T�K�|ذ� �a?ܹ����{٪ ����[ռ�E#��y�k>��_�T�)��UZ�jv}q[C渘�j�j�Ph[�ͨ�����0:��fQƘsu����� ���>�R�]�@/]d+h�4W���<�i�b���@ȰL0��gA%=�TbW�]Mt�c���p���T
T���Lt��m��M�����{�@�i�B͟�����O���޻�B�uZ~7��՘��,�1V, �4������6�9Bs���5{Q�s��C��T��y* �p3d���2eW)�T"�Ѧx�=0hD	7,�eݴ�`W|��i��ъ	��,�U<���=�'��px�A�[Z�g��vr��j���[ؑ�K�~ڹ��\3kf9H\�"�n˳���B�L�k�i̩��i�⁒��ٕ
g>��Eh���K���� �I���� �s����^���'�x:�_2�xDy�g���L��Ą�[���m4��R�yz����M�e~��r0)�?���u��w��඀� h�N�|����yy��7x�36I σ�gT};w���>|�fp�
�T �Ƥ���%h�O���06|���t��K#k�Pq+��hK#��J!�e�
a Ĉ5��H���1s���V.��Ӄ��P�jh�h���5>��3ɲ L�R֒6@A!�������)x�k˕T�yd��L�[]��"q�Q;�4%��m�<�X��k�L�Z9L^r�2��L��	��HʴhY�q{���%�M�5(D�t#>���j�C�|���6kx�i0@�-1��n˘��AC�s�|�H�0�5��m���w9C ~����1-!�`Y�8�}X�6�&$d�pQ2-�L)�[���z����gׄ	��̗Y�u���	�]@2��۔�T���s�=�h�# 6	�/_�o|�����A�ǎsv�����}��]N�:�zh%����ք�����B�G��P*82-������c]�F���R��\#�\ �	4M�	�I4Z��=�Z$h�v�-�^s�r~g!v�n���mq=���,k57L��k�[%j
��S"�~�_����5��W�����'��be2��%'4Yr~x�7kxam��ε�5���C��i�h8�7�Se�*=l>�6g&����?s�6�'Z�ݹ�=k�|W����hS��Y�ft�6RT�O����|[)�-���n�&x����;�c���ZMa��zP��rg}n[���U_�l��"�= n�hz1����lE�Ps��9�m�ƈ+k���ڦw��=�����D�/�M��,���7�ɟx�[>t�Μ:�`nY�	B�b�Ic�(��ɠV��q�И�ӂ-e�ժd�����T��I�d�s �^|�y��W�ʦ�͍�����ݕ���� �k��]�q��/k0ͺ�ɮ�3�JP���QZ=�Qe�Y�ʚV�����V��6 �{��|Q�����
�r"1R�� �����8!"�Ĺ�g�G��CCx6�u�����G��Hn��Sm �CC�g�q��4�#��<�1fpƩʒ�2K�?�fkk���PZ�"�>� �I��qX��_��4Zt1��
�<p�(W4�G�f�H��0��?d��I,���x���������S�ˣG�yO�t	���|[���x�9��+h�a�8�zX|a�I����>�����il�\ p�%�1ח��z�?4�0S����ʗ_���n߽Mm�뱴^�Nn޼����$�q2)�Lp`�^x���"�4&i�06(�p��%��-�{��_�����E�k�!�}�TT��.����E<�3X���$�T�+`o*nU��XU@W֤j��jٺy��� �-{��Ήk�R �3�8h��F�MV�����9,Ew�|�i�p��oޒt��n�h��[�.�]�qFD���X�~����V�%���]jf�/c]�zF�s_>?G�7��`֍��U�̳�`[��H�t�'������N�:s�K,T�8����wɏ�w]����֗ZmD��9ō	e��,`��Q�a�N~�u� ��-�,$P���9%�T0�
�aʊ�Ls� k������t��1�o2�ב#���3��ݾ�e�/����F��ǻww�>MsnB��M-\����߉��6an]w�w�]0�m6�9iz�"����rw��{t�̷�Rs���;���>@�c%H�wq�l��+��d�.K[�*#���5�R�~:SlF�Y�G��ZU�UMT��Ϟ��gV@"&e�l<a�4����u�;Bδ�F���?p�,w��p8��&��/�?� ���T*d%"�e<l�O��P%飏>�4KYѶ�*�+}ǵZW�Q}��w f��﬒Ռ����wn�a�����M��w�<3E�o\������ v��bФ��0!�4�I�����#�HD����+ ���)k�`�F�Vb��$çش�h�U ���l9Wٜ���;\�c�U�Ӎcǹ[�,��:0�۩�x�mM� �)|�|�h��ڪX�]F�/t��k�'\!/m�go�6<��s|���h?�p.ڏ���{4K���/Ds6O��9^�y�� �|d�"���i��/��J��9q@?�����$t���7X8�9�gI ������$c�6�̥ ��3g���s�>�L����~}��=]���x�������Vܟ���90ycL��a�d��F���4�WW�\@�8��Sl6G!� �2����k�b�lҪ�K����I�#\�� �f�{��y��%�W���P���`�-�w� ݀q���ފ%���-�����n�cAۋ��������mcąh�����b.�� �w���������f�
PL�&�X�2�%��MO�Y ��#sݧ��_{�g0���Z\@���6�CJUSa����k.(�>ENm�LY�mW�D�mXi_Y�`��Zs&n�,&z����� ��z���V�BMWWC�^�&Qv��P���#�ˆ�m��@���7(����qi��.=�J��Iv��E��8І�[w��Ԣg`׀�a@Yֆ�W˾a��<�y����"�PZ��k��-��r�άe�px����uշ9c�[�_�^�=��T�&�z��7��U>�@%k�9�mlQg"����W6��O��o��I��1���c��'+*�a2{�Jeq��!�1�U�������E�$�)��iC���7w�F�|�P>����tJ �x8��V��aAI��MÁ[O��n�{(Ć�n��ԕ���>� �R7�q��#\=�W_����D���Ĩ�8GL���ށ�ݻpp?ђND�����' Achۏ�~�U�^x�E���� ���]�.�Z�ϴ�`����0<���G�hǽk�h��Nq��n#G�'Њ> ı�����<�@;`� �f�_����(L�]1�j��g�*DS5e� ��y��yje���Q9�χ& �aw�٤�$h*4h��˼�)� v�F��A��S���L�W� g".e�҃$�:|��	�j�Q�e����F��xM�p�r�2�:��~�>d�ػ��0�j)mQ��8݊ Y����&j&K큛�ի�ص�n(��LC���T�/����1�6�T��Re�;?���?�.:M��ʰ8�P\�W�wt͛5a��t���4�,rz'>33yq+Ѥ塭�<Q�m���@��`mo*f�
��x���S��ǜ�l�i!ֻ�-�g��E��ݴv�4 .,ȃy(38p�F�u"��i�ڦ�%T�(��=5�0���uسԇx����M�y>C��>x���'e��I�he�-�ϻ�5���*��vLhb��5��斄��2�����8�͜������M���x�b*fl���s���Q�W�3u��c:�
 q�hK
;��+�Q�Ҟc��U��L]���!���y��W�y�m������}�����[w�({4�T7���#�i���������/JA��`/�,����n����s��#`
�U��{�FZ0�,ZQ���!�@��[����g���LM{{���->���ѽ�n��̂���P�q?�
e���;＝ #@�}��ߡ/}�ef� O���G,U��9�}y�����������MOӒ��L�/N�o�
�������Y�ț]7���� R�L��x�ΦZ�v�@��/��m`���%�/�P���D6�X���h5���ӂy�?�4�:���7��wi\L��*%	�4�.&�2��6���7tFV���/9^g�,�C��o�gkg{���U$3�-�4	[�Q�DE��/�5�f���Y����>@m�VnR#ڍgA� w�)kfsfK�IsBY�B��ґ{�&7� �%�=�5����p�PZ�<��2$��n/4Z"si��T����0G#�)�����b�@��Ttf�97~�Th��6}�ہU��->�[c���"3[�#\q&�|��G � �x�]��������2���b*9xcT�]ӌkق����yS_�1�#��I!ziϛ�Y�4g< ��/(c̭ ���5��=�#�u/�4�
��d
M�iY��Djq�dg���D2~t�<�ƥ�}\��;�Z^�E��~30��0ך"�~�c+rӼ�Έ G>h���E��.�D%�l�H؍���W_9CG�:>\i[�om=NAx�M�5���֬�	�������_{P6?��-�g��(DZY� I��M�V�Ix�Ԍ!��X<	��$�w��Y^�VQ/�H�V\Ȭ�ߔ_�k��:\AKq��l�y�i��+������[	����Rɇ�A�zQ��M�6��0]��X�@�#�R��[�p`\�UA57wY�Ҋ���cyy9��y�k��͊$)4��\Y]�50��/���^��\��`��5��� �ao�GE��{4_���nU��춹�)	�������^��������c,Z�ڡ	�y�W��v�cr������t�`N�R%Ѽ�)�E���͜p ��"ͯ�3!��o2���X��$B�G>���;"�.��2Q�	
��;�/��N�B�{	�5�b��)����m����
MK��_hf���	�BCT���;��N��0�c�Z#0<7C39�l�@�AlS̜h����ܲ2MHN�޶Y"�)�̅���tIO&o�Ѿ;I��`���Ș8y�3�XJ2���r��I���c����p<�	�6I0��i��q�6)C,yfඈ3j_z�;F�������/LB�%|}-A�X%���$�{4�|ȥqG
�E+m�[�q��0�ݒ�_R_0�h�!XBX��+Y���X9^�Ǜ��e�8���2혽����K���^P\��'��5������^3�;�����Cdm�$V1�'�5�IV��P�;n��4y&*Ƭm�I�=�o��ar�!����νt�N��g��C��Ӝұ�'�t���GlcI����P �
�~�Ѱ���Rk4�2iX{�(M�B�I�d|��l��\���ם�r��),��y� E(%�o�l�z@��>~���y��St1HՀ4�k��47x0���9�u������t֮#Gx<'Z�ۂ�@�� �a�y��im���rə��w���k�F<��[Hz��ᲆ|N����{yP��K���ւi�֭ͧ�<�N Κ��,9D>���ń�F�[U�t�p 6EJTg�Ν�#)���zh�qLӔL�$!:8���{���
V����T*MV�r��y�S���(��)�eٰ����"vm�5��?�?���i�+��i �����PD���1Ý&i���p?huۙ.|c���rgȵ��L-^ ZU�HY$���Ee��g��UM�OF�SD̜ژ5�x���w��X+;�~6oPlXH��D�!uE������&)R� o��i:Ә+�D��0���śZA���` �)R�i����g��\�v�s�6j~�1���(�jf�b�������=u�2���Zh�l�VR���"�=(q�eo�0 �Ӣ�ΤK����tҁqp�H4� J�\  �',���0[�e�eBaժ�+�i_3����a؁]׺��k�������ۮ�����;��d-HP�4�۩�.����gf��]]G=����X�w��k���Ҽ���	��E�1
���|�.SJ�C�����by������������\z�3:�5j�-�X��Ҭ���WA��1F���`�h���{[{��]{D��щ���Ӭ=��a����|�BS\�l����@�K=��A���ǀ���T!".��	�b��E�6ZڤxU�u�!+Y�w�3�\��P��g �*�^S\���J1~��ɂ��}@�4x����&��+���#@y��h��i�_�������g�tWI�h�N��*a�<�v���wV�΋e -M��ےU%u��an�"n~��ͩ�Nq�4a�"�Zί�X�k)Y�����e-$�<���8���zڪ5sVk��>���w(n��~��&pzx��]�J��vQP��������(Z�{/˅���~��D��I;�qc(YC2A	��og�	66�/�pa.0�;H�@�������pؤlf^�t��	�O��?p�����a��*K4������F�R6Qp]t!5�'���6�`,<�zd��S����#��Ҋ�@N�A%d@'��ix'[���ӽ2����ةl �}�}ܑjPP�us�H�`��ٸr�S�'1�ۍ��@A)چ�f�����$����t���t���|fp�Bi�l���R-�`.��-��2��ս駢D���d٘��}�f�=Ә"��ȦkD4�K]f���u���M�)��ŤX�(�	y�8v@�͝���`b` $���P��V<�q����#�{�U��А��u#7/�/��F�~��4�Xu�b�!G�K�3"���Q��Fg��N��-�7˽�<�1�n��w��{���?犵��=S_�Y�-�@�l҇|B��H/�z�g��cl:�53�LK(�X�%��,%�G�{�k8e�����9評��>b��
a���6�_��-��M&9o�4����rjOj#����>�lr�����뺷�B���F�2�+kI<A��M�k����X�=R��׺	���<J2��dw���_���Z^]��i��+Aʒ_����X@Nsg>�8;R�F��FL9�j��p��v:W� l!��p�:+^4Q��\�C-u�c<?x/y��+__�Al��]@�E�g��9ȟׁ�m�5���3��Tn����N�5�bN���n��g|0�㺣��+����)���f>AR�u�IcB�<_���k����Wbɴt�e/Ģ{-�D���-[z�m��)]ũ=i&�����A�gAg&�+���)P�<3X?�nF�[j.	}#2��S�+����f-�2��	Q�_�ו_䴖5�.s;�JF4����r=��a3:~��wQ���Zg�'n�1C|O�}��"[=��?e�p��ՊlF���� ��d��?}��h�[Wo��vg=E�S��Y������OY;B�i�`�}^�DY����Pu$+u_Z�z�����t�)�6vLeX��%��=;�f/:$d�����<N=�܋��=h3c�9��sY��������6�+��#�-���#�X��F��ƞ��L�r�cΚ@��x��n:kg�v��W���碽��;�b��]p�`��
���{d~Ֆ���bb�Ӕ�[�>�C��8�M��ӡ�v�iW�=� r@_�d�
�g{k3��F3�ȵMyo5�؏YG{6S@����#���v.�ͩ�m6$�5Vu�m粨7[1eT�@�'P�e�v脛b�z�4o�[!3 ���9~�0WԻyk�S)O�~��ݤ�?��}uď�n��IV��s�+�֍���F|*�A�uД��k 3�.�� ��\y���6�h�p���*֣������P��=��v�u��3�̨�H�����g�%n~���<� ��<�a �%Z]aPl��G��d*�?'cU:��c��ifW�(�� �t���o�`�"䫕�	���I���5*��hPE~�b��h�=�_3�rs[1~�"f�kZ.i��cs�����������;pv�W��j���0M��ތ���g��_�|�������Җ����� �=��0e�:GƬ��������UބraG{��� c^Lx��/�b�,&�򛙴�gm��ak,8�������3E0Q\��r���dR�Vsؔ�b���,n�G�;�?�Q������'��ݯ��[�۟|B��Μ��9�}�&�rF:��Jr�wj�sb�2}S���z��z>�u��ϛ��Ɲز���N��l���Ǐ$&}�~g�xN(�����M`�5J%YsJaem0��R���@AV�,]M�>U��\��W���դNF�D����tW-`f���ԶEh��2�ϕ��g����|�Y=�8��]�蚅�����0���_�fV�uC�4�LbQDq������h�%@��������(i��7vs�1��� pn|ŬÇW9n�ĉct��ݾ�9�54��ln�A�%xE>)��f����Sg9}"\Q���)�ɤ󇪵�#,s:� fg�s4X�ۨ<ϭdc���B�@'�w2�vh�L�HS�ywq˛V,�*��^;l� Ѽ'�u���to��Ԭ��B��������\�4��!K��
���>�4��K�6�཈�wt�a��5Ѝ�%B-f��e��G��-*@����L��	���G�Q��j]��H���o��}�]���? ț1OL��t�.��g��c�u�b�=$�Q�;2���'<�F�G�w݆�Q�a�z����i�'������?��|Jչ:]ϟ�yJop�k��{Q�?'��U�CAbG��k��T����6J��Q�m��g��CL� _�Ӿ�!C}U&=���ՆuPm��xy���@��4z�n��d�n7.���Y�[0�4� ���F��&��od�N��!k�է�^a�(�A�?e	�\�&��L�K�a�X	�V��q�u���g�@8���C�	��= r��)P�o��W�E�,�[���=	m�x"Ĭ�CjŎ; �@�/�2g�AaQ����$Pz��q.����Ak̜ s�P��������٠�(��r����-��8�,������|C]Bޭ[� �V�"/�;G'�c��?��.ݿ{�]3X+\�Or黕C%{��M<_9\�j!cy�L�����&�Eu��kc�&�K�i���ϙ-����-e����p
�i:X�>d�x���i�]��jA��ej��~����xc�=L`�6X�����u����[/���b>���&���y���<A���Ag�̂�LSdN�vc��ݢ��n��y�������{ ���Ӿ���pdP�n	O� �����+�L-P�-X�1����co߳����8Q0s0�VMH�-�2������V}��.6:�ׇ��v-O�a�/b�w�L�-����/��Gh���k�bZ�SX�Ib�ޥ�uZ]17�
v؇v >�0����<㇛�th�0k������Bݤ��x&�3v�>Q�ܑQfgg�U%�i\E0� �e  D�#�ӊ��b 
b`a���<�f���)7�i���K�����h�!?��jK��Z�ժ�'�ǚ��"xuP���N1�\��s_��S�*��i~67��3��"G8 ���n����;I��B*y�eM���V �0!��#��!ӷl����vb� ����˓�N�����y�����1fk@�8h
J�Ú�38p��mC�M���h��|~�V���dC6�Jp�����F���( /�`E�w�e�%�g�~[I� ��i�SOq��<ɖ�`���W9�U.`b��O�C䘣!��P�W���5-��J�}}v�FW$m��1��&шU�[]�s�.�����9;��J1ݾu���@!�O%C��A�D:�ɭ�P�W��z�o�� y��+G�۠]�VP�Im:_|�l�3ߕ����=��DSWE_����=�����T��;���^���3�?�M	����G�ۢ�6ח��/��(�j�T2ؘԀ��s�s��D�u��w��E���"f>�e9�d��ĥ+������7��S��:<��f�>����'Ο��.���t�^Z���N��u~�h ��(�r֚w7؂5ې�����1�MM/ 7zB^+姂r�1
��H@�f�V
�@+�񍲢[3���jm[�L�߶0 �z�h����*Y`Y���ZF��ips'��|)���i�cttڢل�,��N�I��� ��9c-o��-�{2T 灇�[�<�6 AF��[��GQ5�V�P2�k��\�j����d�/�o�Ļ��3��Ii*߭Fr�/���t�� E�nd��K�[���c��gy���r>.$���7�����̋J��m#�Vt�#���(���m�Yx/�e&\XB�Ƴ�l0ۈ�ذ�d��A(�[���7\�^�M&��n<d���x�_hY��F�EJ��i�}����>.]�D�t��I�����Gp>�cos�����! cw��Y���ls9�������bKf��<�LJw*VMS�zrԍU-,��7���!v�l(��tM�,��e�gv%���y��dOўG� ���m�e�P�p�ޱ+�-D����j�]%=�\��;��Mu�}�<qw��hv	����Q�� xc�Q�D�\)��f«�$?�̢13�`>G͓�$��;:PUl�Q�1���a�Ź�V)g����%z���g�caZݎ��<�{�~A���6SaH�'�
6��x���_�ݞU�%�pNWP(��=���D�l�k3"����"�փ5%�=���ڂ����S�h�����>��U�ot��w���22]ſ��z���5��L!�'����=��#����8��1�����Z��-v?�ܴ@>;F��l��#c��8�р����U��p �Y�����3]( �}���C����Zs��Ȧ�'ߣ�4M:�A���	Ų��S;������W(�"��D�y�a_�
|�h��h�ෘk5��u@���mkj���g�И٤�v���{O��;����t�(em����+H�S2�o�c�MH9��.v��o�o���?�͍M���l���vk�KT�iy�3�J�)"[),�fx���ʒ	�����Y��rR`��{��I��+^A�,�4�r[���I����,	�.�1��3�����G��GfR�e�{�����ޡ?���1<��D�pek��\I�e.7����G���p�޽4��G�CoJ8�.������яńg��4mvL\v^66?���j�y�BFX��b3TE��#H�6č�t��t���!��eP!L[�I>�sS���1R�Sx��������4�
���,��D���[�(^k�'N^�
n���9������>�S�?���T���/��Ya ����N,jw/s�=�W�t���Gx�;$X�����#�A�����P��s��ܘ�n��Zy1�����hw<�6���T@aǐ�s�����}>�e)�k��[fߢݕ�G�7�?!ϲ1�n����%KF�9�=SĲ�H��2	�b@!2eS���H�ֺ���02��J�-?�콐/Cǡ������M4WCf��g��Y�H�+eF۸2�|�/uw�8���wT�b5T�"9a�{�Dn~��jU�\Ѣ�|��nd���:Љ�k�6��N��L|�ҟ�_Vi�u�gQ��h��j1ĘWk��d��Bw��5���^h�hi+vƾ�F��Y�A]�y�"οo�ޣ��(��7���t�Q��2��A+�i#��UbyB��Ƨ�"�)�^� K9�bWl���d��J@WT-䴙i?Օ�e��y�)���*!���xq��99�^�-R�n��&��oQ�p2��P��Y��CS�N"��r *��{ s+-���:/���H�Y�v��1� ����j����э��]�$`�B�`�y�+g�+Y�@�s�=�E1���f�i-��=�ɫL �Wal���1���Ȅ�J}�J=``���
�I^DT���ED,&I �X-�c��ASm֠��𨌍�魆�"�n����4E���y.<��G��{��0��X�CBfmG�����U�?ǘG�Q*�J�[ǹ]F�+���6��tr*P��=͌�`��4�ԽM��m_���i�M ��y�}Ώ��%r�O���@d��g��-%sM���ϙ��ʊ�s�V�fߗ�Xdpk<4�j������?��[W��!@2�ʧԲ���~���`��Ӟ����{\�2�M�N�vt�87�[(�샾>���=�\#�B@���w�Y(3+�)r%5��ݱVd�}��!v�`�x��<�S���T��� X:.̥�D��p�k����1z�fi�ֿƤ�Lﬠ帾����ߚ�>�]c0��ݶ�ֻPY�q.�'dK��g�>W�2�ls�{G�Jpe9���:��ި�x�,����L��Y@~��׽r�
�\�B9]ze}0Fm����t�|Gą��z����myi�iL�CM�����F���Vr��B�2,h:5k�i�=}�F^':f�7�+Oj�ki��p2���m;|�d{H@��ɗ8��@ESz��ߌ=,߱���H%x�J�V�z�L��um�پ�{�g-�"����������fDN"�͐u�]W�Dc�=w��������,(ŤoNj�1����_��� ��w�Ć��Ex��ud���oe�ԕ�%�486�����ݬm�/=�� �������|�|r��u��=����(V ��Gw��HV�|�7��'�f�$A*��B����t�A^���n�lc�Q�<�]Z�7��[�f���#���X�ZwQ�C, R�L�=zL�)���+�8�Y:�]���N�+���wW���&XBu�{�c��vY�{��;0
�h�F�H@m5�d N�r0kW�H��� !��;׬h*0;�ٽ�Z��(��л��{�7����yP����rkӥ��1��LȶV0�wr�kE������{��hCm2Xe��>u�@��Up��IB�)}�*4^/ @��춭	s-��B(��`M�Vi�u��}r�B��B{J��<�^��'.��fl�׫�l�^Dv�.ͼ��Vrmlk��,F��].ȡ�ؖs�����j9���^]M�3�9�)�jT(*�[��!7,�>͕d�0�i�dA��� gF���\L����
 ǘ#���B�[,�)�Lq|=���
u�m~M3sѬ�g�HX0d!��M���~������_3��p�~� ��#�U�S�F4砀q�O���J���3��=�g)�q�� ��A��ʮ	�JM��F�ӊ�ȷ̅EX���?�4`�m$    IEND�B`�PK   ���X�䓶� � /   images/132fbcdf-34e4-44dc-827d-09a965026955.png�wT�Y�/��QgPA�H�%PP�tA@zE�&]���E��@�H��~����ݵ~޻�]�����9g����}�9񉸡�u�����赫 G�#'/:�f`�(���5�C�:t�1����z���k �w������)?3?COG?�m�u�p����� ���JS:�@�E\��/�{i SB����[�?���s�?���s�?���s�?�����
c����A��?���s�?���s�?���s�?���s�?1..l������c����DQ�;1����9[%����-���w}��.'��3;�\�/|���Wh��ж�w���t�i�%��_��������~�j��w����P��S��OZB�v�3r�r��E�8:`7�h֤���`b�\�o��{"?���s�?���s���Fq�� t�t�k��iWg%��ZQ���X���9�G���N�Z����谥#�鏀7z7�;��]n[�PQ蚭0B⏣��/���t��/wetiD\B2�Z�QF�:�+auY��f\�@�;j����+������'F��~ӣ�+�qͪɱ����E$��@k�]�R���.#}��J׽��L:�Ʌ�?/ZE(W�A�*�>��,�gT��.���V��`/�Y6�l���g��G4��乄��6K�E�k5�	/��u��]TfTz�MDڝ�==����D��T��y���
��=���]��|�	e�i�f���k�N�O2"����2hە�,^�S�Y@�&���2zf��K���y�ۻm�ʵ ���sm���Ȅ�WT�J�=~�	Jqi���.��g���r�u�&����&�+
2"��u�����}�۫����<g��:��sB��?����
�m݁k֢�97�����F����KؑQZ��v��6?QTj�M��	thf*k��}H���C��ߦ������^0����hKR��AKC{�{|]9��3j{4��������Ur�t[Uǣsml��o߿l<���"Vi<H���xb�lr>%G'�+�`]�h�O��6�rq�3
�gbxN�\��il� 8�Kb�iՎez�����N�]{�Ҕ�-I��m-�dTy<,5PF�ɹ�hX�o���md�^���s{ç��~��~�,|��; a�i�7#��ċ�SB��:�.b�vUrs��Um�c�ٹn��I4/"�Y���l��0��&�U�ptY�MY9����T����v{�ڞ�}O|�H']�qA?�.#)~�J�.}�n���F�H��H����S�u�O�}�)u��Ӫ8a��{��%����;����m��k��SK���ɺ�sYw0�������,DsUz�l%�
��ʒ��q�G�1釠��``��m}��Zz����k)%i�򣰺��;�M�u�*�/W����z���I%1ԭ`�@��y��䪧�7�SmƮ�u����u[���\��G�Ud�ב�ڞxݎ�4l��M屵����{�w�h,�b���Zzc؝]��	�#����Q:)��	��^d��Gv7�����I!�q
��>������ƞ� ��`0�Z�-��%���F��ڒd=�,Rm��WvG�A
M?W����O��/�;����-U� �����x����ǲ�^ 7%b)޷R{:r]<��N_ ^�}a���� ����Xw��>Մ׌��2I΁/]X1"g�2���@΀�jU�ۄK�"�l��Urn4�&(�&���/V�����K�[�����7��>��D���B븹C&�/�٦(ԢO1jk����P7��Z���봵IN�����v�:I������mEZ5�=�3�b2�߃��g��p�����Hp?M:��9����v��;b��Qw�Rz�D�,c�J����wF5�z�sʪFW�}�ޢ2z���`�̬�J4Z�(�2�r<.�&��K \R���>u����is��U���O��J� ���Jޱ������!<o�KVI��\�9���/�1UF{Z���=-1"�)�H���h�P�F(�ȥ�L	lB�i�d�bՑЂ)��1����#��~r�����5s�/L*�$�}YI��l̵Q߀I�o�4�2>��IXjھ���x����p4��᲼���$$��7���i���s��\h�o���ڤDBC�ս�d�u��u"Q��4(�_#�U�4���˺��2O�s�A��V���ᗛ݇#d��+l3���pC��̮sc2TE68�Iq�BD_@e�Y��I����-�@�H/��
s��7�~1]��s%��d23�)ol�v�֏��)"f�l�o��3��������jD��Q~C�i#��#�Z�4���������F0�G�1cط��6����VeX�;��>��>fy��Z�v���|¹���7�d����#�
��d=�2��~ߵ�Ξ��L�U��5���O�����ۇ+���#v-�TM�/L�&�V��ѥ�޷tB���[�mh�9��V���D����\��|D��v�X'~�1�πY ���)����� ]q?�Ӕ�����<�6)�xz������Z��UlQHG�y�j���� �G �IH�/�
��5�@��b"M/y����7M���a}<g�VY=7_7�`���&�b>`��e�P~�Cy�lm.]}��K]�}6Pt�V��"#筬vr�;�\���T�UȜ�� ��C;H���T���r઴fQ�js��&�V��y�e�-�G�`d�H�l��8
N-ib�����pK���S�Sݳ<y��mo�u�� �LN����2m�d��4�WR�w�<�azcc+���gz���u������V�e����.9xy��u��A-�&?U�U��j{(r�D^Nx���f�7�$���u�LȠ.�~㘱���ҽ<�Cg���'B�^Zz�;�=���S���E�U�A�O��*�Jn��<��a�?�ܐ? 㿯�V0��kq=:Sr95���h��-nԘ>^6����:�J���4G�����%�u<���
Y'�=޳F�u:�z���%���U)[�/�{�*���V|��>�4�e3Rrx�K������j1| TDH��dx�+XfP*3M�,X (�`+�2$ X�f+��pE�zf �������Z 6�xx)������A|�[JUN]�.?ʯ�3�>쏣ו<�p�v?;�c�dI��U�Cbg�L�����1�Q��3;��]�+�_�],`�;ژ�Ņ)pu"�E{P���j���5~4��GѿC�A=:r�q�t7dwz���{�E�ȸ����<��_-�Лo��׏%�4��8mD���>��{%�ш$Id�[�eYk0�m猧d;�t;B*��>[y�-��rD��[�ab:˟�ܨ��|�x#pu7������}��m��=�5�Y�
���|f��5<�YL�L��TbA������u���E�I�U�A�9��w�SlM�3wI�����L��������S��qU�ɞ��ۛ�x�L0O��T����}j#)ֽ�`�:N�ҵ(��\5��Y��um�=�"�I��J�|ro.{�"4�
rI}�����ux�Ln���[�q��g���/�u��\I��ғVY�Q���K�!w�2�yre\X��'���B�*d����"����ȼ�*!F�AΨ�8�B��鹻z�G�M;萉_���!��OL�������}��3���)0�Γ+gA<5����%�X=b��C��`��лk��=���[c��{��އ�X����f\O����~�Q�����0aru�*�f� N$�\.[zh�p�5��˫�E�Q��
�t�Ū�p�o���s�q�~��5N]{�Ŋx���b�ߢ�y��<��dԣ�j�_�G�������a�R�}�$c���5gD����������#;{�;���a�R\�o蕱��9����)�BBҏ$+���D�1�!�ĝ�8��T�1��|�Y+x3
��65���o@<\��,�0U�a�kJȔ��?�u���XTG�N��{m��
0ZH����U�6�Y�պ���&����b�&��\����y�y5����e"N2gK� k��0�xPҩ�/��]k�WYn�]��@m�E�^]ꍪ�~�Y�frF鄩�p��0&�;��{��ڸ����W8���6�R���bb�:�P�#6U��ms$A(N�o�6(nU���[{��&�<{�pV�3��W��$A�:' �0G�L��Ě� ����<��U;�6����z�d1N�8������A�ʃr�;1��s��E$|rMu�7W�y��P=������O�X��q�Kυ�'-��#�{�x�$��c���=M�b��MP�Flv����������ݬ����`]���'�Ω�s�V+D�5T�v���^��f����j%m����f�� �A�|>Ӿ��L���d��L��v" ���r��,_�f�Z��?O|��j���]z�����<�������w�!������n#�05��lo���6Q�^ǿ\xsP��^�I�4��xc�UG�A3�O�dݹj%�/���`�������(����ҕE��v�}��*��s�m��`���wz�/'^�N�!�p65G�˝��Fj_��s�E��w��ǫ���Q`�*e�r�>L@��VE�A�θS.��&��P �]���LT�e�Y8��O�)�I������8[}��,�Q6�.���.t��.&e}//�l��"��]5�	ZSIE"F�����D̨r�N̎/2��I%�"4��+]���c�Sv|�(0�ۏ5�U�M�ߦ�x��q��4��C�,��uEQ�x�&�¿�$V�&ۖ(�0Q��)U^��Fa��4�Tgu+���sC��ͳČ$5�Y`dY�|���U.{���X0�1�1�>�2�/zi��xl�I�M��G��Mh �_�\VG�,�D3ކx���ƣ�0����ZI?�'��J������F��Ѷ������իn��A]�E�4��j go�\�H:93yBBT�7��Zn��Pha#1�>���L�j(�*x��ڌ'��+TEQҹ��Uв����{-��0���g�m�O@̖,T���mE,=5�C6�(b ĉ�E��
��L��T�R?��M��V�|3��I��M\�UПZ�iTF�1��1�1^�'h�CZGl{e�,�1��,���^�d8 �u�A�$����N�G�αCl�ɮ��Sv?����˙�g�A�NX4�]���o�!��쌢�wYA������&��V~�܍�Q��`JϏ�nG���=#�lf�ٴ¶c�`w�X��� ��x�ӥ�<A�KOC��x�@,��#�s�vO��!�c�(V���r>����}� \U�;��d������j˾x�^:nv�xN���i�Gb�n�p&=2�}�(.�!7�����[ ���W%��!��zr��D��!��lm��Z�rr<Q�?��B����#���o��+�[�nA�}!�7@��b�>~�/mR��쵫������s�y���_�`-8à>��q�V����q���2����g�r�n>|��f����Ĺ!�BB�cm�	3r��kiǞ�\$��e���/�.*�1`TغJ}u|�Qa@�y?�̛��Y���� 2�F��|O�"�C��BRa�׾6X�aF9�oV��B������Ч��	��4��<T���W.��Z"D��\y�������ƍ߇�i��#Jz;�!4���h�}��E9��I"��
G}x����<�E��g,�0���A��
��.�SE������
�A�l�}�6g��ةS�uk��>�ghi�=+������>��k��c��|�Y��1#n��8��&�N�<<Oj�CC+9�+K�WXᜱ���R���>A}�B�<k^�W�qW�4$���'P��B�a7�q·[�A2<�����VSѐ��z�B[�V2{sȢ���|�n!���p��)/&���ΑU�W���w�6��_u�E��]�\���O	����)�-���I�B�y�́_sԮF��)5_���9��ܢV��sͼ2��˖�U��U�>��dX?9S�����F *���'��:
lg!;눻����G�B�������W���쾿���H�sV�A�/�o�Q���MI�=����J!�tWl�U������F��&�y�A�NB:��%�Tf�#��5�-"�����^��_��z���@����!l�F�'�(�X�K�1*��ދ��dN=z�p}�$wE��G�n��+��- ��0	�=��2j�Z,*�-z`�	ic�hzf��R�����om��^�����Q��=��8F��$bxE5+H�#*i��1���7o,��޴��s�6��]�ƻ�Wn铲���U;� �e@��-�͌u���(���ֱK��v�LV,rQ�rGE�$[	��<�7�k����N�ċ�myxn�.r��/b�6
rm��h�{I��'����|���W��%��}N)X��o��P�z��X-�:�1}���{�����A�iH�	��km�{���t�M�^A�D��A
��QNb�DO��Q<2������~I�����g�7��P_�N���E��x>���@i1��~:J�BU>��K�\.�(�"��ē|e�^c���@�� dS������4�3�{�'�<k��=/�>$Z�AQ�-������GĨ����P(������=�$���9V�qp�,�y���o~�]�)=����	 �ziC���u�7����J�~�JUE\M�T��Dq*j�^ �~�N��T�5�L���O��1+K|[�x�s:�Dm�My;�W�����~;��	�zO�Ჺ����!�2�bc(Fq]�<b���v��*!#_�ַ�҈%��]P> �E3h�MT�
^8��ӳ�~�6g'�#\��\g#�7������v1��������\�<SG�_[ۏvx��J���d7���_� 4lご4��.$��l��Wn���OhŜ��[V���a��gM
t2���%S�ĬF�A� ��Bo�|�[�{GN��߾i�~��2�I��_�"Q�N��}���^&uf@�W����� d�"�i�,���z��ؙ9N톀,�`�mF������I����o��l�4Tx��W1�M���?Cn��W�7����;z���T�glŜtH�ߝ��'C�!��?TP��C���������"
)<۶�1���4����y�^�v�yw~�t�ze�f�5�{!�Aslgc-�Ge���@)�ϡ-��z��*��8R�����Q9��[�Q������L�K��W�%u��}18��v@ա�hg��}{{�GyF�Q�Ql���7pc>��Z?Z���������(�\�|��$���5������wh�G6pg1P��8�c�?'�u[=�J9{��L	��I�-���ݭ��?rk{��܃nھ�X����@P�p#���޳SB�&�ˤU8�ؒ�?`=���Z�$�8F�|�=�⋠���	-Y����у�^���}$�u�ۊyj��yx-�`�Q���Lp�Q\*��@��aЄ��t?���jp��DNj$�LqV3,9�R���O݆��;3q�(��5������n�x�b:�!$�a���26����(J總,�=
�0'�ϋ���!+�TRPPWJ/�>��T�L��m�~@���jnI�݅{�4&D��
��ܔ��4�������$À�"}��q(� TAG��4��K˪���p���A,�o�\j���|�D/?�3���y��@>`��L�9�K+��W��Դ虬87�ڑI3�a����$}��
E�,�
o۷xŊ}�@F�X$@E.\��rf���R*�1���x���>���\�L�����RSM�Q���yOX����C]DlvL�M�s;���cW�p(�ݞ>,Bw�^�?=��+��%d��}ˠW�Z��k��Qx�3� ��o$U\]���u��l'/�D����VP*q�`�k�Z�ݓ��V���i�D��C�N,GJ����)����4��Z�ɏ.\�2H�j��I�.�S��h��5��M����ʃ�A�)s���읔��_��q�uC��q�8w���.xm[)pm�bpm�I]�~=w0jZ�t��e���`���A��A��~T�>��j
$�mYМ4#p�?�#rg��'��Yh�;Hj�eWd��w���W
6�{Rs�[�`?�AMy�#:6�lyB��� q�ի��}_��6�=܉���j+)��� �L坏����j�)ۼ���3;��Y��I��7$o��������ZicD �l���ksv���VjP��l��&F���pd�&AM��m���-MG��*�̏��B��N�v��F�9�M�C�	�#�~2�����CsH��Q>3b�PڎSna*LY���;ڮۂ���H���"��O���#���/��K�Y���*��P�W>���k��m}iCkH0\r���	w�:��ua�3`��k�w1�`�~�M�U���ـ�}�!��;�`9����Pw^�X7�[�LU׶���v�cKѽ�a����!tf�NYL#Yv�	Du��#�y����̭�_mF�`���
����ka�ƥ�W��	��dj���T���ؤ\�[��\�W��]Q��תv���ci�wh�!�@Y�d�B��LU���5Ņq��Pw�Z�ж��^���a.�*%� �Z���rߑ�n�����_l�?��x�x������o��b��u4{Z���v�����αQ�T����WN��W�&���ɛ��I^۷Ѽ�Z������OT@]$��[��0��K5�@a���ۂ[ƀ�v�0K�F�Ԙ��Ǜ���˗�H��Ru��s��DH��/�DR���9�F��jS�A�&Md�f{U��f�M�B@;B���؄܌<5�/���:�+Bѳ�B͙�zaB(&Bf�F�#gԅO4��Ze�]{�n�eM9N�ʁ=U=�uKc@,#>�n�l�H:����f�Ǩq	4m��>�g���=��K�yG�^�~eM���1��Y�w����^��7x��V�&�����'#�8��=������rSQTQ�6hs�eʓ�\m�����gi�=֜~Ec_c+^!C�݄��?S1�""1����U��l"� ��/ w��6��Kk��1\.�����%� ��#�j�#72�C|'��l�����M�-w"������7�0�����h�#���>_cc�7+�����T<��0կp���l��^�6ȼ�:�r��|�m��x)����{U�;ӗÌ�Ƃ��vJ$��ڟFo"�¹�n��H�[��`��S�@;��$M���Y�V3�cY^�|�X2�w��wْ��;�p;F��jo}M,2x��FuǺ�w�@�=<��Su|j2��R�M_A����Y����$e�%�/9v�6\<9���8��@�m�tY��2̺� xmGvGi�L�J$W�[�����6���&���Q��Anv}�S�pb�8m{`rO��\:�N$�nT?����w�i	�n7�O1��"�;h;�΅~5�>jj�[įJ�(��J��e�/��}ȓ��=nAC����).�wd�V���,�\ś�������4D�p�vB��аo?̟k ~1M�&
65c��C\@��K�.�R�郹�,1�H�r`F��J�,�O�����G���U3wgiB�L�v�D��\"P/�6��%�f7Sm��+Ӝ)��|�g&��qKި"L�?��4���u��r�>T�lu�b�У��=���WoS���M_�F/��KH���җ�6$���(`��a%#$�Sc��[;t���9�~E\1q�b��'�0����@�e��|c#�i�+�]k}����j��s�h�W��&�@�v9|��J�֜��P�gZ���V1[�٬#'}�G���R��}��ؘ~5�mȚcJC�<����9������b�~~-*������2�5���K�*c�X�=Z�R��س���3�����^�Q��"J�o��sV�V�b�����dB�e��_��ձ��,P�ٝ�T����w�����kaJbm�ѱA]i���hK��ظI~y��G��&0$�!ɤ�X���9��d|@�Mu�3��0��%�@�Ѐ���X��a�	�&����N�we��M8k��~�<
�PYj;������?��t�ϱ(!�}�H�4 l��{�x���Y`�j�;�=��C�<��wd���&�{�n���POM%6�#��q�>�0#1#4���:��!�X�0U|+�Lo���A��3���Σ"��3=�t�z� _ꔭ�\�;���L��k�3{��d%��,����@p�U��}k����w� ��o.!��8��ɦw`Zh��wؗ���W:���}�^����z�?���@��MŁ�I^2���P<^�IcB9��������w�"_�S!'S�8�7�����P��
�EO��\��xbuݰ+��qߚ��;�<聲[�w�VS���{��� �N�f�@Ƨ��Eu��qb��T-ǴD�݁�$1����T3c��!�V_�:t���4�c؟�9`��ÖlObN=/�5g�>�U�6�Č�Ȼ[R�^f�� �.���0�{�=�(A��Q��k}{XkN1��X��`��NU��h��0Y�f���]=��y��5GoM������x�
.�t��F�v��.�F���� �e)z@��\�&��ʼ�}'7-qv�)������*�u(;չ*7gh�AM.E�!-��Q}Zި���e޳;�Y,�۴ẽ�֋����|�}{N"J�7��-u��T��iO����q�u�96c��{�|��
�N�AHk��m�^�T�X�'���x�����0�"�M�a=���Wvk����'�q�k����Q�:�C��.���nh��zu~��z�z��h: �-[C��6��N�ǻ��a�`�l�_Ā�q�:���2�i�F�Y�K:�Z��S�4�6�_E����&W�k]��z��I���g��׭��[�`�=T
l;�g���֓5���ꤍ��r����n���4vٛʦ&��*4c���q[:K��/�G滑8�7�M��=���'�m7�K�A&o�Lu�I�S�o�4���&���(�J�r6���W��o�?v��@��iWY���$�Wty^���eo�/U ���@����Q�ٞpG�{�/&&���=[4G��\p*�p��1l�A�A_��2y�3�/շ����r�޳���������l��.�\�V@/��	����?�/���_�R�#�����'s��]�x��[? M�[U,�'�3�u3��&c�ga׹�j� ?�+y;G��_oR xg+����՞	���Cg.*�󒇛�,�i�1Vr!P��Js�>��^]ҫ�؟�ZC�[:�z]>�R�,�<t?�K�`��Q�^r�]��]N�N\���&%v8&���I:5��aw��Ƽ����fڑ��N�q����=��zN�|C��g��c��?ί���@��s8��~_x�n����kJFy��Z�3^��6@��S��U@��_l�%���.�l�m�-�=�l�	8#9g�lX�۱9���D�9S*�:LDx��2&��c\
 ы���35b-��`�iA��l��F�Y�:��}P�ܧw�G���ge����y���0\��7\EG��e�*�CP�罟��N�<��z�k�uOLӝg�a�P	�+��;�r�xE{�}�F>�xQ����$C��%?��l�g�Li��X���)w♴`�ܩT��/F�)�@�<�����ש y��w����ea�a~����
(����Nb*���v)\�~E/	H�ŭz��?�Ԡ���^��}���������^D&7_���>z�-�� ol��8Oy����}-�[�djGY�� �9�M�'�-�~_��Ě^�U�z�}�o����9I�ᾈ&T=
���/7��*��"n�!]-Y���/$v��
ޯ����i�f�ݐr�^��!t��<��T���2�j^oQ_����u��߮]}'$�w}���j�\�@+n�7��$�VM��'2�!~@6R1��Ȍ�r��b=���f��J��ә#�$�K�-4ݒ(ޗ�}l��؇4�o@Y����߷ �����A �Q2�>��#e�[G~O���<R��!��n��*�케�$p���W_�2��zƌb躪Dj�1������]Z��G�J�eX8͕��U�Ž���M�a�ཡ� �p"�i�^Rm<!�T�S^^%g>qs6(�U�K�8�ӡ
A�~���^�p���o�I+�A�
D����8?EDM�d�"Ԗ&�V�Ӯ�I��a}����-L �M�������f$qx����):��"Fف��j����o�7���K����#EOJz�sC1����q�P]|�$�l-�bB�����#�gX�%d{X���m,��~cw#(^)謱�nMl>�@���yT�S�H"\�ˏz�S�VÇ��KaX�*�t��`䮘_B���>�X�Ȕ�ں�~0��t>.�
mj�6͎+��B� 6��n���bf	�Wkj��L��pZ���&�[�u���*���p�m3m:�-���q�D.�d6�;]W}'}�ϥ�Q�)E�۬X�j�>^�G��G˘�p�@�+�ڬ���(����ΰ8:O�J���ĖL�y�JC��N�!�T��xQ���u���[l�A��O�C�%j�<�=����B(�R��l7�
���`�uf���\ bH8L��������I�r-Mȉ�*RPw���]��:��~\\t���/�^��zD��ފ�e��0��-*����۟>����9z/^��!~N��i�E6�����'�S�U��=�z���{|�p%����U�OMvU@	[���!�$���Q��]�[�{��biU������+�`�)���k�v�7��u_ؽk>Q��~�%_*yl|��a�ca����TG�577}�����-h��k�+���Q�jq?VY5ഝ����3`+�d*,y���,�[y��nN<��J]D��)�U_���� �~`�NU&�s՚�F@�z���������qS�� o�e��yJ[�*Jo��5fgO=��H*"CwR���� =^L�c����	6�Lxu� ��|��R1�b��'B<k���M��&����)����	�	"PO��~ rPγ�nO%h���VI�okq@E�g�ԟ��U`��*���L�xp��
�"i���HiA�a�Z"�ئ�ę���O�cZ��cgp��h��Ls��LT�R�2��vnI_���ǈ�܏{�� O�ߨ���\����o�ꘝ>���.��8��Rw8sJ��kj.u�5�*/��\_a˂_�=�?o��$�YC���w��lC�B��R{8�[�\�K���E�*�w���7 /��U3ơ&����0x]3�e�,C*۵ek�B��X&Ǻ/2��c���![Ҙ�3@-+zاK�-�_�#�~��
�/�i��73������gp\ԙ#��:��yb����(,�
j�L���y����%�@	��@��ˎ���2��}��.���?�j�j�˸
�8.�ߙ�ژT�/�ߘ�<P�������ŻN��	�-A�t�}�<��i>��tP�L���Y�ʾ~�2.�7�{��
�E0�V=��=Ӫ���/#�b�t�K3�1���N��?`@����z�D���$Ѱc���� ������c=�Ы����׏<������<��Z���c�;�2��!���� �u�Z#�ef5/W�`�m�'M�;�#bU���2��p��ѥD#�`/w�����~�ꈘ�>K=O�ݷ&m<�j���u��n~�����\�zt mp|���`"����1}�D�+2�/�Z��l_X=%^l�Lv]�&�}Ï*\aFj��ǎx&m��0�@�Y�Ws������&A�>�1�Ui/qs��Wb��UQ�s9-����}��Qf@�:��B����lA���2��͌�y��m�5;�z�޷�.��������ahm�y?#W������!�3�����T	�q�ά����i�Lu�|�h�3�c���U���M�?O��̔	{
}C�zu�s��ۂ����Mm!}(
�������uD?����\�����s�˙��{�,���:�XШ�}g��@APVN0�����մ�E�����<��R��GV

R�V~l�ϱ?�^���O)����l�<��:�����uKĵ�'��`�$��dr)�.��FID]�zP���LНC��/�\���"(gv�ٮ�f�o�S��A�:]V��;TrkZ�~��A�@mq�@���i������m�Ⱦ��yfMN�{S�U�Zd����V�%��`^���Z�Ic'w�����<,��^L���9Lb��쎑����(&�U@��e�io�!]n�ȱ6�(Gw��X�!b�)ڦ�xTTۨB����K��l\�/Z�o�q�nW� �l������&�,>����2��U�(�M)���?��{��xY>Gt?�̠%x*<����,�(J�R��+��oL���+Ø��c��wo�|,p(3Y��y3S¹d캣�=+��1����D�_��+�W��� 	����8��$bhF�v���aoj�_���y�I��ҕQ�X?f����;� ��R׶��������'�4�	o��6Kܻ�q�\���_��	a�k��6
��a�ʳ
��v��!��k7XD�2�y��P�İ.}4H�\�&��ˏQ�(֔89U�~-sM����M�`�x���Eu�L c{l��Qg�)�v��?!<'�)���*R�q�� �dwIp~�Pn���X�%�8�e�-�4�4�����&-��h�1�]�� ��t�3�ke�=�.���ϗ�k����m���@M��H�m/1��T!���>��Ie����3����u.Ļ�n-f3�J�:�ʼ7��0���1�8��g��.�h���Ȃ1(��J�ŧ�c��PA�Qǲe'���IƶZ���j�52� A�������xO��L�[� TPM�6����.�Q�e�}��v<�S��
^?vN���������8H$�L+}kbJ�Bf7cX�B�\l�J�3�����ȷ��M�ۯ��T�~P��T�1Y� �zo:V�8���v�~p Cf�;�>Р׏���$���p���jJ�5����I/P�{v,���^??Z�*u� �2բ�j��.�"3F��<s��F�<%���<z
k�8@gnX���XF�X�*�!sZ�퉙0WO�@��_�-�[2O�[�^��=r�+�m5݉y�>�<[�NGm��Z���VOn�+�$�G҅ 4R�VD|Ջ��o��ʄ�H�!�}���x2
$�O]���b�t%��׻�����!S���yB;8��OGϘ�p�Z�97t�h�ŵ>���!�2,����_�i�B.��틳/=Z�(d?�H6f�&�9Z��vo[�hL;2j0���Sb�vS�N�FG��X&��v�C������ e�R���'`�BE�;L��x�7�	r���~A�������F���MJz�Ci���(�'�,�=y��SW�0l����ۓ�RLY|u	�8�Yh���nf[�X�ڦ��
1�
��sUd:����E	��<���<Q1E'eM����h���}O�;)X@\1p�4j���AQ(� �YG��91�z�����Ў�H��7됆�H�:4x�> �ɱ�ڄ<C�տ EP�)� K�s󔸩VZ�[�)�#r���T�pӟw͝�P��Q*�W�
�#��o�����b��]jo!�̬��
��w�)k�G*r$�2��J��ǏQ�`s��!�?����������r�A����;�UA���<ٞq�A�x#��V�n��r�<�͖�mWF�
�L3n&j����
��
���R%���:Ef��J��ÿ�5�O�ɂ�]�q�@qZ^�:FIFW?��u��ILvC��M�߽V��;�#<W����I�N�"�z���})L�d�∃���s`��9�E�X]�C ����ՄDk�T����z���~<����J��Ob
-z�9�K���>S�ٟW!����a�6�<p���P�Ds6.)@Ԧ�٪�p4r�3 /�u�$��ؽGf�t�>�ws)�x�L�fy�A����wF�oѸm���N�F��ɇr�AL̎e�(oW���$��hpB���p��<�H{�ѿ4`�}����.x�?���-�Kѫ�/�m��v݁�?�5�4��Xގ��&L)5zW�`ypD��5*���L��su����BP��R�<x"L �x'��t��t�ٟ��(c:^��l�3[�}��;��uz+���4�$4��d�<�"�j��m�Y*g�{�9���<�(�����!��+�>��|%��8�Lz�j�P~�����&�:����ڋ��ֈh��̑�@1�C��.�I+����,�M"̰qS� }�Rt��U�����/��X}�̭��]�Y����xө3s���R�s��_ؙ=_s{��ʎ{{�����k�ɷ�)5aW�VQn�@ӥK���/M�X^c�Ŏno�j% �����6h&�=�j��j?�V��*�+/��n]r&O'oT�>δ)��5}Գ��2�NW����o�[q������.ϩ����')����M�e�Dt���_W�<�	���?8u��(0��T�I(���ԙ
�!:u�[M1�ߐ-��L�8J�׌rX����O��ob���P8�W�c��B��Y�>�	���7��@Z�������ax����� 7��\�Ce@%I�+�?p E���H�ItcV��U�/-MD4齾3�G[B�t{^ ,4&��A]�:n����y1\��ÌߗT�2K a#��;��hĘ�H��xU3�NR]̀�]�2�_��6m����M7�忸	��n֔��K�^�UC���@bZ}���9끨��J %�qE� ��gpYm�[A�zq�7�v� lۏ��~{�GE�7-���F|���]�������:�X��	+B��uI�e������뛽Y�.�R;�g�|�<Eu������ e0���NdJ���K�,[t�~��Ij�O��*��;�ܷ���g��F~`��8���6G��3:%�?9�l�g?%����{���'���#��ב�SL�M�__��xkd�YFh�]�9n��}i*L:�Nղ����t;���VJ��\�`ݻ�`�D^G�$k}�5?=c�cn�2$w7n��?r�c쯍��JQ鯩��E���Q/�!��%�1rtS��I����\��EL�K��r���\Q1(q�cH]T�פM�c ��|�nU_�*���Q�1Ǟwԧ]V��.sS.㴳�＆�ɞ�p8+��dE�+ O�ʶu����=a�:�i���4�����^3�5����\݃��w��Źz�����m����h�D3K�D����fy7�?EY1�]Ev�9Z����h]&Bp�H�/�QK�HE{��^�\Q3I(����`��f�C�N��ޝ;Zɲ��Dc޶ڼ��Y*|D��@b�4a�l8uى�6��������T�Σ�����ڠfV�f���@�zMm�z�<hs]��o����b�\d?޸?�C�Ό�.�qJ����ͭ�H& \�]�q�T���?�����&�L�s;t�l�?�����m��
�[���۷6cc�=���fhv4��������z�x���|���)KR�$%�%YO�%	!�d�'Df�t(E���c���5�0ʞe�����n0����>�������C3���}]������z�/
I�2@�◭(ݎ�פQ�۽���*�ȿ���f|-��[�V��Wo�R�3I,�I\��J�8�|�5�Wa�Y+�J��]���[�T� &:YRH���`7��n��H[������h<�n1�u��!��&z�}�����,f�?��V�u��C4���)k���J��d�������.����^{��gǪ��6�=����s��G�Ro�H[�ͪ
p�r^��P���r ' ��[/�#��.ژ�s�uc�B���Ǔl�A�up�:�Ԍ� _�m�q�XU�C�Ҏ�(�}���ϩ�����fV�P�I��a�!BUՙ���@���
!��\ۓ�c�o�ܙ��.9m�=��^�D���c�j����� ��&u�w."�W=���&��d�\�f]����G��Y��0.������F?*��Sk��]�wECx�;>>�Ґ�;"1!ٛ����9�+�VD�k�XgZjA�/t���d$����z����j����O�4@�A\�����8�5�Ur����@�@
2l:�*��(D_���:
�I����������j@ ����Q0���X]��I�E%�ox���3�p��8�۠m@<o�bPq͓Rv��Ǉ�[�#�"HlH M<l<������=r]C�rt�����a�L!ߟk{NU�pΌ6<qq1կ�M��I�N��ay����΀RQʧLX��;����2���\��-w)�?��'U�K�?0Rs���C�~�0P��$Di�+��L�Ҿ�TlU�� ���󠫘�P�	�drI�4E�[_��X ���B�qV��w�h�91�^o��l�fS9���S������*��<@+�7����s����ty�̥�� c��Q������ٲ��^ԥ���"N�0�<��xrU��t�}�����7+9��S���C���:�C�EM�v$�(�ٖe*\�)0��Â�hYYY�c������ID�pY�@��*%�m���jӱ�z���u�!.��k�̏w�y7�u���J:C���#��������z����&���a��i��������wUJ�=��mӍJI�gfc+���h���D���$�ښ���c����0�vPo9/{��[�y?cx��!�������L��b�J����vC��������/�������1K�s�į`�qBE��d���i��s&{[4?'ޅ��!Ấ�ib�@�n�.�r�Z�c�Nr0���~�����m��UNPC-m���-�(��L>�M4Ց�G��,Fuj3���<K���͸C��}"�lc�zI�`���T/����Q������L��⥖�۽�$+9G��0��ǾZ�h16�D.=�jϔ�t��K��Ѯ����L6�3Wl��t#��{V�3��!-D9�������(̄�PAa)�����˯ɥ'W;{�dw�.h
|���ht��-oxK��������50PB0��r��>-�?/7b�]�	�h�Ȣ�c�Hv�G�O�ٗ�6���T���q�O�q~f@%=�fLdA��G�	�7K�U,9��̍�׽ �S����6�z���d����6˝�="gc����yLZ���[�}>��#�/V
n�]_i�����h�p���^ �[�%ĉ�/JsH����	JVɰ�s%�{~
��L���=H3�Eή�a2���X]�҈�O��:�z��M�8�X�����y�6dOv�}�h�K]a���� ����M�/�FR���Q�'pu��J��J��uDD��U$-/ծ�7��1s���;�B g��B������!���_���{6��P�v5^ۉ�Px�K,K�8���ؕ�����.�yn'��T��H���_�C���Z����*X�WH(s{�^�֛�֩���̊R��24��<����}�����E�c���;]2������j���p5yX��y��|G���j�0�(W��e)�SF� �tKj���h��7 ��*m�%�C$L?Eo����\RX��g� 6]05卝���5�߷΃�<=��󥫫��(��RW�;��J��B?4��1���K��L��I��!��cL��ǌv�7:d��ʨڛIo���^"�=��)!��{�5@O�p%ۚ����]��T�XI݋ʀ��/WG��IV�+t���[�: �<��F��5ݩ�v�?x�ִ���[cϔL�N1>�E�����x��|� ����S��ҷ�S(��eHQԪ]n��?g�����_$��ٗ�J���|�z�#W,#7��i�O����7&sY�)���ߴ��2o��kl�
�^��b��mպq�Q�S��]�:���/їL�&��
��vO��6ٺ��"���'퓸�����Ih�I����}������{��`���3��w��Xt�pＡ����J�8Y��浦��{/OJj��Z��鈌P��4�.��/������9�Ō	O��2�VP��5r�0�j��|��Gk�9���7g��9E���aD*����1�d��Ȱ<���H����Zީ���m@Eu��+�'S�vڣ�j� �/�ڔ�\Is��@)�t�A��+1������be��=s������+�j�m	H�]<�ut�.�������χr���+̭�Z��H���q{6�8�漣��n���)���V����с�i� Z���z�<ڽ��
�`lѩ��s_�=x�}��*" ��F�OhiZ!u�G�j������\?�\~?�(�$reЖ��)W�'Ⱥg���$�����4و�W6��;j���l�i�N�`M�N��+ks��93�ӹ��I��F�m�s��SF�'T�)�pk�f�$� �R�p�dc�<�t�*D�*#"��i��㼑�E4�N�`o;��	 $Zi��H�0�[z���q����ߚ������9�%1GҸ�밬TI�ҰR9��)쨧,�S��f���f�91>z�yiB��7���9O�w����]u"�/>i�c�G�Ba6Z��d�������.�������e���L��Wh6;G�U`us��g+c��YG��k���ƑS��,TOH;�%�)���e�F$�A�P7�oM�Rk*-���k�����
;��XDA{Z��Zx���3;���EJy�	T�����С��E�*���3��IV��ӡ{��>|�λر���h٭�:�z��Ӫܾ��V�G~�8@<��1ض��U�#K�a�hVK���9G3o��2�b�RW,0�1�B3sd��c$5��Q��@�W�n6�xy]�_��Nox�~d��3w��Ґ��T�����S�>T2#�P6F���{X�B>rH�h{�|����R�R����	8 �]�=k�W�DG#�-�/�>�@OK�E�x^$������I[aw��:�ph�C�	�w���8�Ì��D[���=ȩA����5��[S�2�P�c��-���}bɐ`��dXgSl�5,�aL�+<�(}	a�����x[P���!'��,Ÿ[M?P:��$�-ӂ$s �s���F�(��h'��cƯ�
�mW�= ި�1\�X�?Tk�)JE�u<i���ǌ5_�c9��cհ$��'t�}��>3�"o\TS�^�%�,IR��_�^y����)��s8q��F�/��i1辗:��È"��3[ߛGX�����xU���H������=�=�B�!G�hFҋY�qC�g�j+��S�A�R<C�%6]98�����熘�_�
P�`��o�S�_4;�;N�ũ.?>��-ͷk�����h��Dm��
*���s_����a���:Z:�$Q��Q�����Z�PaDF�>����5`w]0P���XV�U4&���mL.Hx�;~���X\"� bs��>!���a7�1����� E��:�S�6[� �?T�<�����*����[)��#�r��N4���=�D�J����`���4������YY�̡��ry�ķ�&`E>����k��˚���ƿ��I��؟�2��V*���t��Y�i�d��P�b^�L/����'�����f_ʕ���#�弲d�� ���ݪZ���8�_��:i���3F��1�ՙ��z>M񭄢H��L[���+�KoHeQZ�<𓻮x�'O_L%of��N�	n��~[)#��	���Y7
��k���3��T�*��]7����D�*���g��g-?�fl0�<�4�\VF.���]�M��HIp�B�>��Q�m@�'��rgAjd�m��(�,$XW���5C�!�l�>q������2�Ƕ!
��^x��%�?���~��_>�C�����׫������|��|&D��'�j*�e�Le��k��;~��@'�E�0��`�����\�^�1t�_Xaы�@��z�4�Q!��̀��0�ڐ�t:�Q��BE��F���2 �uG|���or%øV����A�5�@��h#LnV��.��1mX��\9K�.Ķ�c:�S?W��TF{
�E�e��O�l.f$�8l��|����"���(u�����l�?���D��Z�3!fݿ�ʘ����H  PR�Q�yώ�N݁7y�2�S��1�ۈ*�"׹��k*]���x�@y�������{��,���]�(r�w����06�>g���F�l�ߎPI����%��(�V�J����$0؜��N�47���Z<ƪ$�f]45d�G���f��sfQ����F�k5ǽ����)��-T��#�5*��7��d�wm�ƗQ׸s��Ŷ��J'�[�A��ɮ�[Wz�\��U���	�Y8f]��"fڲ�#���X���!�2rsZxE��Y�"��"��Iy�Ƃ0oh��Ȧ*柂m�����_K%ړ���!���H��3�}�j�u�o���ző��N�1k����>��Tk��/������M�!�`�ᡎ��!:H�����?.�����=�H��6a{�}� ��O+��̣<�� �#_ͦi�0!
�.<���x�Ʒ�)h/,p%�=��UȜ��]u�c�4����e�����Lu	�||�޿��OӀ���R����&�g�]��o�r4ix��ͥ�{/@Z�5��c����k���g�yz�,���4�plZ7�.aw�>�_ڢ�ɿF��Xmf���(��Y9���n/�l��5�%��ɿ�a�G���)��)�[{}M��M�Dwm7����[�l]LYg
|�{m�|�_7�����BEqv�-��-2���'{���2h�E6І��r��� N���Ǵ���/j�(~]faϭ�
��o<��.���Y���#�Z���͌,1ԑ�V���7�N
D5��F�z��$��L�d�����)��Έ���Ԑ`�lU�F��9���Gzt�\¶��Q�~�akf�U9��b)oKB��>�M��b��-�O{�V����P�%����L�C��c�d����iP:��iC�§��/v�>T���~lk_�����������B�y�衱�y��{e`��k.��=�#�����AN���|C�hL�����W��M�҂��IY��m����#���'OQ_���W���|��'���0��yHN}8I� _ ���J3���͸`�] �����������9��`K	���O��T����M3R���Rٲoǟ�sp+�?28d!$Ӓ�ٝ��(=v��\���~��%�36Ç��Gu�X}�3��7�B:�Z�`H��W�FPiq@�2)Vzi�����>�]v+��3��}oTˮT���4%F���ݧpdn��G���~��X��Q �bMw���
��TLT��}N+�}��VИ���IUv�\���}_F��0�z_W�D��������t�bQ�{	XE��@'-�o\�a�лGy�UJskP����=F�����+�y�#����L�'}�(꩹�Rv��|y���0�0'\.]I%[H\����sD�D_��X�ke��T�I܂�(0E�
,�K��|]fW�A�U)8]���4����^�oQ.)��_3$�E?�7yY !6 Q�  �2x���7\���t�J���hz�jB��\5� �hh�������F��]�2t<��bJ{ߊ��p���Btѹ>\�������̒�|�v�.^7���b0��	����#�s�V��37:/x��$�d�NH���T�@�^�"%U	��X�WK���XcF����$��wDF��#y����Қ�%�ز�I���1C��|hV�h�쫬-���>�tN.��	��G���z�D�ҫ����q�d�]��ޓ�k�[r��B{�t��P$R��W[:NT�d�	b�W�l�N��5���{�a�#�|Ek�D��_]U�n�7�::Nn*E�a��(Tw�9n�H�σ��˿]�1�K��,p�..�ݨ��_;a�`>�k����YS�Hmf�z��V`R��x�L�2�W8ǿ �{aȷP�
Tԙ4ϩ*ϸ����ҽ	LzF	�cs�=8>0����؟�N�Z�ȧ,�Z:�s6��̻Y���I�%�I(�9Q�Y�������[�8~p�Wܓ�Mh�s^�kX�QE��`��z~��w���]u-C|j4ȩ���*��qc��F Ή���p
�.���V��d� /{��Y�f��e�傜����YY9�b&p�-X����fg9��ղ|�S��Q���G���?8������j��~G�b��lw]h�a��A�ä[�׮��z�c�Q���κ�Q�hC�ʗ$,=�sA�+�f�������Ok1I '�݋}�����a�f�B��U�j�6B�����A�X��-OMY4�:��3������;�yٍv�<��KPh��)�
@��(��q_숄��k���mX��ސ��I>]�o4k��4iWK��!j1��U�X;�gL���j���&S'�Ȩ�����-��ʃ���$�����h���3��$�0��e~��
���m�Lt{��;�]�g���4�>���y\Ǟ(�jAb(S쳂�&C�)?[aP'�M2�y�iwV	�5灴��Z\qvG��q��������`o�p�fP��aft�E��s)Ί;bF>c}'�mX��!�Ht3?5��.�x��B����\B�*|Ԕ?zj,e�KH�\�c �
p�GV�{$����c����;����������BuXJU��pi(������b���=I��D�#�{V9�� (f	b�u�s~�O{��/�Ma([�}W��6�g��$w���^����Р5�j�uޥ�Ī݇���sZjIg_�Ѐ��~ebH�<ƛ?��U�]˃{���,���a�/l>�����H��څ����ޚG6��p��#�M>Q���Gv���!5�@�!�Z�m�7ߋ��Y�r��&������z�s.�q;����!�h?O�F����IQ�*��s�h�B�Zm��9��H��4�!��	�L&[}��0y7��}R���ܵT���9�;�Z�K��9O�t�M��{�쳥�(5y��{�@y;��@�f�h�ĩK��`�5W��'䄼�+�G�]����`?%h7x� dN�]ZfKv�Nc��7ukx��m��uU��^X�Uǁ��ȇ*���94A?j���+�+?;m��-<��}v��":�sB~����3`C��"^b&�	6_�\޴�PGzO�@,\wJ�:�,3PN�zZ�DdU-��q�%&�߾:�% �m��|0���QD�ۯ{e>��:��A�/�*�DÊq	k��
w�U�ǝ~����u '��}l?��F�y�Qh���w��(�9�E/&�*:��e���`R������FfB��黙�F�,7�`i�wJ��CC���t57�ӽӼt�\�Up���C[D�J+-$�oA��Z�B��������2�SO5��Rd�Gi�B�y5d��AB��|�5���/������c_�v��z-�y���o����}5�-!�s��������� �ޣ�P��a�+�����ot��k�>ʽ�h��Y�} �WO�*�C}ǖ�rG��_J�Q��6���n6��dH���2���Y���+r�X�+leCW-!VF���F���X�+��]��a �$�D����q����v��*2�Y���M���ҌM5G�����Ի���N�P2�1fIe���q�G,�D���|�ĥ��Gr��k��'�}Qꩀ��m�:�5]]t?Q,�a�4_gCx���wp�mB�5��~\�V*;f;q����PkB����͠��~�^�P9?�2=��+�~�A��tŚ���T�*��x�AI���;����~3�#��*�lҤ6�2����ir�,b�l��aT]A̡��6/�#,/�;���afiV��ˏ�h[��	��_�����uξ'v��<"���&EF`��h�t�X��ȟ4y���գFc����������u\�>r��q���|d6�	�n�Y��L���K+�G-�huU�+���L�䚂F�=`@1y)��}�Ku�N�
�<�$��5��?��q�*A���]	�^w��� )O�(�yVfk6��������;��D^?JCp*ߛg�"�c����*h
�.\EMb�>���."�
�}�v�����ǅ|1�LDf���%�`���~��g����!���O����]#�|���������R�G��,L� ��dCQ� ���-B�?�3�bJ;=E��rȷ5y<��R_��XI�{�ǳ�ɞ�EW-5l�����A?b��+��[:�j~ .s�P�o�v�a��m!�?�\�^/Ᲊ�Lyc��qGD�KЩ垫a{�Q�x�.�i�1����+���
���<��~���'�'��\N�Ʌ�]���u�����۽6}�3�=��U! ���﬜a���A�t5��{�m��l;y)u3S�RL �lYl�R�F���*=E���>��X�*���^��K�q�b��#(0:'�He��7�J2��eUWaom�FH�m�nܲ$o'��{�1HS�D\�h����3�!Ĺ� �Ѕ��٫P�!� l�ʢc�������g�0�Pz���5dm>���NF�j�!4W��Y�g��3[AP��G���P���a���_���}c��4Q	q.Kjd�C����G0�*�ֆ5�|$:�[��k�t��*<?b�>�֋3����"u�Y:V��!0����=��1���~8��Yf�� HC�����]�BT,��yG�p���"��x���7�W�(#t���݁#P�����(Ё��
��7��y�i���W��A��029��"�N]��L�d���e,�e��T�����~�;���������b(ޓ�
�f�Y�F�0��n�I��xEA��?|�Ȥ�E��>5(�k���[xiDJ֛�y��r^�J��f�˚�ԑ`����/���&1cv���=	��T����~Mr�_�"��7U����Ǎ�[S���kå4f,BZ�s⇛j���?�Lص��ۦ����>�v��f�bI��f�o����<!��F�i�zL���3�c"b�LH/a������u��Ь�n^�+z�Q	��w�	�X����u�5����,�O�#���knU}��sR���� ���h�T�&ybm/BMJ�r-�V���'#H���9*�X~�(�|Zjp�6na���� Q�n�)��"�j9%���~k+y>W�H
���)�5,We���'�eq�9�����8EV���c�\32
6*�FҞ;��C���;�L�����R�w_%�%�qy}�v��?�)4��(�"�WB�
�S=���;B*�fe��Ǣ��q�F �����y�f�4���x���$�M�o��.�@R��#���IRV��3պj��0�7YC���p���`�/=��	�#���PFy��_7،�N4zg�X�2���}j����nm�'��d�-���g� ��z�y�$�m^h�Ӯg�&�8�zW-�sy�D�[���ﰯ�ӍlѲY��k�?z�MC���͈䛐�d��gs^���URG���S̢�*������U��q~���-�=�<��\�"�@�rnl���:�q�� �T��N@Y�ƣ��5V<��O�&ł�yJ�6��f��Y(�2ǳl�F03k��2���.�5F��<��Ai��J��;��ÅRQ�3e�t��<j�F	�%�
ɢN�Eʬ�S��ٛ�wD:�]c�n��R��K\#�a�AA�
�g�;�n�|lG7���|N�˩ 9���!}�Z�@�?�,k[��i���	�� N��`}��5Oh��Z5�r�"�+L��|t���A\٩�#��=b�y�@Za�"�JG�Q��J�O��g#�z64�`b�מ+e��Rp$ɸVձ�_��1��E��
���T�jKf�Rz�Gݙޫ��
�!g��^�� :d��8�S�0J���ѻ�eԕ���;x~�Lb�%��Zv�Ղ2�!޶�r߾��R�y����0����S������s�*��Nt��Fô ��0����I�d
!�Af���J�p����w�}De��u� �>�B��n���C���rj��0P����u���~	�V�i�� wvT���'��D8�a�i[��Z��2�f��د�,�]��J��h}����i�=���k�4�u��^zIJc	-�ۧ?���Je��� ��?��u,6��/���p��k�䨨��9��_�0lR�T."���wy)T D����ًxC�#����^c6�F��5�wh80ŋ�(gm�&�6ܡ֌�F��O��i�+�Fu�|��c_Y�.�?j���W e_G���U��%��0U�������'�=��Q!��:��0к/p����h`�<)H�t�Ó��o���8^�=�ZԚ�6�w>j"���;`��%'�MjBSP;����G]Ea't��"X�U@a���Ӫ�C"�RrD�q��U@�:���~j_2/ $ ƥ��c4ߗ�yo����y
f�R~O:_�]�5TK��<˰4i�c���&,)n�f����m��~�ߜq�us:�z\�Q�Z)��t߻s
��`����fڂ� ��4|�8�㑵;�T%P�G§=d�00�����i��[���=��u͋��Au��� ��½�^Y{[��Ǧ�}�K���]�����6&�m��jI(U ��#~"�O�h��o���?E�o(ik���e]f8�*"'�2���q͸���m@�L�8q��`�#��XB����'R�K��h����q��Gػ^���	r�tU��[t���В=y��'G���y� �����u�R:9��u__-�r14_@�w�0;�v,{�� ��W�'�����g�r�7�T���,�-ͷ�YZ���k���m���ө>7jB����5[9]C���I~���ݡ��#�{��n�e��w���8��I_���c9�^ze��"3b�Fo��X���Ы�Ko�[�>��l���Ag��z�}揺�o	����̓z���J�<L0�agC�h����1{�AN��A�~��g�y��E���e�C޿�� >�Hn3�WE^��d����i6ŗ�<��/��Bе�А��4�̤��]m�M���X�. +t`��y�Qa՛ԏ�~� Fn?<i�2��#���������\{$�lc �Yd�Ճ^`@aq�����p�.k5��?]���ޯ9�Zq4'"�KC,���L����Hw+�Qz걐�L!��OŰ�V�Pnv�sO���ZS�T*9�^s�Ї�Z�K5l\�~\C�� �4|�������(:�p�o����po .z����	B3��6G*w����oʬ��)=��r�Q�~�� BG$:J�a������п�t��l����˵�[����Ea���Y��-
��+1�r;��m�@N�8Si�_c�Aƃ�Q�(CMq�4":��z�#��2��ǩ�����#�0Z�eK�M�.�09$i���|6�ǯ*veVա��O�$r2��r�G2O���t�?T����k�lcbD�. y{	`�p���w���ۿ �,_�L�7���x&�v�e�ʷ���z���L�~��Tg}�pp�c+�P�D<Ŗ*�!�O��$�fg=Ůq� �$d�-�L�UP�ap3l�1y0��R��pBduv$)���5�C��i�/L�`��)UَZ#��_����j3ñ�",��|�W���`t0��]u���)�g��N `�\|T-G
���P�����cu�cjl��|���m��&һ}�0/R���:�M�|�\�]�����z��%@xw��f�i��t�aq����=}Q7p?������_����y ��jȯ���l��v5���5��sKbb!���a&���L��0���-�u�BX�I0��G�"�/	0G��H�(~��z�/��^׈��H|�`�2&��-D��<���c���KHBE�>�i|�r磛k�D�����,~s�
JOBE�`�lա��ѩj���*�r�?������;���3yc	2e9��A�lLZ��1���L$��")�Bc�o69��~v���hU��yYm����� ���pEg�Oa{Db��	D]+�&a�"�p�Cα����GJ�߁��.T��<����Ț�n��SͱO�V#�(q_�{�u'b��߲��AN�p׿'�:D%��G�f ? nM��R{sd�&�J�s@I��5���k��`�q�L|�pn�Pk�Q%�eY>��0L	��X�~��:���{�E�B�K�lt���s{|�r��<C�j��� $�)ʁ):�U�~{+!zb�`�r���@���{��A���+�V*�@��ܟ����>�}qZ��F�R�|
�f��j����a��{�Re��5�6�LE����|�E�a�Ǌ�w����'}��D��~Z��4�=n�x��.�о��{ˀ	�}�ђ<�<��m��\��l���S�	L c�*[�������: t�7K)g�H���F��Q��A��h��Did���Ah� ��@g�F�DѸ�5uJ�N/9Ы��Y����FO�#7�#���<5�����wf�O0�9�2������}��iԂ�f�r��2-��j�ɣv�}�x��;�"l�R3���V�r����/��6"@����G˯n��%+�j�&�x��W�-u1��x[�]Wyx��@�Ia�iP�Y���>����������j⟬*ƚ�9�s{���D�g�u^hĴAUh��t��dj��&�����`��;��t]it�������FP�pfmy�~Њ� ���J|	e<X<;��F����֕@Y�y�F��r���hϲK܍�A�݁�N�\g�H���S[�2�� ���&��@����e`�������� oy��AC������"B��*�_+>Jq��_=��u��l��sGBZwT��%8k�X/��RSznа�������0�KAT�S&�xtw4�A���;��������}����1��o��Ε:���S��i�����a�c	����0�8�9(���R`�,��z5H��W���պ�p]������5�Q�߲A �K�F�[��t�Z��%T���JU��~'�n��Nz���h�@Q*<;A���B�U��
�ː��e��{!�*����N`�U^Z-xܡ9\�jr|D�2	��$[���@��{p�KC����2z3��ظ��<=�*�u��a���X^�OE�����ᣅ�ː�ǟ�~�H覙��s�2�-)���YN�������9�o��B�!M��{��W���{�5�9����Q�/��M=���N�o!fJ�#r��Q�IAAD&i��R��Qi_ ���<��)g���r���㹱�.A��3��k�� ��kW���6v�-] ؚ<���}�W^hI�+֧����]�d�����
n��G'1HQ�i�*0Ob�I�ӡ���@7���{�%�O�\@1��2=fF8�&��d����}�E왜�jL������#~�oߟBd�w��G^MB�n�(��5�J1���HL-���EqA�B��I^���K�{�$ʤ�(Y�ğ���n�e���8ㆬ
�Q"Y��������^ڃڊV��Z�����^(���i����Z���=ג��2�����
�#��H\���_��d�T40�C�	��V�%!8gD���5~koY����$��ˀ�e��e�y-��Eh��y(��!ɮ�a}5{6'5*n8�M\���Sޛ���I@��;�NZi3	��[���:�Rשչ+��t]R~y�L�3X�͉���0?I��X���;��%L6�zo��F����y<r����2��3�|������j�*w����c��B6����$�4�eu��Ũ��!A�x��9'��GUN��m��_XK�-ޜ62IЋY�-s-�{{�.Q�H��:�0	���O�\_��M�l'?�V1pe��;G.U����l����v J���R_���!��k��Y�ި޶pQ詩:߷��1/��	t�4�Iw��:f���{�^��m3��hS_���-���*���Hp03�X͓�:�C�w��;���N�x�B���xa�������vVӪ�����_r�\Tg��Դ�,f���V��/�۵�M�n�x79g"xpk���[DB�Ϯ[�������:��~wD|���ծ�ׂKg��)E�=�_7����sԳ�H�����8�o�@Ѫ|vb�S�Y�i����,����<�ÇǢ���Y�'�.q�ah�9Y^E�!���>���{5vغ�]���ͬ�}�k�=/M��Ň�g��x,7,&k���&̮(��zk�R��n���sU��ͳe.o���<���	�~��⪗�i����,f�����v�L�	��#���<+���H���\sf���X4��KG��	C
�/U��o9�г��e;�%�����1AucC��3���/z�)4%�-a�M)˔?�� Rm����血q��fy��[��J���۟f�P��Z`mZ�8Y.t��vc_��Ib_�R]gɭ-yC]ͽ�Gڊ�����s*�_��KXaM���k�L�ه��6Q��ܬ���NRae�C�Pu?�8�#o��d��ϼ�ڂ��˭�Ƽ�Vd0��w�|�P�d��Z�L`�U^�r�i�X��	�S��~ARy��I�ƍ���J�ک>�s�H!h��kƹ��{UIj_��>T�g@z�Q��G�rN�Io[���r}#����z�����J�^uO�'�*G��GW�f�{Ͳu�U�����b�����e�GQ2�=��.>��:J� �x�H�����wF>!�Yv%�Yp�uH8����/��=��9��K��-U�ٿ}�w´�vbX� �O�����q.�o�v��W�o_��mN�Ζ�t�ԄT !űܓJg�W�+���F)u0��S���L��\���{�H�����=�oMc'��4�N�����	!C;B�t��R��t�HncM���,�����7as�b_�J���l�J�����	@����.�	�3��d#��C��[ZOD��6�$�f� qЋ%7T�r�D�[~7�����^฀�L�Jy���b6V�5��`�w�w����Z�I,��⣀X�G2O	"�J��L�J�t�8J� "!��������������:��`U�Y�D7J�����ݿ5��KUWI�̱Q���sU_�1P��0wK�!���=���e��C��m>u�D�J�����^�Ϣ�|a-�������ؤ�U��ٳ��"��[c�8�r�C�]U�
�z̬>a��o����Ć�cy�g?�kr�r��'��~��p� ��b�����-���8Y��;������-l�L�wS/q�>}^� v���� \1@�czο'%�ױ�����P�-{���qA9HާR�DN�g���OY�1u��o�9?&�a���П<j�@�rk_KWYj~/��_��;t��*�)��7�'"'������6�ߚ�5�v��Pzk���L�ɭQ�B�4�.6L�w�4?��~~������Z����g��+h�5I�=jn���(�֎�����6���'�O�>�T��3y)[m	K��;ԕe��f�&����Cs��b'k�^8����N��S(�,t���p*�c�w�n�)� ��I*�kO�����'1?2_��p���c@=���~����P���h]�z��7k̕��,��AP`y�S��z�\�u@T�n�/!
�&�ylXW�4�
](O��k+���G=/hv�BBkX,
MJ�Y�^��%��9���6�|�fN+���u�� ��|f�U]���o'F���B[��Sz�Ϭ���z��N�����s7H<Y�s����@>��B�/Q�:M8l ������7Z/��F,�����V��#�3�%���3��h ���^Dܤ����Z�~��I�hP2$WV�����Љ$�~�֡��ّ��cl�ky��@}|�V�=�/�U2u]���>�"(S��56�ڧ�͗ҶU��S_�a�SR�|4_���D��Wm@g��Q���AD)����!Dk�k1�����gD>��ń jWN�����iG���8+q� �De�*���y�� #�!H��+����-KjV�d���r*�X1������Ԣ$V��L�|��qNeV9���2|�z|���HU�-�<䀛�g%�zQ}����dTd��;.+e2��Ig���;�Q��l�)L[4��ۑ��*��~�A �<5��*�0m���-�N����%�ԣ�|�s����w�^Yn�\x���;� ��,��'����n�G�x�aƧ�g�r*��A�1��;�Eԏt�������)�"N���%\�B<}�\oyo^~��ڸPg&ǋ*�jb|�N���R�����A� TZ��a⊭���ۮ[;���D�U�S�-��+��uET(~v��t��-�x�l��kؽ����&��N���<@J�4Y ��?�	Z#u~U�O��k2�)����7<S���k׈�KIquȧ>�if�{�b�%A�N<%=�ґբ��<]���} G��E3�P�Ͼ,x����:]�W���?��h*�w���K�Ebm��arx�>}A݇��u|��A��4�ؾ�Fr���{c���cv�(<���K;O�_vy[�g�F*S�:��nJ8��
W;qN����5m��������j���@+�.[o����z�)���p�G�2���3L��]]B���;^�������P�q���"$�w�"co��0�~P���! 잳�l���7�>���%�pu��}���׹88x&��t��P�� P��q���,�����^���	J��A�i�נ���s�i����E�j�55���[D�^!��MA�sȻ��Aد�ә��;���f��1���_*r#�s�Ҍ��l��i�@�*r��{ԴM�	\�3��dOผ�� �v�i�GV�Z46D�:n�ZLs��Q1H���V��c��y�a%����/��᠑Չ�Ԛ���b����W�(?�z��R�e$�^Ǻ�@ft��Es:�B�!h�!&�{:��Y�V��n���a��!�;t}����5�������Rj���� 8��
��i����M�����S�U����@@���[w�uj��&W��u���E{��~p�n�`�������:��ײiϪ�� r
eIEb���y��: r��{�E���82sE0��8&@�J��(H�aT@��@���q�$ �b���t�A����6�dhr��9U����_��/��Z�.ƪ:g�����g�*��16��#�>B�ƭ4O](�D��y*�W�s�Q��Es鄉�:W�?Ij�W����������l|��#OU䢸���� 5N�Ӥ��Mx�!M n
����/&&>U�F?�Y�8�>�	��5>�Hf��v-t���Cv��u�Dɳ���>z���'z������L�Q
�D.��j������M��hc�����%PN�1��I>���^�׊q+O����!��|��Z��dX4����� �Z����(�N��ڬQ�����vv�	�j�A�ϡ�fU���eUA�~''oA�.�$u�fs�ʇ�R^/-F>�����Z���A_Y8C{F��~0���.�^X���@R�Hq��H�C��&��7�[����(˗�i��� �j�?P)��ZCQƞ��4�F"�͌��)��1�_R�ߢ9/��ާj��C���e�Å8&�������G95@� B�I�8��4Lw��|� ߆�K{}!��c/���A��-���N˧�xl�|>e���U�둺@���	����.\8���֧�t�g��`��kLl|��8���A�����&�Z�m��q�#7��E�86�н�����PY����>:o� V|�&��1�c[�����|�mBڗX��:m}yױ��HȒ=� Ś�q�}Q��uh�x�xg5tv�Ә�9/���ve��VQ$&n���8�X�n�?���qA�6�+(7��6���2�Kq\:L��1�����tn��.�$G�����{��)�/���F�MT�-�����E�s���pB�^y�,}
�g�o�̺,|������X�N�;����]�ƛ�HJ�7�ThtMAr�n/���j~�~4����P(����(�t�p%r�vH�@>��~���j���Z�=���:�͔�A�r8�H�@�M�����9t��������?A:o��)��ǫ����zty�u"ȴ����)k)c�S=�HsG����U�Li�N�����Ȭ�e�B�dz��5���ª�w��ɚv7P*��G'-�*�� ٧����n��c��oe������4��+��<���s��*�lu�	M.u7K
�zϹ��k�d��x+I�.���bD ����&�Џs�0e�u��N���}�KA$s�x�	s �v�k�(��d4�&sG��u6/>q?n���:��v�>0��� �����Xؗ�M��~̧�k�ae�b# ��_�����P^2�R�h"��l���S�ڦ+�=�O��}m���?N� �-�vay�*�����-yF���!|��#Ӑ�_�����<NG}���AX����9����C�&A� �Wޟ�(��:7ydw`�Q���RՕ�gzz�\}�|iq� �����$��@z��\�r�U�#ਝ�o�������vY�G�~R���@i��;s�별��8��Ey�]����/V�|o��]�$�����+®~㠲6�j�w)����{ޔ(#�0��s����d�����j��|��N�/�nϋ�W��ԓ&��j��WN�� �Y��Křƛ ���jεq����	�╫�"h���%,(=�0iw�Ջ�H�w��#�������p�����g���C�U�]�ۖ��{�QU�j}=�r D����Y6�9է�Sչ��%_J��̏ �	�%�,x(����[H:ICtS�&��.�y�[��s��_�207��W��S��f�Hbu�.�OD��Cn�#�* �����^���R��Rl^�U��$�P�{.i���W�#
R����1UP*�<K�{46Jy-{�����"�����zQ�~k^��O�Q"MZ؁� 5������;���:*(/��C��k��(Q�g����MoJ}gG���S�}%L����& h��AR_���6�__�vr�RP*,n;�s�O��MM��9s�> �ȇ��������W}d,"�#��Tlr��]�ڰȿ �ʾ�N��.�e��N�$�?B�?zT%[P���T{��K,�7;~K���q��-�������������'���ؓ�ҷl�������h������cN;NןY���iX,��o���^�s�JYӣ���f��n$q�Qy_%�ڽ�t(jjEU�%o��u�m8��\]�4�ƍIe�76_�n��6Vx��Im��9|�[�b��3�S�[��W�,��p����A$Ҥy�Ło���K��`�X _L�rX���t�h1�����7�8Y]���&�~>�섋'B�]�k�Ȥ�Ak�M��i*H(B��*�1�e�!I��7���bV?�Oۓ6�^h�uF{Bq����	�U�N E����N��)p�6]�����n>�E'�8��S���!���>���۞[��I��EWE�"��Yx��Nۮ�>d�9FuG�ĵ��"���yu��K<4<��%���g�K����V�Y��S��J?��lEsI��v���'uS���Y���Vm�G򷄽�sm>[@9���ѓ�9|���GWzT��)�85S�͈l���D�����:��,�r��'��%hv~�n�Y��4l���Nhp���\�l�Y�� �'� _8�#'�Z�/�#���ا��9��[�p�E��v/FG�7��>fe˕\OJ���ߟG�xNMJ��e%1ڃ`'R&.�S�`�B��.�Q������-?���i�w�oD���?@
�0�x>ٙ5ݏ4�(o�m�{MB<�:�v�{�κ	��V��Y)��k<����n��o�^�K�B$���&QFs�u7��i.����ȁ��吢�6�!��$6j�i��،QX�X<:�� ����y��l�~��gAα��!�-��_����z+l��m �B�?B�*��Mg�n�:ru�˄��n��]�>^	N�>�f�����+��uҙ8_�''�zW����&�]l���nu��Ǔp����;�ޭ�F�|ҝ�wϪ��/�m���C��L���7���Y)s���'�YI�E���0������l|�!2��:���?{��q��sk�r($�ԇ��48�~uJѕ��#�p~��T�C��l��;͢���z!6^G��9��҇�:���u^H'I�H滤�J��s����$7.x�:?���kI���y%�9Зڱ6zQhf7�.���L��F/���/`FjQo����&�Dy[�f�_I�O�)�]ob��߀����F�6N���]o+7{�������,���g32���e���/f2�"$12���yO���=	�p���U�Z�riv8=���2i�2-��[$~�߱���]��p��BFQ��rH� S̦ӓ���	GA��壟�k���d��- rg�p`WZ�DMsE�#�*����f�e�ꕽ
ܥWƱd�T���)1�(����7T$L�����Nn���|d_��z��z�����v���q�1��NQz��B���k�B��]���G6�8��C�J�A�{I�y=`k�S�A��B� ��w�]�?��/��0Eo��>��e��0��c���Ŕ: �;+��$��o������O4E�먼=O�6mH��<��%������%+���0@_M�	'��M�;��?�I��p�$ǧ6�F�	� i�]Œ��UQj8G��с��y@�#֖V�����z4�P�y
t�g@���q���!�+�S�N��y���SB�̂i����]��2�W&��خ��u{%o��x����;E��ԣ���R�O���J|[�@��P���Y�q�Z��-��d�C�ss�u�-�Ps�L��.A�Z8\��g��Kb-�^fj3�,�31��L3��bq�z5�_q>�t'��3 ������,X�@&[�Y}�^�Z���.�7*ڡ�aa٘?��&��UVeFa�T�.Hfm5W2oI�����3'#�_��LB�\�d��rҭy�6�4��{pN��C���{d�_�G`H�X~m_&A���2Ǖ�fq�3)���,�/��.�u��	����.]��ܩ��+�u��՟Q�˷T|Q*��`��(�&�������(����`���9��{�F����Z��X��<�����=���R �u������y�*��:$)	�o�Q�R	�U�����he*\����>�Q���c;E(ݥ$�4)�q�{L!gŁ�͛	�E�w��D83x����h,,��/i:�A�@�w"�]�u]�ׅ���63����|ݾG�,������欌����B�A�]���i奡��^�A_������3���ѫe�7��<(@����	�9�Q@�M"F��܀[*=F]J՟���I��׮a�1N�%-:��T�䖿p@�#6�v�~z��0P���߯��G��f��~�"e0�qFSO�0�Pl��ˤ�Ԫ��`$�� �J��S?􍣀�$W��W���T:?O�É[Օ��D���m�!}�-��ֿ�[��B��2#�9��>�g� �n.p�(g��<�'����B���0o�%K[��a^��2�Sv[���a���[ ���Y��ֳҗ���MuB{�Sq.y�Z�' ������:���Z��J<§+O�AUZ����Q8i͌����'p�wO�_���~,3�N����@��a��%$��/�vP��[��u+O��i
=��r��ڧ���D�r�mA��#�-�B���d-���*��S� ������,�2���L�7�%�����S̩���C�N Q{!�̯���T�e��7�~�N��p]�ج%E��I�pڀ�jG2�����*$��]I ��$��E v1u�<®��;�\_�E2lC
��vg��\C��K�;o#pY��g����g�k�J��9X�j3��� E�\w���g�*�z]8$��"�bg ��o$)�Lʐ���}�AI<�i
w�$>Y�ʰ��}� ��:��?:|�=�ϝIN�ݏ�D��v]k&A�d8E>�����|I�͋��K<h�v.:�muf%�:�58�ȧY��b�6Ԁ+<du[�x�q2��!��[W��iB�<�� �iݮg�����ӂm��� wn���ɬ%�\D9��-_]O���h�uM�b��� /��Q���_F�$�!.�jZm���w����_qu�K�ɡI
����	�=��,��Q�v���p!��,����"NN�~ѵ<d� ��RAx���=�����k]�ɇ��tt�
+�뷸�;�S=8�L��@n����T���֋��R9�u�#(��M��j���T#� 	^�Oߡ݊�C�=�i#�����#Pa� G,!��}��7��~*���������>�-�b ��:���.j��FeoWQ�j�-��e�"[n�-���Rn:0�Ӎ�^�$B��^�(���6$ܧ�V� ���q�t��b�U�����pokK9@�:*�j�������Vh5���Ay��)��n3�X��^�iZ
7p�J�ƚ\P�A��jƢ�oc��c(���6��9���ihX�V9�|c> �M�z��3e����+��8��Bn#�w&p�����Z�d�yU��,������a�'m&���~4x�RO--�+�N�3�N����E�D�"��j+�D����j\�Bg0l�=5�(g4�ts��+�>��2�Ek[�	�v�ӕ�od�*�L/��i��&�/�f��;�p��$�f���j%�9��
"`�2�duzm�()m%q�4�irr��0lX��{8&��৵@�������ڳn�l�2�����+WϾ��d}S��[BK?��o����Jl��$f)J����嵻{��C1�K+�*3�cZBJ����@�ì�<���89��]C�&]w�4��Z͌��\���cR����E�~f�0���U
�������BPS(�cRj����-/�dBAQ[~���A.���4��*0� b���w��0��n)�_��K��nvjN��%�҆k�>
~��>7k�S����~q=��V4�Ք�;<�����ͼ�f��#��t�#�eU�����g<�T��B3��Lj����aM�' ��6��k����/��o������ �Uc����r>	��P,~�罤�$����G�m�r��
d�$�/I�>�=�����B6�0R)~�����(�ˋ�l�S🖟kY0**hU�
X�%��e�R�(�K�j�>�,ml�P(����8p���4$r���mEd���x캤�Jc�1M?{.�VS�8�(��+ �Ճ�����6Ȋ��K�.G��}��\�|������uP�(Gw����?�v��l�X�ȧPTV���sf�	7Ɉ#z�nŗ���C��n&��ОH$w�]~���P�Dyt�w�C����g�3��t��>f$T3k�9�A��9�<8!R�R�gpf��:��Lu��F��:D���+�����u�����W�&�1&���6C�)6���c�DT	w�By��8�����~Z�z�!&��%#�]���$P��w���ؿ�I��/�� ř9�A���֬��%�Z�{PJ�RJ*�m���*e;*5� 
��U|��P���\�&o$���<��a't'��.׿�����vγ|�p��ˏ][��>n���FҒ�2�z8���_s&6Qޖ���w�we�5���u�"�v4��Ш�Q	��T�v�����p�'�]5i
���q,;S��e����dD��Zy/�6%2!���˼�|o ��:y~$UG�Lo�7�[w(A�	[��ʙ�	�A�dX	�7o�dOqԨa�+����#_��d0��[]�KNÎ	�&�8�39���}�gl2��|���|GM��Ʒ�*�=b���˾���^�%��޺lo{#/�-�$O�2��Q��݆ks<
*D�^�~�O��T&��8ny��c=t���Lv��QH�^�U�f����w%<���<��δZ���<o��w�.��!)ÉR2��B\���݇�SsAƾmf�Hې��~��Oq` �ѯ�ߟ�;�x�!]x�	79\�������d�Ƶ[�Hg���s\��:M��D��g�R�<y#�㰠(|I�e�,m���b]�T�	ŵ��2��.�}�QA2;<�n���_�Ar@u�9��Eƪ-��7��7��Ѱ����%ʿ�i��DK�l*MH�i���"�k�9V~�
;�3B�o���ʖ~��L0��$��L�]sȊqa�/?@&�؜�ޚ�9< �N���GM�7�n��b�$Z�� �4�Sϟ�愘(��*X��aO��?r�PK�EFTJ��������!��O `��
O�qUd�ۍ�W�5�9]�b�LR��G�	ܛ��Q���!h��o,�|-ކ?��@|���5��[E���a�v1���Q��*ʅ�-rی�KC=���@���F,mzE٨xA��ī|���p*�F��6P}㇗�P�_\1���������N$�k�B'���a"w!+�k7o�8T�P���V~7�:�i�U������ЉUO�p�8������t`�o�Í/I�+p[z�C���7���'@��`���cΗ���3Q���D�(�*1ݺ7?"��[���O��p7��U��H��#/Hp ����3�q�<D�|B������w䳦F|U=Yg����̚�\iN)-�b߳dt�4?",~�	x�f��g^t\z<���-��~
�]��vF1�&�B^�|�_����"}��(Jf�qqwo�6��j�,�qH����'��I�.~�-�= �~����Ȧ��D�W�#.0�w;���Ӌ�07q����������)w6�־��($�M�������Y!̰3]H`��R��0�;!՘�N� -��;�LC�i��g��_�Na�2=rF����m���-<�&5�2*D���������;o?L7S�F����p�F~�0Ʌ������h���&��#�!�թ�M�_�o�����1
t�9�,��=R����_�+àl�]P����{שZ��H(e�ȘC�x$�������M�����<� �^��J��_6_j���.b�Q#���۴�y !E<��<Cf���#��{�<�E�p�����ʰf< ͊�˜/�S��HNS�1*�P����R���������d;7D�~�Hƒ�9) �w@��[8��ҧ����r��Mya�nٔ��i]�Br,�'8�<�y�ϓ�֔�;����j���V���`?#9C�ÓmV?�@QA4J�n��	n��Gc�.aw��,D�إn���n���Ƀ�=IW�P
��?�b�$�l`�W�D(g�����E{�p����s�Cۆ�|n��,���e��tDqq G���[��=�0S�뛋b
�y���m(w��R��iE]��|9�i�9�j�:Y��3��Q,If]�t�%�q��T��Ɂ�46�w{��mvK��0��5�0e��:��(�c�f�����Q�$�.�2��E�#�rm&� )+�\]���߿ϴ�W�A�`����*�����^���2ZO3�>h�U��K�������K΢
�T6A#��8�.>�S>�9�ӧ����B	SW���aH*�V@��N�t���X��&�����Cn���{j�C� ����zv����)_m�����n7X�k�3᝻�����L�y�8*8j�x�DW���E�����y�na5*���2�y2�ij���_�f���c�qt���I��6���f���S �Ct���H	f��m��δ��7`%#�e��־��Y���5J奾���)���}�c~�!`�	5N�������EƢ��?��d-�c��OTHUeW��G`���Y�� ���Rq2��<��\���
K��!�֎��i_L�Fk����Rb�|f0�?G$�����ל����E%��@M�$7֕(g 翲��^�G�d�~��BsBWT�H*XB��ڭ̕h��f�5z5% 
� ���7(��zRr� ͅ�v^5A�]=`��� !�grA<�!�'����im d ���@v/�ε!�kg��ȡ�������3H8d��O��ѵ�(	��4�D�s.b�M��
�D�l���,��C�zγ	�����郞'+�	�fL�}s���*�����}p��?,�&����T�w��f1�N n9�:8�N�?w	0�\��W�
P���Eg��@ß��m����Ⅸ9�~,|�+*I�T0Cҁ�<@�Z�����G��a?��fDٯ���ֺ�=��2$�"�$�L�h3Y&��O1j)�{���ֿ/{�!G����1���m2�.�����o�#԰]$ې��/�C��F��{r݌	T�͉W!ַ�'��)��A�1��5l���x�U�L���fp��-/��4�@m��6���܃�2�����'|�x��nm�6�~
S�轗�s�K�@6�lLu�ԏ#�9�  b�yzm	Pa��b�� h��'w�Hf-+I��j>�7�6��R0�T���œE��-BD-9ņ�5*�`-dVW���P3[+}�F-#1�M
@/=є� 6�B�_z\�{'��`�������j�:#`X�d`�%*E�	^�z�)JZ8�
 ��C|�w��fd�G3��R-�� ٽLȗ�	ڇ�����N�:���*d�h�^דe�"_���icV���`�ȔKX����"����(�h�Q�"��xBsY�\��P�~dw�^e��|�SE����,S�n^:����3mm��$+���vzX�E���F�Ov X8�ι ���45��O�e��õ�d3�G(�C�I�:c��m֮!�P��\��5j��M����}��o�=��
d=�9FC���"�]��)�#`B���O���,�8�z�;���;�ȁl�q��D�̲|����[�A ��������:>�������c��JK+Z���� 0�-���Y���Ϭ,� ����,�}�\����}� )֞�}�����������
P.Cy�W�K��k��,��v;Dz��M5��w����E,�"����f�S�|�" ��?���j���w  ,Ew�pml�`~C�]���Ba�L���z˷�g��7R��o���k�t�e�e��ۃ�'�1�o3A�� �H֝�����"��7,��n�[Ѵ=�I�E͙
�"�{U��k��]sr�qS^`�~�r:�>U~��o>iV�Di�+	���LO<���4loe��=�hL�9C���ٞ �\u���?����@��!(���DKuI!���򲪢���@V����Ϳ�௷�� ��w�&�G
GQ]�o��L�{��|�����^w�j�N��[W������bs�"��`^ 5���k�Ji�Z�h� F�?nY7�_�F����ЮV�@���-W@�;Fq��;ia��~j�ϯ4��v �f��jAR���/��a}A(�Q��&���!��|�u�M�
>6{��m5|�du�pd����
1��] ��A���鐏�7���n/lt���|}<�7��O�|�Ŵe(��\���@.�H�Ȕ�L�Yl#q(�.����m�@�Z�2�i�:2j�ζ�>�fBy>#�X����}fT�p��Iv!�Wˇ8�OUz� .��u���$�a��Iݗ�Y������~|� ��oi��fQɧz�Wm��X{U���?������XW-�����^ܳ>�b����=���y@�Mm�	j�i`{)�olEr1���&7/�6��*�2���+�w��}|�Z���@�w��I���F���[�ea%5����pdgi(硐�ζ�F^p�һ H����������O'< \�U�� 1��`�0���#�O���?��Nb�1=0��Uo�E���i#����b�"L*:}q�����`��6�г����8�{|�hw❴��1�8��\A�Z����#��K%MjFAq�L]&C{�}�$�F`8�埳��R�vf���Y��UJ��!s ���p�z��8�1(�E��D�,� </n86�t5�H�~�pfN�|�q/fk(kSdޅ��P�a%��?�e��qf��)D�.��<Q�X>h�X>&c=ٸ��X{:H8/����㏸HKב������������xwD�G �{ԗ3F��ڏ�o�3Kb��o��K�H
�Vב-��K�,����Pi�A&�b��÷��Ϗu<K_�K�q̺��S�l�޻�9OՈ���������4�u���颌��V�x�\`��Hz�wF��uO�������؟�[�d���i4�/>6�惘�Qr��pȪ��r�kౡ�(��kgb���}h'�ߊw��/�M5�h�ixAw]I�u9�Zҝm����D�%ŭo\)S����K���?�t��	����˭��-\Y��9�t���<㿲
+��+n�=o}������er�Y(�T��moV�)��ɠ>4z�]�Ԫ=�H�P1����y,>���n���(��+���x;�Bn5 �*rn�
Z��+u��_`d"�'�,s��C�(���5�~�ɣ����Nem�W�����5m<G���TI�x��=���	تwe�Vp�;S>�֢� +��n�Jp�a<��1�v���0���oN/x���@D;.��8Ca�|ES :eߑ�f�?���(�_zI�Ɇth$Å��t�k2*d�Ζ���'��]Vti��x�G��f��|(qu2�7!LN�cmlhq�,#H^�b�����B��C�48q;���^Fc[��
������ן���&{]5X�O��V9��ڏQ+^7{�J���=%
K�M�x�w۸�x�p��@�o.����4�b �DT�-�'Ʋ�M[�<�u<��dp�PEc�2�%����-�(��������s�{p�����[ ����yY�"�8ye�N����^_���ɻyfI|1 N���7��7��ί4/��0N��p�����~��{}���h�i���Ӱ�k�|L�d��;�F!P�uߋ�p-����zCgI��q[������`y��ȹ�+�3��3���t7���.{��6��
�w��xq��J`V�
h\O��t�ֹ�0��S��]�Xb|��Xߵ��ɼJ*���n7J��3���QI����ڱ���ޜ������?��W����^�yt�=���ª����ǲ�����<�M}!A���#Ul�+��^Ge3��{1�� ��0�g��_�8�0X��?��Զ�bm���	!J�9h]=�����k��&?��O�d, ���1� ���6��a6L���?�o=U��2nl2�pP��h�x2��Gb$|��/��D�y�I�!#"1,��7H���9�T��H�A�j �;ί�6��v�>M�������j����c�$����g��4����-��x/H��O����"Dʥ�t@��q0D��5��?}������c~����#_�)QG���9q�}�9��·���ќ��z��p�!F��j���i+�z8������S-�	t�{K�a�3�YG����x@��n�+�#���A��X �?C7�pZ��S$	pySC�|%�+�� ^��?��Z�8\?LAG�~�a�!���k��������y��x��+߀O(��s2�����u��o\h��0@�2b�ۙ\������x��9dq �"ұ�x<��5+�NV��	�v�9lNSX�� �@7ކ�S�>��4!���7; �Q��dV�F���y��c5��d�<
�o)�c�!5}ݡ��,��8ׄ�_J�$�5�y����\��)O0Q��↤b�~K�����N^pm���VT1B1��!�@�R�_��2B	�e}��T��1/����8Ǯ����r\��(+ �5((�I�4�n����i{R���Ձ�ޚ%� ���*���~t�	�t� �sdj@1�x�'#���R��c%�_���梻��̀v6��Dy\�����3mm��u�"y�m2��?)�f].y0�Q a�8�j���y��ZӠg�=<U�փ�jc$SS�=��A�ǁ���i<�i�W�2��] n��ټ�T�h'���mX.�(8���o,����3߾at���Sl� ���X/3Fݏ�V����«����Ҁ�H���[��>��3c�.�/���0y`���?�s�t5���X�.���500d�1���[7[��V[7,t�Ǚ$8��y�gs�hŕbƶ-tiw��sve,C�^���!��7�����PX���)��9TƕE[AS�X������~	��3��;U�%@*f7�?�\(�����^gCۚ�$ ����d_Q0�'��>Q�ɯ��dC�����kD��?�vz��g��\��Ji�+:�z��x%�T��_ +�&�@9��2۰��r�#��_K�8�P��7��.�0m�w���_��/���'�e�Y�d{�䍜$gDQ{]n��m�
�s-@,gvt�\el�B��X�c�N�ݥ<͏����]��G��������L ��|�����$b�Tݝ�c�3��6~�dK�&�u�������ף�(Y_���o5_���7L���]�Y�1\��^�Ȟ�	ѩ,��?G:'��>��Ͻ?�d��M��(>o�F����YM���@"�'��T��]�e�Xμ<���R�� .m����X43.��im�!/�WGǙ9jr�|*O�|&�������O�(#��BP�����vp&"W
�6Z�#R�#��,v�-�'9K�q+3�C�wz��!�'�������o.���s��c~�:R�:-�3����Gz����4M��'53�m�&gJ��Cc?P !s�LL��M�4�Jsy�">����^��:�=��pѵl�)�:7?��,3�����b O��d�:��*�A	(�6�?xB"񤦟��=)^+��U��,�O��L�]<���D,����l�R�]�.7�����e��*Rp�<I�d`�s�d�I�8���|	s�xTz�Z~ .���I �:�e��C��%���	���N@�&��S� 边��N�r�@��n̡���*�F~�1X�9~X�� ��]�W���L���9��?nw:�����$m�q,��݋�r������,<��8�`���ш�z-���oy?Hm�\�<8�G�����ځ����3�+�{=�� N����n�N�� ��^5W#���5,�N4��| '�f� 
����3J�N�����E��.��%�⧰�q�E�߫��-���S�$bo�����G)�١),���Ӂ�M�bz�fe��?_+C�~ѐG^1FR��Y>w;rv1(�B`ڢ��j�ߙ݊6�e�g�{��~{�zTWQ�����*�G������kn�vLicU�?��	���r�zq�~a��4�8��CsX�w:��hR�z�8��u��*%����cg�a�Ȼˈ�D���b:`E�ϓ���*���<k):�g�cA�8I��n<\w��֤V<��Z?r��v�oy2�~wo2�W*�<�ꛩߘ>+��{z|�R �[��;��m��,�c�x��A�7�g�|�)�a�5b��6�p_��;������kPlOT��ln�I�nU<n����������`��ڊ>�ەG�i/�x뤒�/{��b�	�
4�q����
wE
��I�tȦw懟��Г[[0�nk�+^� �=bc��jP�g��wѬ�	���]�H����*6�C�>|;�����������c,��l��f�Оj�)���B5|>�����V������X	�)Po��5�Tb:؋G4~;A�������dc���0r�?��*t�"�ZÛ��c@�Br�vߛJ��{
 K�O��u.2����#ι�7tΘ5�A���$�?�������)�Iy�P#EAv�	����u�;"� ��}'��,*���z��<7�����T�Y��K6K��e�PE�� @��WbZ����� ����
ģv��پfXϰ�v�������ez�j`�B�~Em��{@4�Gc���)�I�u��ZP݇T۬2;vPOy���n�@pUzw@	��̼&��h����Dރ�wv��^�=)�*�w���� W{���h^-���Z'-E�|>�.CZ���瞧�/��她3�<�ł7Jk���5g ��,o�za������`��ʛ:�4������ b�q��/,���@��یi�@�k�$�: ��l��R��~P@�x�Ik�/{�ˡWd=��P�s�5����оy�߾�Kʱ*���}D�e�x�"���e�nO\�{<}m�zOm53q�MQ�i��.~��݄
�-�~�=����1:(���U1-��7J��8� �C�qO�� �0��oJk1(�g�(*߹��˾W��N����!.��a$�c��I�*�n5�BV��3#p���4���"&DT�@�c����q��66Z��>����P4�=��p���@�SF+ƨ��M�L�1��_�ts0�7ԐSEn�B8��?�A@"�wLm�V�ؔ.!��#`��:̝��������}���_��ڃ����.̑ˋ���ĤO�O�r��S��i{��x$Y������>o��ҽ��l���m��uL2�z8.Uc�D�<.L�9�caVg�( OA+�/~���F>�^{c1���3>���Ը��P`��ǫ	]�j6�Ԝ�w��5���ݫss��z0��8M��LT�K�ۿi�߱�r��# :���Ƅ�v���>5�J�R_!��6h�0���h���X��|$��b*	�M��f�/3���6���U<n�F��R���u,I4$t��n�
7Lyԙ�3�"m󤷮H���,��R��@m1�o/U^�,|j>��"8*�
M��hsaǤ�d���pۂ#��/��X�v�9/	v�V�kߣ۽8�h&YC������=��w�M�X������O)�[W�k�����,��s�N�Zw��!B��
/���v�J�e��ƈ�!��%�b�fmJ�j��xE
����7�M�J#�
y�8�c�\:��(�����T8��lM�8
 ���qv���@<�S���8 ��7��7�[�f(d5p������ϧ��o���a>��OAPcZ���`+�P�f/����? .w�ߘu��}�佖�祡h/��g�?}~���q���!�X\���iv�����M{���� �d���k{�����
���
��kl�Р�x ^�WK�#��0�`Q�RM[�@00��0+�$����<:D�d��vlˑ��� �T��@^y��@����i����@^�����Pn�3�.[pS� � س���W�hۏ4T�n�������gp�A:3���(�������d�{����S���ỹ� F�%;��-7w8y^(�yV�����h	� �ΑK����a<��Ǹ� i��&Ĩ�����kl��d��8���_.8P�jY�9�Ϳ���?	hh�����-pa^$@��x PD�aU�]��;�N[��]%���
�tpF̽�y=Bv��A�Ї��w�����v�;��B��u������V<�GZ^='�Y�B���D���6� ��fS��d�1��4���M4��]���g.��9������HE!(b�L ���ߴ#3R$Q��;[���_݋�E ���ƤV%y�k?0�� I[��l����3*b�pkҞ��h2p]N<��ɿ��Y�ҽ��r��j�p/�k�"��"ܲApĀ/ۨ�kSJ9���o�����)[:Y|7�P��B�6   ����?߶�򛰵���E�J%��qb��~B�/Q� #p�4qo��jİ�8�F�1XwOe���z8��w�̳��h^�^�S6y��C�2�
���&+P�Ȟ��K]�.�U�fT��"����0MlCޫS9aX%0df����`���6%�:X�B�lO]�ƅ9uo�">%��T�ȼK������Fm&���S��7��E5�/3��[��:��c�/�`���/��w��L)r.:%�V|�n�����z���������mt�^���L`�	*il�
q�n��Y��nĐ��xc3��J���n��b5
H��'ɛ �Oype���%�,Q�J�X��R������5��6�TÃX2��?�����R	�d3H/�^�S6*1�K|�}h�vԭ�R��c�7~�9���Ak\�n���>{���m�Y¾u��.mB����]LyL˨w\��?�[w��/����v/���`��"�d�ҥ�P�����e����q�?��0̠?�[��E�1�p��@��]��K�w���.t�f�&IoK����g"�+[V��5�����<t�y4�d�3�b�����uK[7~���k��g�2�����:������w�5� ��G����������������_c^3� ��J�y������_��E�ڛ���6��C��%�O|<�oז��r���,�?�aO���6֤�˒]�s�C���4�(�ZG/&���X�:�f���-
3-�R�I�W71���v5j7��਑Þ���C'.�B^m7yl��{�˵?�n���,�����9�ܽ[�s(�ȏ�<�Kcm�I���xfs�~����~Y��;���c����.�E[���(��6���y�3Pcs�#rq���d�0u^�B�����}�����7�T��p���W9��>�P�W#�R��af�o�,� vDxs�waQwi��o�ǎ�m^Ӿ4<�D�{�9�U�N�ouj�sɲ�VR9���ț�6����(K+�e8e��k�7��n�3��BԯJ�����87�x��D@�޳=AAqHG="��ȏ����uQ����D��d"}�^�cs��n��)�:� �%ϴ�:�T�4=�4t5�ƶ��|���|�g��w�nZ4H�s�^�2!��O�<ʑ0�ԭ8��-��iz���mw����^#�;�x��,/}��qm3�����j�!�_jD�߅Eg�SS��jc���jsH�ѹ�Q�X4��b[0��#�?D�&�of��KM]��G1;~���s�~Y�a���
�^>q��;��84v���z6��3��=���59=M�72���h=��j�9B��&~wM��U�K	���ٵ*�g�W��v����V����̬Y|��7�.�vQ�'˄���G֙EJ���?�L͐]��^@�+���;<7��a���E�2��w~"�c%����ˌV׺\P�((��'�r�Z��b�l�߇q���qo�oq%�#��=S��2��v3�J�A�!��*��"��q�k�ʬ��~#���<q6�@ڙ� w�ԁۖ�{h0{Ű���(Y���oRE���;[zyG�z�7�v�d������p�-�:m�҉иk�?U}׌�D@n4!���Tz]+
��H���M�d��u��J�E���p��i�_Z7�9(�9�S���l@���Y�ny&3,�-aZ9����[��p?�y�,v���g��(E�%�?��k�+������|W+!�|x �5�N��'����ŕb��Q��B�.U�]�2�������7�!6D���9W����lH��j��Z9�F*z�85#ńH�(��4��?��ѽV�zJ�k�
۷��*|KU:-�D��B��|��u�m�󙀳 u�,9�9Z0��U��M���R��%�&4� �	ŝ�|�<��*���:�ۼܑIs��p
r(�ĸ�몜�mb�W~f��>�/e���A55�$��¥v�x?Af^�j�Q:lKD�XR���V<ݿ��BP��tQf��a�J�����m���
5�ʖ6��I��BJ�Ⱦ���R�P	�P)ʞ}�[��k�dwqm�~���]���<O��<�{��|���y����o�6�6ba�.9���&����e���0�Z$��3��je;k6�Kl��X�?����55�ܥ�«'��Kf�r,W��N�i���ͷ&��k���L\�����7���ǲP��?y���4�0�D;���y�+�#�����ƫD�:�X����������Y4F�Q�J(��;�j�����M��-��:y��qb�a�H{߿�o$�+�KzM�-QtM��w��n�Ƥ�5��UD}ll�b.�Ո����kRZ��P,�2��L�sơM��U,��D{�� s-�h�;��Y�c�H�"���bQ��;�,��j7�5ʻ�]�w;�/k��wTM�L�s��zl
��t������] �K�S}��_T|��ܓؗ�1�dd���?�=��Mm��ء�T��5�(	�Y�@�i �;S�_ؚ�!CT���Ua��&���°��:���S�h�Yev��J�Vx_Ul��S�!�Ff�vOms���4�ԧ�Ш�9�a��xZ�X�H�s���f����1S�cv��&ʁ���	Ղ�>�Eɬ$b��U1��&w�R|���n�$ߪ����`߄�C�� l��&��V0p��2-f�|A�W3������+Y���J���Ҋ�.5��=<aLq:�v�Z�&u�~`n>�i���Ǆ�NF���XV@}�����j��)R��U�ַ�Z(�r�}�@Ǽ(_�x����)�\�}�6
K�/�:M��p���L[�H�C ��oQ�`N�V��\�᳀/AL���wiX�\��V�W����"L�S@KF[�\ �%"����/xQ�^�$ `~�����L��<M-�HqMUZa�������V��\�k����u}=DQ����~
B���i�A�9�����b��c^�	C��l�VӍ�t��rW�8�~�2���]��d�>k8���]�6#��YHu��t����^���:9c�F�^ڤ _�����hN�Q�uu�h�����¡�R;\�2mc3�F߆���4�yg��H������s��<�,P�����W��*G8�Ԅo�ų���"O*��e����eq��KDԈb~8w�kF1{��;/�X|q�әj
?�����`m�@@0���3�7��3�	�b�����_��������?3x�1����ѻQ@Z�(H&�Kз��M�n��1�����|�L�˃E�8������!'z5ج#~H�w���M)�u7�7C����[�'o�����uFSs_�`jX�d"
��P)񒶷��///@d�Vb
��	ӌV��`�xn\�^�C�<n���t�8�4�N��Y�:�W�Au��ڝ�]�R��)�jX��sFU5ܔ�W��Z@�IĹ�Cq�\o�����qV\�܆z(�9ځZ9��*�c�.G[����`��'��F59�A�Bt�����k����fYi�޹��o ��U~4#-�N䣘�R�͊Z�,�8�HG�P���B�,~�V�*A-�S��و�4Gr��o+�~��v>���%p:���[����~I�VB��y���Ft�F��A�L����#���l������zR&i��+�O�����@\6Х�xO�ʠ�"����pK�6/�0S�r�罺§w2Z��k�n��!N�u�x�W��(�W&�������6��P�t��f��<�����L�����z�<�8�JX�\�[��;���쮓t�s�U�4}L���o�pܿ1��Y���[�FF~�x��4�6.�l�������x����Jt�v�T�p'R�@\��g�@�x��f���z�F��y��A�1���;�j�%c���v~�����{�~�M�YOR��S��Z�	#\�"����rfh�}�hj�i`��oR��6�Eʸ�"1�ҹ[s96���$��OZ~Xx���I+�p��;��V��g �`WT+E�b����^���Fr&VH�*���|$��b�I�~JPw�#e��Rh�\OT\܁��B�11�j|��1s�rWtտ����>@��Hpz9�i���U>��e��dĽ 	NT�fƛN0a�ʵ�j���c�fO_(з:�$F0n�*o!:5!�g�t�%_�[�ZLe�ۥ�c�rϟA}���-�5��/�)��1ȟ�rkc��V?v
��+%�G���H���&��(d� H�F-���[ǜZ+��YX"T ��₳ ���D����!4��K~�LA�3lf��$&n�gd��k��,V`B�������LOv�1�uL/1q~g�V��yP֣�������G�� N�X�Q�c��@K1��+�A�-O�U8Pر����y0`:)~��d��N�>��fe��k���FQ#VyȂ��T�VP��ll]�!���u���#��x�Z�fy�)D����eȮ�a?6Y�r�.4���C�iὂX�R���?���("?�~���S�.G$��o��y���f�5����:3SZ'ԩ��פ�b��6h[�ܶ��3�f��At6��(u�k�� rg�.i��E�t%�ƍ꜑�T.��>�H��s`�)�En��tN��Fu�=4'��8��*��4���\�>��'�y,����F�����Te�y$G$6�=��H!̈́� �˜�൘����e/4���jZ.��˅p�����+T��bўˡPM���N���yw�����
Uq�q�wW��C����ܿ����#�Ν��@���h�񕩪\�D��
��eo\ܙ��Ƣ��

�6�b[Or������I9�6�@�@�����@�"�7Q�y6AVAf�ys�㞹.i>�;`�(�q�ڍRMd\ʀܨ�2�VV�Ke�����SK��{�S�����d		�ƙsx�鴇��-�ɼw
�*z]�}����Ź�a
��kp[��?�Pe2r���Y�
��f/�!�z1��S��PX�Aisb7����?j�z�Ĺ�@�,cCn��׹�������`���Mqǟ|"����f�����2�g��^�s�������b��/��M���8C�- �̯���Seݮ�?���?B�}�_��{��8���  �����6Y��ŭ�Q�5����\� lg��t^��L��$�)�|��:�fj@wVBWd`�g��U�hn��(�R���� .gR%��Q�O��d�~�����`?�ȥ��b��%�tDN�\�dOߞ����ƙ��ȓ�����������:����"%�ڢn��I�'�F�.w䴆_������\�����7�G�#C~��fr�J�:��u�m��{?<e��jG���~�vm[�zltA�X:��j�s�nW�Fr���mɴ#}�ewI�k>�a�ϻ�ϿGn������Ѓ�;��K�^c�I1�G��h
,%�k��\������( �le��\S��ڭ�'X�����&�2��%�FY�br7�|�;���L��v�p�&��#�'��Lk�O�Py����;z4bXd[��̞�����+9w���TJ��'�1���Rp9�:�6��[rw�?��G~�W�W��?Ż!FԀ��R�L�\��Izy*�ea`�)�t�kBN�^69�a��Q�n5m��skc�45�R�n8�ޣ�?�B�3�G	���$:Ɲ��e�Vm��'g�<'�^�>���ѷ���9E]ޢ"�[��ߠ|]	�-sɥ9��$�ǫ��4��3m�R�'F�'�:կ�4dw�|���[���P�)�T�CJ�]���#��[�k�C���9�����	Gth���:�s�Ĳ�����XWԃ<V{����ϣeiN�af�w�\D��������yH�� V钰>�C\��� �Y(�Ny�@�9�XE��3�x m@z���&�"��]�Y0�p�c89�\���Ε�O|�*^�Oy��x�a�l�	���i�S�{A� ��������3o�)#d}�\�r��#�Ȭm�W�vPf3�A�	��0\�G�������Ƈˡ����Y��S��n�_��[�d�jy`u�s��3SN4�y�Z`��R]a����|���xJD�{R�/���1/�*`�1�����lk���5�yxo%�tU�� �S������3��FHص���h� c'y��������ӌ=MPl�;i�5V8)�#|�"�떳���{h��;�v��bg���� t��,�K�B���ˌK�Z�R���܇%��Ʌ�:��M�U��&�!�"���ܐ���U���_.�--T���ڙ��,�������/|A�kתr���l���>�����̛�S|���©"&�(�:�xK��D��iHH���R��n��a�=]�����_>��j�����>,����U��|�{���x���O����t�:ک�\����	{���� ��>c-E�qc��}�������KߊƇ������IqI��V��V�s�2���߸�s��Fw���jIMߏ�s�Cj��������*�[K�[Ϗ\��+We����~�ii?�,^�s�БQ*����`y��i��|���k�v�C�iw��3�o����:7�Td��q���5��}L�.A%���<��\��������:�˻17�=��A�(���"APuߠ�����4@N��UQذf��f��S]6�y_S�a���"9J]��Sk��*\�Ȧ�WO3�awid�hR)���L����t���Ɖљ��<���������B�!19�L���ʬA'/�cx�{���j^{{�!a����
볖�)#����W�Nc_�R�W���a�A:b�̐oκ�k���A���[ŘR�`��s��l�֢��"�q��Xg,� "�-�,�&�e�2P̡�o���8�9K�e-������ľ>� dЌ��]z�5��ؐ��!�7��\ʫ
�0q�[^|ѻ@$��}+�ڧI�;'�A'�O)F<����_�~�T4_)E��M��>~���0l�L_��pu��9C~�����Gy���\����ƭ{X+ٔX�@���K��,��Wb;a9W�NhK����*���'�;b�2&��_R�.'ks2r�56�˫�;�5#��G~w�֡6�B2������x�
�ƒW�=�b7�ڽ�J[�5H���&���(5����>?�4Vh����{rO��d5I-K[��ܟֲM�7������YS�A�Aw�+
o�֚j�na���{|��}�6�0���&��d�d��q���CaQ�~��Q	Uf��4D���{vŠ o�1�'
i&�.cQ��n��t�o�ʉ�O���(���ɫ�63�4*/����~�f��%bS�J�Hj��{4��v�Q������T��C�Z����Vz��0��-��P{�֥�%����y�*���j����ZOk��~����jk�А�ֈj�(@���xv���H�"�ܙ �=��)"_1�,���q�ڼ[�|kA�\c��]�˃��_����;*�z06zȓ��<����WŶ� �Q��3q��$�r�M'Yo�VQk7�zSsF������\�'̗`����_M:RY������n|s��W1Nt]��4�K �)�i�*������'V�#x�b:P��������	M���P-;|�|�j���lF#�>��}�N��iY��%+�/bpsG���w��i���d^�v���Y��	Z*Nr��~<��D�^5|�e���P��'XN�[w�{�>g���jp�*�DG&*�N��!�����z��	T\vm����c׭ڼ��|�� �zR��0��I�`6�y·1�����3���Ip��7��`
���q����~���r�����X5�g��9k�ņ���o>]�Ҫ1�3��gY�n�"�19��6��F��*'�_�>oR��%�K?�yY\Ԭ̝i8Ծ�OcP���}�W��m#������|����T�����Y�R����wc|j���zF%�J��;NNUe	<��L_�$l-�a�iy.T�H��Խ�N��]z(!y,]�1�WeP��pV��>ڕT�١�HG�hܦ]
�nƒ`�	t�\/�,�)��l��W����%E�c)�E��h\S�k�a���̛��Z��Z�xd3�P�mq���Nr��Nc�A�c˱�,�VJW���9w��@ޤJ+�]j�Y~�R�㢟��C��9(�!I�_<å��p��3+ߣ�!���q�H*Z��jM	�h0g�%"*�(͉�$R�s�V��{#^��^N��G�r��~�\��3b?ΨKw���HmH~u��U���5�5�O.r�]������,E⨜��g�,�%�!�ʺ'�+�pn�×h�D�w,PںI��<���H|c�%[3J�|;�����\gnR	vJ����V�H
�6#þ��GoU����"\'���S��z"���q�<܋��T8���`�EzHQn6�:&��C�͖lǆ��O��ݪ�����y�l���W�-�޲�دrq����?Bf�0���S?��P��9�tD�8�}��%���q�s9j�dɃ�[�X�������P݄��.�D��EYM;��3��ѽ8���#�����Y�PJT{�x3�+v7JJ�����;��5���g�4����a~���%=@朗,u�w����1�MWŮ���ѕj	��
ot�>
eDޠ��>���-�����\i�}X�hWoIR����4�H��L㋏�Pa��3�r���7y�0�G������2���#%�����*�3��ɪ,�n�H>��[���1���El���������R��Xy��":n���oo�wN�\����[�?E�xO�ڛ�-�פ�W�D�MԟmQy�3pf�>/�l�A�x�g(�cz6}�2��t�CQ�� ��VE/��D$��dGN.��z3b��Y֒V�Y/�?�����Q�t'���Q2�\�
戤/�x�'�E����;��q��G���1.���9C�Zu܃,�W#��䯏wU�w�����mZ�
�be���O�i��{�&k�\�9hK��y�S�X�&����8)�<!�/h��x:���#V���nbuZd��|
N�E�8�u�N��ب@�xs��G5�Q��{/�b���r+"��;����8`�\�M���'����4E��hSo��o��{9>�-@�x�P̳��1�S�^2i��,'�[0e9O��cյ��ɾ�T�݁��(�-�����4p����5¬�nH�䙗F�e\�Ëw��Ji��������3�u�&[z.�VX|�m�;2�pN��&bH=�)�}�^������5Jj��2S�ac^��Ɩ>���?	g��C3�A{�5�)=�F�5Cب&��V������D�L9��k��4��=<Y��Ҵ�)G��)u x��ވ��>��.C�L��!�4b��7�Du+-� �������(�<^�h���wu��?e�v:��|����v��>S܅~�O�7����/ѕ|ƺ�;���L,w�z�M���D{��]Z�i.�J͡�������x�}E�Bk4;G��ڏ�ʁ_@��'�4sRyNM�u/�2hAـ�[���e�Zλ���}l�e0W�nc�WY�@ [�9)7\ɜ���ʊ��K�ca0C�E3$8)g�Kb�K�$�h=]n�=(�<�1~$�u���}5����u�ʽ�BAW�t�8[*�k��I�ً�Y�����R��rƸqo�s��ƌ�.l��KP��KާB�����^UCN�E�)�rhE�u~������TM;�`Ne$��>*2 ��k.E�E�8Xd>�7��ZaS_�M�ٿw"�B)M���k?HL�yW ��*�5��D�L�|l&���N"Pj.M5���2�X;���y��M��Y���Hޑ���c���j!�Ŋ6	�2;Fms����RA���<$�/>���r��ċ��H�r��dXT#���+2�9&�+~�c�0RJu+(sX������a���J������O^��n�W9�l���ف��w�_�tA��Tn��_�m�x������#���>��[���y�i�v�Gh�+u[�>V"r���4(���q5IMVYs�%b��`Y��r�;vX>���V��dx��`K<��k쟟S�s�Wþ�3� �Hf@O��Vw��U�-:����)�=���c@?��Ar����n���f�pN���]	��M�cfr'ܮ_3�5-�U;�;��G�2n�Ug^��䶴�/	KX6D4��_p2�s�C���H�J1�����y+��I��~�H�ے_Uu��*D }柿	�C�w�� c�̜A϶b:4("a�{haU��B�C��ϵە�h��:+���;��@FB�����G���]�a�(�����vҼ׊F������?�Y����ӥ;��ɍtNZIN	���#S�C�V)�B�O|6֏���E��U}�'�rx��ǞO�Q�;��u`]�zvu�E�p-��������;V�׊nbM}@S9j�,#��V��Y��:vGMџK#}3��b쐨D��b�u� �ʣ�!�l��w(v
^��QH�����=yKV�� \�I���Q�� 	,��I�7SX�Kg��n��Qуd�����R.=�V&�u�:	9}+����!_6\Q�cݘ�O�Z�����b#��b}�\n��t��L�帋>5�ƴ��p!�5��*��䰺#�T��`�2�<�b����1�s�-|v2�6ND?g
/6��"�h+O���e��˒��ZQ���-3?�9j�ʑa����1���G[�`�m%M����X��=�s�nNy�����v[��z[��*��T�����lE�T~��;�KP��%r~}��%t
 䃆��!n`���Vڤ��r�י���; ����ٲ����-N�F�\s�I� !D���;�'�0���W��$�6�vG���
��I��P������+�o&����N~؉Uў�?
'�,&��V
!xՔ�'\�dU���X���XƱ��� d�6֠�X*�E;1�R�[R��ȹ�g��f�![���]�D�����εl¿�1�x�X|NQ���꟧��-M�!>L�?�|?2\��G���L��k�f����;~ћ�K�I������^e-$nWv��m�鶵q_�P�����'e�<�I�.;eǎ�-{C�܋H-����e[�-�Y?�	��v��su�����ׯ����Mc//�䱗32�D�>]��á1�h����H����G�b��5X�3,Y�=X�/����Q�Kf�0ӭ��e����W"��z�ܟ���Ũ�I��p�����1�t&j)��^��E�(^����ެ=w�G�=�i*��R��-��E��}���G)-G��l�B���<6�x�����~U8��C�pv����S�K����`������--1�.�K��1�gPfa�V�����53= 7H����)vO�sd��I]l�k���k5�s�%�w�t9�B���Y�[��l1����ɞk��ac��^n�A����7h�blV�/���b�V�?��>2\8�]��Q	Z�s�Myj�ި���b�D�5�Ǘ�����n1����$9/�q-��w^z���Arx�����ݳ��Z��	Q���R�q�z�"Ӹ���h�HwU�E�?=Ό�;{����K��:Wáq��F�L~ɒڥJm#�����s��|����࿨r�ԝ�e���
1��z�uQ��{n
m��,{�fyF�d�r���1�0?�����]��EX0O]��{K�x�ci_)�⺱���k�,f7d$Jԭ�����g�J�D��&K��nرn��8G�Q�M�u�>�2� ��S�e��ײ��X��]�:�?,F���N�/H�xL,i�١��i��ҽ��L�53��]�бīt��T֐�����̏~U�Ut�������=��}�{g�p"M�t1�D1��W]_�?Q��O�/�R���L�nmٕt�p�*�Rf�JT,���� !��e�0����e����cӺ^m�3+���?me�*��+N���? �e�1S]#c���ެ]���d�K���Xb�Y�^�oWr�x��쾞zeކ�����`��R�j�����e��J��i"�T�v+���%�-K��OmȬ���q��䑒�-J�����ǘ#y��ړ�9(���a�Up��.G�L�.��h7X<C&���11z�މ�߇e��?\�^|�l�Ē�,�%.���G�\�X>�l���1�ǃ�ڄ�>C�G�6�z|��hG��<���_��U���e���B��dk�B)���YY;����VpEO�:ñk+�[����FO��'D�<�wk�"��]�ٟ�1@L߇n�̜��qv�p�55�@�Gߓ�	aPKC]̊�3l�Y~�o�3^o��T�ڔ~I�T~lm��T����xM]Y�d3��w���n��.l���/���8vo�o��)�~q���"
O�6�=�h��|������Q��ީ-�i��p���zv������F���npa�Д��%����w�����-G8��BT�1rz)�@6^����՜T, h�u�*R.��ͯ����A�i�n� ���.}���6��;�dY��4d%Ir��7����t�/�]f�����z���-��?�|��z�2y.��wh�]ea�"]䬭�����$�I���c��ĳ��ʭ���u�7U����1f��W�V�x�DA�Vo�,ߝf����O��7c�뼄��o<�=O�;�\��K�>I���A#!a9��SC֮��ȇ�����tؼ��EP��
��nj�+;R����H^ogo|�4�A��x�ɬ��R�&_Z�쫳��������H�}a�ʚR��"�t�ȇ~ZG]E�ԟ	K�����s�ȑ��"�Y*�[\�UHF�"X���j���A�R�,X��3�q���*ƒ�p���U*E�y^�$੩�A;�s�;Ѯ~h�y7j��� S3!6s�
��M}�c��Qʺ/݌|p"���fT+����9<&@��*�Ƣi�l��`�w7Z�(�C�{Gl^����H�%��c�>{�׎)'��!Ə��N:%�s�;W��63}|f 8y$�F��X�%i��m�j�xo��+MG]N;N�eo���Q�����!x������ʦoK��ܡ =%��a���;:��ۿut�������'��q{��;����*(�:t�W俘��q>�??g��h�=?�&c�P�$�w�,�Y�S�Te�zr�*ƥEa�8��}*���u`�m�I=�g�n=�1��p�OW������k3���O�#f`.R��h���n��紼�L��>M��|Zs�nތ�%�����57��c4�R^ 3��9
���37��oEmL�!�^�(�tQ���!�E�#
$���]w���N��V/z���,~-��j�� ���ͣ� g�͔̈qD�nQ����á�Mj���j@�.{�EL@mм!�1EY�MS&"G5�����85���tՋ�¨I�	
�پ/�o����9YǴ�r��5�{U��>�H����1v�-('���o�aKs�`��`�E��r���m���t���[��ln��)��nW�#c�Ò�Egѵp{�ô��ؒ�-��zܢ��'@O+�Ǐ�����TmEAe���n�L����w�>��s�����G�\!t������>�!��ѓAU"���[f�*�Kq4���1M���,J(o#���E���eǦ�)�8O+g�G�OSs��Oj�,iG��x��ސ���૟֓de�OY��>dc�2�bÕn�U�tȊ�Y?����8!��>M2�_����K^�{����I����Ȥ�FW9Էױ!C4ҷ�,u84��u)���}�[
6a���{��vq�����)əmb��}��r�ec�HQÖ����&�ǅ�|�4X�:]�"��p����i�<��U���lA4��p�Jb���2IE�
wT}�N�(NcmgP�Y���o�(0��0�Ø�|岥�=�=�|��=2�xf���{:�����C݉�g��RM����yG㝨ޅ��ɼ,�~8��	����9A���"��ݼ�@L�!���˝�}�}̑���hɼ�	�`g/Q�+�0�N�<��Q��m���{�|4j�
���l<ґ�!�yd�>�_xR�۞����,�,Ag������&HB6��V����IGbo��gz�l��� UXp�V 丹��cp`4�E�͋�
>����`��5���6���<��>@�@�L��
��[/$�l�Ó$�5l����䵠�[�,�3� 뙷n񖎋����C^�4u5ZR6*�����?�B�@ �.���_����H����N��w羨�bb����K���O.^8�����p#F�]�J���""�P��꬗�Q��Bv|��1(j�R�dM����!�\����&��|�H1I��X�ՆЙQ���K�
m�L��`��Q��V*��0���K0��Dex�XCM4E��r���J2��n�{��K����1[Ϳ��哆��M���b،f#�6"9��.�Ab3�K[b�d>�?uG�=6��:����Э��v�U����NI˶� O�ݱr>�O�f8y[�ЀL���c��T5�g�W�Xo���[p'� ���&��r|8e��,�߱�� J���Z�j\Q<@d�8����ӷ��"�߰����h��j���Jl��˘��}V��S��8�`vRu�L"f��_� %d�%Ǘ�+�[��r�����?;:��4GE�:'��_����O3��ġ�	�\`��[a�ۖ�R��� ����u���&�0ҁadpI�WZ��VڣfM��d �䥰����I	��mx�1/�����G=�"jp��`� ���Qu��U�W��)f�����а��ݻ��5W�A����ڪ(��C��+���4|b���TϞ@'��$�`X]
��--ݝhg�v�����VS�IW�Z�w���V�:�ڋ��}
b��	a�Ӿ��.\�I�q�t�`?l 7|�&n{��U~QF��*���&[�,r������=��]Wj ksw��`�y�a��3�9�b;Yf;� ���O�	���1��W{F) �g2m�� Lm`m(�ci�=z����Uzz��<��?��䄚�Q�s�B��,���n馘�{./��[l���u�є���d/�KN+�46��jW�*6�rM�^���x�5z�bG|{�����`ׇ9aǜ�G]��Ū�Y}�.��6#�VSo�� �#��M��r�I;}A=�Q��0v����I([�����A�k�hVD���]��1{k���M�:}����lR�y���AA�u��=�H�����,(b�̺ӊ�r͞6G�(����A]�o7�n�b̺�e_�5�7�I���;��#��!�-Q�ަ������(�{�6C~��m���XdS�\*�	ˏ�(L���_Rs�\@}��`X7e�/��Z�p�yшF	T�HП�d0!Wk��q��P���! ��M�����	Eb�57E�����f�[X1j������&�PY�{ڰT��Su�䞇N�c0��6��>��l�f���L��a��@����N�#{�v��[!8���*�;�DΕ4�hU�E|�C�T2ѻ4V7�=��°�Ǝ�)S�d��G�GЄ�Xs
\mƭz�%I���g7�~9�܉O���-	`>����h�	��:+1Ú�@R��I Q~��?�~Is��e���;�ݥU\��9��F�A���E^�.�W�$�[�¿��2r~�J�;�?�:!��	A������&G�Qx�EIZ.)���`/&خa��YE�r���&���eW�7 .�� p�� �@�t2�n�fy��+e�«;
u7��$aW��p���BMzo�K]����g��T"�P(v~�z0Mw'��l��o�!�X�;~"\;�N=)�+)�#�s���2��<�*!����Y��f����T�!04�{J�`,i�����B'��uL�@���~f�L!��&Ͷ{x]����-Zs`���l+�
9X^��5�\��$���?�Qo/
�] �q%WuM����~eG�^�f��U�T��qƑ2%w�ى�J��tw.�ůK�]�#E�-�c3/�E���9U��̫�L������|��"P���B����ECڜ�#�N**�l�T{M�D �"�U��j��m�$::���~�NA��ċƨ��g_^�|�\��Rۿ��9��#�2Z	!��^M/Q�Q#��dz��n��f��� �%�)Pv�F�Xj��d�O�b;c+��0�ՠ��ler�ho��*����#S/`����C<KG��Xg�`�#��ЮW^Z~��=��6Z��{���Ŷ��2W`ji�ԵLWյ���(.��ۘ���h�`^�׎�~��7߉��\�"&Ѕ��׀���x5���WM�ךLAޡO�[�[E�/[�cjV�.Bf�6Zp5-T�̔�""���w��8�Z�E��a|�*t���v%�|�v��I��z�
�،�'�*�EO#�<��78���{�Vr��7t@�F�\`�Z�_TE0@�i��w��/�
��B���2&|a��ŧ����W(�NY6;µ�R�a�8��('�#a��ՂH���� rd�$�2�m`�E!��r�%�6�})�|_��;�
��'�[�#�!d�~��R��\C8ƺ*�~��`߹~��6��W�
r��&�;�Ծ�\w����/�g|����K�ĳ���~��t�ɉV���/��=����@q����v�������i3�w[�o��-M����5-h_����3:���p̴����i��ϥv�XT'� �h?��x���W���p�k7Z�I��4lc!�X��x3%�-��Q�Հ`�F���������@��_����l��By�]i�a�=iF���,�h[�*�D|#,��y����̍?���dV�ykߍ�	6��b8���A�?7Zl��$C�������>8]�g`��}4~�}V�R�K@{�k�TT�?77Є �6�fʲl�.�@mxSr�Q�xIL�Ƅ��M'�/}�r����X��r��iR'C�6R�sP;�aÇ�>� �0�{��P;� X���&8�E �F�n2�蒱��:L��@��u��Ƭ�:��������v�?������F�`�N��)�f�<N�)[5(��ϟQ�~	�"�f�(�V�-�!�۲�c�+Ńl�M
n��➻�taq�P	Ƿ�@C%�moڠ�t��U
R޵�.��{�t��&V��;�G=���n��Kͣ,i�k�YIM�'s���R�{A�V�k�H�T��~r���&T��"���%0̴ ϥ�zݫ���x&b�碦v��~�Y$Q}4�v@�q��ǃ�-o�����<�P]��ź�`'k]���A�!��D+�]x[������;<����OM�'�3c��ı����Cs��h����ǟܹ7XȓrX2	��,���%� .*�q8����� :uO����0R,�;�����LN�6�OpĶ����>��2��˝�tKf�:Bg��{��J�T?͉�Q������S������0���C4�
�Cc�7�y	��#�{Ba����/��x��+���k�Fy/i�`����y�DE�A�1+�mBG�������+�|��H�R��-w��.�u��?���B�YD�/�S��ʜ��L�{^����3T�?�/�.GI4wd���ೲ2HB���4�/�ލ�����%Y��Gɀ��2x��7T�Zi�s�p(�A*M��0
�n1<5"�㴥q�� ��)1��]>{��$ġ��5���o ��<d�?ZD�z�aDz�i=�6���?R���4�Z7�`R�z�z��:-"����}p�3
�������i%xe�E8�A��/6Σ�-�_�������ǟ!˟ݩ:�l��Ʒ�]�N�ѭ��\[UN-���
H�W���_��֟Ӱ��K�`��0n;��k	��oCT���X&��[=.�<��������$�zal둂-�^�
3�2�mē����O��a�v�T�ኘ���v�?^���o%`j{��Q;�r~!X����MҚ�!^��x_��A��m�?��~���-�p�3����N��)���C5�I����-����a2m���_J_�v�m��p_����K^����͟;���Rλ��T��ol�uc���S�ߔl/��V���'%�cMsCu5�.Q�3�W��$Q�8S������մ}��T����߆Ҍ����y9������=�7=�n�*>�lC��6�۸�6;��;���-��޷�bY6���Uߖ���H����0�'4��#�W4�R��r�f'�_6x�����t͍4���E�zd&�zتɼ�WB�G��}C���Ux{��K���9��V�#i	�3�
�=�YV����َ�$�{�3�-���
g�kG�o���Ic���	��&�8�g�����xF��R�2d�˦���XW>v�?S����TZb ʟ5��q?��m&x)Ӎ��9�Yκ�E��Mv��7�+�� GP�܎x����ʫ�cw�.�2��&�7��+�g�<�h'm�w�8Qb�S�ė�g��(��p4���zd�a����=O�f�C��L̙f:/$U6���������D��_��O�zw���
��H�9�>�'.��Ĩ�A]�y؍ʕ�|��ɒ�Z[��(|{������ξ�����#�ʡ~��[�g��K�ۚT�t;�eKY)f��yN�}�c�B�?��2��K0o~D�y���Ҏ��-�z&kx�"�2�o(�n�$��ܻy��=Lz��w�??Q�U�~�j��[�E������-���f]x)�}Ӗ����@������'"2�û�4�3�����XbO���[ҭ�\HԽ.Xm�}��07���T�~��k>\0�����?[ұ��<���*9f��L�ts6O��<W���~~�e5�M�L�0'�'��ue_�m±'���{�+�FZm��\]i $�6e��x��sgG��58���g>�� �^��w��>�
F�����b�0]��:�:�:�O��ι���Bp��֙���@e��f��Χj+ l��g��,�	�q��)<Q�#}Z4 b�K�2���nb�r�gs<[���������3Y'�-�*�pG3W���=�7���`C7wu���\X�YR��e��$��p器ù�&):�8�iQ�&������z1���k�	�ҕO��t?��� �[Q���m��������=���E���:z;jEe8����[/�G2��,D���7=��q�rp����l k���U��d(p<V�������ժb��X�C�\�i��B�KiGfs�C��@<^��bϒ��7|(bS�zq��UE��k��@�8�Ù1g��<� �ZyU_�V�V����P��b�zp�����h·���n[�M���)����$�qbh�r�y���DW�G�N��u��N:|����4TK3AP�dxV�GQ
v8C_9~���a�L+��N@%)�%<}��%�ֆ�5�yBz�wo�[y�IEa��4c0]����v{!��ldĸG�7"�lL��i�Е�����8�ȉ��6�m�� ��J8�>��')n�%�����r�c�:b��<�^�}�R�#]�ie�I��HGIԽ�� ��+��	w<�,|L#�[=��������K�S�L�S��qEd��7��ᛧ	���gx����1�Q`�u&�Vփ�I?GͿ�2�}��7:	�"A����h��BH���A_�<g�ee���>������;�(К	b���1�p���XKn[�F�S�{���_�?z���8V���H�zQB�;�� }hf��{x�t�鵛C�{:[;��@��Ղ�)=�G�#
e�'�{ծn�=�;�d����pt�'��>���l�8�4�p0Eܜ�b�c�����g�/����eY�g�����wW}�Y��]��;A���C� ��˧.�.wJt銔u�T��2��B`�����؟���k{�ڢ�ޥَ������eVb�w�����)�/�O�5��?�z�"�W������{	��=���?�x�1��(��TZJ�V7�v���M�O������K�i�rs�9�m�>	�̟�����&���S:	)�e�I
��iяmeO�Μ�><�'u��ڊ�=�Y������r�F� ^�*������>P[b��2�
�<F�'R*��C��s~t؊Z�&'������Vҥb~� ����9s�#x'�_����\�-��@\�W�k��9�D��j@G��VkĐЋ��~�Y��v�����6-��8o�����Ȟ8��	m�Ԗ��_�0"-O7/�}��6�g�"�4b/]�0>q.�RT��D��ƿa/J<�vQm��%�<�g B���������GB��ľ�ס�]q��������g��eM]�v���~:r��{Yw��4/I6�^�z�g~!�W��[�w��`��>����r�Y�z������>��p��1�'M��eyʊƶ�A2���R_����_	��P|�S��љ�C"��R�B��$�3���\��ů3�.N�=|�T+FAd�B�6Xj<c�����5����{g��D���@�K�mpeM�g��W�< _�+�JT�u����/���lbn�m����}���n����g�m�����w����)���i���"��B'�Nԫ����WY|P�'�i��'t���w�sp�bh*�,�2h&��n�$4��=�ljm��( "es����^�]ׇx٨9� �/: �q�#�?I��f9]���ȎK�%��",�A�d�5qH���/�E"�E3`�]�)k:k
��l<q�ϫ����.�,,M�{��6B��#�yl���>�M�>�*�HG��ͷ�͑v�d
�/4���ׅ}C©O)��R���/h��/��^P�Y����f�W��F`�$�z1�:b�ˤ�s�ٿ���VÒ�9��b��k���_;���ہ*�
���*\*q��uRz$ބ��:�6_�}W�f���f�g��:�g��I7��{	E�Űj�ֹ��g"2����!ߜ�Q����k����S���	{�菸�����~�|�<�u���r1Č������Q|�7?������Ū]���m��3bg����-���9�lBBa�������=�ePq&A�߆1@�FPG�[�G��&|9�J?�&(2�h;�/�����޵�hO�f(���������G�&i����A�>�OD�+QVd\+�q�T�L�%{fo��yCƥ2B�#��<�9���_�y�����~���sι[{�i�7l�R���m6V���Ϝ������ąH=磨����T�c8G�A�X��LcsS��Sr��1��{���Dt�A,��u]k�ZW���;a�ᔃ߫��˘ā�T�?0K��$�������ˊWeL!�@b�u����T|���хI����1��ar탯{J�B��+����H����Y͙t���h�U	�oŨV�*�0��YM
����S˥Bw`��~�-4PUq]z�@)�7s�S`�p!�,c�Ѩ�c=�+�y��P��Wa���i�@lxj>��)ej�}x�7hQ�lNP��qQ��R��y�%�Tp��Nvs�m���bV@�i�<U�L�][O�'J�RM�����),��5ǅA9��*���ٚ�>U^5�����O�I,�5A�����1�#F�����n���:�@�t�tIfF����31;�9�0M�_�:,Z��v�n��_ �wHXn��	Y�%�0e4�-gݖ��4�A�ᾆ�ؤ�M�9��dr�w�����}��-򺹽�s���{`���V�7ּ:�l~J%:�C�4��bkdf���ݜ.���s�u6LH
��`���[�J�/�<J��Q�ĝt���ts�{��t'$�tF�ӛ'/ɢ�v����~")�:���� ��j�)@YʵoC-������~]硍�!���~k�	-��\��yBi�� �i��N�k�d�@�d�����Zݑ�0�4�Hb�zOt�͕GY(c�e�SML�I����K[���{m|�ۀ(n+F�`�Ԅ��H=�*���b��3�
ܧ{����֧WA���e.�I�ra��p_��i�s=���"Ƙ��&�N���`� ��.���n\��ӹp�kQ���e3R��~�8�df���mo�Yi��YC���垐#e,/o~s`�� ��+f]������	�h�?����!��\S�����<�y�^�=�n�ӑUo4k��D�)���S܎�Ro��oH/�7��~�������[��W��u`�R��~f���k40�ţ&���I��j/���ANB�٘��R�e�~	m5��^���:���r��0xx�^�-DS��	�ۥ�%i]�y����9������Gz|��RX�&������i'Q�׾�Y]g�V9�H\�6ZB:�^���֛J������t��ц3��ym��/���,0���fG�����J[�j�����1��Fg�l�=���)U-dQ3�A� ^K�#�� =�mU4_Q���Q*Q}o�kc�,Q,���R�}y&T���|�Y��G?)�n�j���%c�mW�}�����Y�?�'����L前Oe�G�"6�a����H{|���^]z�I���XK�v��9�f�t�Y�o ]��_D��������\����9�F�U0!�`2���V��_�������.3��Ҡ��C���G�^����ځ������F��+)��Y�<0 �,�5�W#x�з1
R�i3��/��W-N@NB���(m"ngH��rn5����tτN�.vƶ����s^0�7�W�d�Z���x��I�[�@�"�1�qm#�d-b�az~��=I&$6����1�{�'�s�dx|����T7|!~���T���{��}�dK�J���c�� q"������cd�[�!]57jt蓠�n(X]�ˉ��ل��t�������U$7YH����*(~(�Y�,���a�8�>��މB\X|�:F���K��zbQ���_s%5� �ԁ�|�2��Z�#e�O�j�D3�9'�j�[�|`�Vy�]����ϔ_��5�"�IVob��`'��&b�|�eE�^Ԯ�瘝D㼄n�s�/|L������z������� ��a��
�4KIa��3�0��q���9���m�:�6��~��K	}��ʒ���{#X	+;��R�@h�ϓɂ�{���o��2˗s<��t��_023��O�৞�9���(�ҜSP	 �G)Vq��	HE�ޔ �����{��6�Y������{�d��y��g�缌�򯙭 ��5K.�#L�.
Wd��D��XZçf�]���̕��Bpy]%�YQ�"Kg��b.���L�u�nΎ-]!SU](��!5�i�\��+�/��Z��FN�ʌ�`��n©�|�3'V@��y��m�G����밆螀�f�����Ƣ��5 %K����)U`ԋ��2QԢ��PTk��Fa-����f�I�=���#P5�O�"�ܘ�?��Z��j����Dtn�d�!gv�$����� �F�AC���.-��6o- sM�*���\ݚ�X�l�c�����)+�f�F���)b"����>�e����K���v��H"`kC�����57~���&�r�B�Y-H��0�Oί��l(º�?:I�$��V�[D�iL��]�zK_��m~`�T9�%VW�/|�XNx0,%�Jb����^��Wd	ء��f��m;����?�"��|ZU��R���'����\>bk�uQ ���)+R�"�:��]���?�@���.
�]�L�$�X���[/�����FK'�pn�����I4\�N�k��9W.��K����`�j�2N�̩��-�Rւl����N�I-为�ǁ����̸����V� L�ꀔJ^t58�D,;�9HY}b�R��9�=[c������N�so�ZC�&��-@w��,QC$f4a�;��&A�m%!��nW�L�m�Y��~�<3}`k$����L��S�}��|gS6�����K�R@Z�D]<<�\H�y׮]v0_�m�U�P� `R�BƄQ���?��'1jm���#2n�@����@�_��<�=����!�����"�/�u�$&x����SV�,J�=��
*j�;mF����BL$«�;�J"v�n���S�����1�h�1��r{��0��AII��-�,���Yz=/��W�-�,��;,�f�*�Ԧp����[�c\��Ȝ ٩b�T"� N��8��p����!�s���~iC"����f���&%��m����R�O�_�5~��_,%o~3��Et��6s&�mY
�L�#bn��ρ�O+]��Z�8�)���};��6���f�)��H���/x#��;9:8Ǟ2���E�I�����ր��?��%�E�?�[��>P{��/��W�R��,��'�F���zg�����5��~��$E�#;��9��΋��Mw@x'v�������ѳ�u�R�~s훫hG��U�ag7�x�c	�:b�]�i�_��}'2�\���P�`��O������.]E�XW��wߡ����HE`�!�ѱXvw{��~���k��w@
�,U� ����_��$f�ӆ_&&���ݠ�A/���M�����"�rY���[�R�	�6z0�{b��,��"I�Q�"�7�ՈҘ�_	Ŧ�/E@����O��5 '�����U
��c��k�Șk�����$��W@H�m!��qN8��ߐ�km_N�r�(� ���5�C4|ڔT9X�h�5o��{�C����ah�p�F�F�L�?w�����	����ŵ�C��d:��	,܆��+_�nm��깱EsWen�a#2{�o�.#sb��%V;Y��B�:?)p���{݆?T�/~�:ǋ9��;^3q߶2j�ۤ��G��XA=��y2�p�E$3���ύk��|W?�����gYP��;� �%P���G힢�6�_���+�&K�%�����5l�Q����{�E+/���9l���.�\��̂a��1<�6;פ������PN���+'�YPW�Ɵ��Qd]�=��W�A��^K���"2`uI �J�A>�p�JW�%����c��̍�W�#�nJ:ǶY@�l���>���*Zl���� k�w��2�n�/p^�x�Ri{�5}��0xx�F�`�N�
��c�����5"�F�ɐ���P��^�>�-����Iλ
H=Ǌ�7D�� n��:��ZlP3I:18���m�V�ѱ�X�I�o��W�	{�1x��nO�4ex�_�Z�����2D�@� /��h�2er~�@[ 2���e�J&���B tc��	+���uz�P�-]6��;tx�ى�SGP���k��Wt�sｺ��>�ނ�g�{8Pk��+5�y�jS�̋e�v�tb@�W<��Nh�<4]�L��
7H�+Y�AN ��,�i��+�t�4�1�Uv(���u��Oy��{��LXk�4L����d�>�%��*��P�z�b`��1_������u�_�y��������K$�����n��A%��<��r��tJ��L}�OH	�~1>`�>�	�+2Y�131zs�\bzN@��cL?�a�b������3�*WU7�8�*�o's�A5V3�>�s���q��?����M'�V���a�|m�gP4��K�~h�a2���>`?^@��
�B��tG��?�"�d�v�_l�;9�MO���N�ى�)������Ȱ9 {x������,zk|(��u�b��/�7��4d6�aܻZ(����<~lML8'!�C��y���nY��$�B�Ha�V�����^j��`n��&�3�s�}ß<��g��<��ˈ�	j�X�*}�"�
��@"��a��f���Q�/-�uqX���z��D`����kxACI,�����F8q(z̝x,�2(T$J�i=h6
ڜ�kuZ�ֆ)�85_7닢�֨����94��L4���
kQ��
����(Ӳ'/;ޛR6����E ��	S�:���;U��uA6^{$qn3Lt�� G��8���g��+�k+����W�w������܃�� �Y�IHQ/7�G�7�؏8�	YU�@�ߕ؋d9�g}�5�:3*ք;R[�D�u���꿜."]�����KA'����ϨX���ª52���%��Y3����4h<B�' hڸ'�3-]&�lA�u��X����z��<���%�TU�W��:n:�H����ǔ׬υ.*����'}��9H=��#�qĘ�#233�y��[���������o���5�x���
�nBc�n3��I�����׊�h���hS�c�W��-�a ����'W~ͦ1n8�%3}��S
�G�t�K}%>�^`3�B����&-��X�%� |���c�G,G���h�~�<R�Q��M�\Q��K^?o�K~*���N�Y�Փ�����2�9�?�3`��c�iG��_|q���e�A7�7����5��t������k�>߿�}+���G�=cd�qf�ɕ�~~�r0���b�	������t��#OZ��X8��{۵;{�sZ����yET\t~����*�ZX=.�~B�KiW��Dg\��/�� *$���I�1�aT�(�Eo��G�3�X���F��ײEU�3�o�um�o���X1Z�~}<x�F����7��c�5З;L��^���0گ��E�~����C�z�E�{*����[K5�uE	
�co88��'�p�rq��KF+SY����?I��w�~1�V 8�v	���åaF�E�7Kf���]���{(ģx�ڎ�����x&пbG����XY뢢J�S�4i���ג�tǱT�Vj�h�^��BU��L�~@�Z�or|�y��@�z IAܒ�x���>��y!K��1�clF��am$O�ۮ�u�.Q!�U�l���F��R��kh��� !�t���r!���4�
���^$P�ds��P�u;�9��_�pA��>)���~b_��C�@o�O��P�[�Eo�VhK���<�5������_��G���nɤ��{��̡Rz�u��f0�8�RD�S 5{�:53{&���m�2�F�{���,��i��-t*v.ǯ�
E�Tu�Uk��(�4��a�I�R���~�P��|��=z��_��FV�5P`$��+4~���1��k/���u(�@�Ϊ�Hv����Q��Vl�A�l�}��K� ����@��|�y��]\Ƒ����B2��+M0!H%��+��\����\��tX�K�t������?5BVyX�f|��$��(s�2e���o�����C8E����ⷌ�L}`'1g ����ԁ�Y-��i���BK�r0�;FX]���_�Z"�ɗ��X�Uc�)7-`�K�����ֳ�߲7����q�P9�N�4�b�2�k���ױ��������Q�y���A�����Ѹ���Xjd@�R�C�q��jݢ`T$��fe�s�G��4u�o��(����´<��aW+��"@�p�`)����f�	c d5�r]Έ���o�:�R�`�x�U_:擾t�?�RG���%h7X�E�Y���<A��V�;Y��KVZ֧x��3u�+���:�lIQ��3�|�G��
�=��&J��Ӯ-x:��^wx��݂���C�C��)��Kt5V����Ez��n�*ǯ���"��M�M�W���<be����-�i���qK�V��y�2O«���u���6�r*��Ҽ�\����ڱ+�nG�c���.9O�B���y��!�Н��k��q|�
�`�:�	uW�2����6Vt+��~f���p]0Z�%�M�ۑ{.ʌb�%�?֧��
2{�,�+ �~7��Vl_$v�֘;���ҙm-��7�ƈя|�K�}!�^˫�B��@׆0�b[x��t�[`��4FOx��/� �}��=�B�5C,o1�{�rӵ�3#~#�1�?���Q7��AĮ�X$�T�m��Z�`"A����e�S�f����2H�L�ÝS��H��G�N��	�c�e[���Zs����O)�L����#CW��[�v���b�T[u@����, @����RŘs4�/������Z�z�	Z�d�yk_?-l���z��&�o��U��f��Y��	̡��T�*/��G�f���+�0�/3�y���:����AxX�?U�X�9�N�	$�֤��h \�2U�Z�I�eA��+B�TG[�"i�* I�����H���.j�Q��H���]\Jz01����}���N$&����z�]4j����w�W?�! ���W�+��N�,����\������RD�&])��/D�F�����j�a�ZO���枈2�E�asMt+?� k���ji����T�x8��@kK��S�?G�a8��7c��Lc�����\��Ȕ�
,h��@uF9�e+�+'�d舖�u����V��nS�D��[t[�5MIԭ�z��Y@WZ�$a���I�0��:���{n7�,��5* y:�"]����8�oRPpw���`w*{๡���e:Ѥ=��������Qy�&f	��Z1�E�H��?]BS�:2�� �"��t�+M���0^���p̥�Ųb&���0�M��'��܃̅V�Tt6��0B_��ΐ᳉J�����T�Q�b�
Ѿ?��6M!0���2��tb��(�nE�c?�m����֔D`�[��^�l�z���攴d�0�c��!jf���ǽ�32�WKO؁�@C�2pڬ6�BX�и�7?7���N]-J�\�řg.��E��^}T0�@3=�B���s��kV�gXf�W�N��O����n���p��WTI&;2���ޜ�I;:�;����UnD�C;K�p�f�Vzm�r��K�ӟ��}c��O��*��dJ����)lLj��c�b��k��㮂Y�R-۱&V�ݑ�bR�'����$0������7+�1��`����bǀ�4E���v����G|�P�ܯ�9M��)�c�Ą����Abx�=�fD�7� ���gƂ�xz�J�݉��r�*�:;;��=�ǱWa9�@`�W�='�=f4d>�\{�\����1��(�:먪�ƍ+u	tD��tg��"#�B�w3*fB`D���-��O+���=��7���~���v�77f[�u |�/�%~؇�w���y�X$1��g�#�"�
��G�&���S���O� �hڊ((Q���T&!+��Й]�Z�ڙcDf ��8�hJ���ݛb5zh�hmZ��[�[g�߸�E���P��!Q]1�5�V�~���*��ۺ`��P��u�*[�+
����;i�6�sЀ��#4.�AB�+�l��Y�z��}��,`�~�I
J2�W�|�)�>5W7гsaʖh}h�%m��%tư�/½���01ȁ`~g�(岦y��������0ϱ�8��ZO�7b�G�L C>���3��N ��6��"������>B�@;x�=p���ş�tb�ɪ�yye�����*ȧ���\�35��?2ުfW�D��4�CFz��vt���^�����2��"T�5��
˂�8�"�j`s��v��7L5)��5�<�e���r5�k��������r�1+g��_���5�V��+�"��ӆ&�t���uK��Q�>
��y�������9���I��D�*@ǅ�0�=��*(�U(�{�F(ݵ��ˌH�=����hgqN���(s==���������4��\XZ���;)��|^z�5��ۗ�`/�K/��E���*ZW'�C\Dw�h@{`�es���A�/��3�y �Ź2�t��[���5>\�"�q����ٹ(��G�CY�A�4X�@�
���7�H�&���E�H~$��B�̵U�k>)�oO݅�����:�7��o�Ű�����}��ol}��ZJ���V��b�J�G�p.��F�Ӝ4�3�C���gy�
����!l�KQ6�-#7 �,W=�����A���췸�0��Y ��
K��F,���՟�������:Y�ΊUeja������=��Z��k��� �9�2x3��Y��j���2�&�xj�����W09�L�M'�r�jpC�����I`j�X(bN8��v�R��5�л����ҿ����w���JA����1�x���(H/RҞ���Ex1��7�G �*�Ot,��H���Y\�Ӊ!0�e��{���ļ����O�2s�d�%^ΪcD5��{��&�xu�E���k���lJV������}�"�
����E�#
͠�z<u �ʯ���Ѧ�����<+��!�X+���B��Y�
۔���	�Ko��(Q7x;,2��T0��c��/\���A�2�)�,��X0�A���/  S�f�*�������M]�������u�.��.Q����]��q��1��:�T��dʆ̀� �@�!a�ہP���w��Y�ۻ�g|�U vI<�W�lV�s��׀3�p�b�\IMך؟k7�>��f�B�T�'���j�7L�<ˠm@$�h�������c�#�g��m�Z��N�o��}�%���y���xa8���r��]m�.��M$ˈ��/�`�(���	�eKש�ϕ4@��\���8��F��:��"���u�����F��%�ei��ޗ��sR����a.��s��a]U��+.P@X���&���!�C��jB^`����I�d-�P
��O#V��,�t��w|�Q>�=.]�S�ص��%��Ӭ��v�q�������`r�M��)���<.�hlN/�#{`�JG-�A)9Ī1%��]��І(	:I�˰�Bvd�0�0��;�κN	��0-�M��3O�����@�����$��:����-�� P����P��K��h���^K:�A
�C�@1:�R*�fR?��v=�z�:���6�q9�_��͵Ⱦ��(�^��.U�d���� �im�!&�ĭG���\��OXA��S����9�o��a{|�j�g-�ݴ�Į	���Wg�#����e�w��vG끅�1_���j�X��V}�R�^|"Ѕ�����F��Kc��˗C}�0����G����ʌ�b�U�0>�j�\���NO�˜���c6-�:�6#�)��I��xr/S�n�|��V�=�o�����?��|=R1ٙ���n�U8���%T�eK�ʆ�;�~s�~��Ɯ�U������Q�JF��⩣��W)_1=�j'4�
\�����@#efgU�@��b�5b 	�+']?��~,�i���X >:�k�ʫφ)K�43�؝kg1�R��&�������<�SW�;�@,s�	ۭ�]�ELW��]|�ؗֈ�������O�TL(ሻn+�"����v�~z?��̛=	rF�R��K8pC��G�N�aQ��Q�d:���H4��SK��ۧ��g���F���	���0�������.�[TW�ɻ��ɷ}ձJ��Ho142�4��ѻI ��W��->��Q~��J2�F�Kx�Y�ƚ�R9S27��}��v��L/]�࢞K?y�rB܉���Q�3��p:{��% /��fϤs��W�>|Iޒ��.���Xu��~�DfK$ 0���X�c��qP5�[��ދc`N�p��bB�C���*fּa����dw�)L_��&�m|q!�}�¤T��\A���Nf���dr�;e�d��7�4MT.��Yl��]�^0W)aW���;�=w�Z����()�XJ׍����+~u��N
�9�MkaǹM�Ǿ������ڞy{b{b�r�&l��|���h@ޗ���������0����
�O|���XR��؊Џ��������,6��ƾ4J|�ޑM1�fU�ǚ��b�FYۧp��_�&��ˬE!�B��/������mǩ��u  ��غ��|�T��q)s�z7��\i^'��U_C�ٔ��7m���I}�=��a1VB�1��j_p]܀Q���{��$�/DF�G�l�k�.��Ȗʦ�t��R��\\59�/3���'����R�b��}kDrC(�b�H�i���U/+��Q�:,$��+��?��m�(�of�����_،޷�~C[��^��ֽ�m�Ro0I���G�L���Ru�����G�ؙ��tg	��&��,��%�z�;�.��tE9�	}(����t��P��� G}jjY�(�'��n��V|7�bۃ�|%��O�`��޾�-*�=Z�=2�ݠO��������������j�@'x�4����A�%�	�b�2���G������w_Y���Mw1���ݷ$)�@��  ��ЏM�76����K�\q1p���Ll<b���Te��R |sp�_'�=pg��9����`�,������~���� �)�'a��>�bC�!f�A��܊a]�8�=�7 �z/��L��A�B=b?��琱�'�
"��G�!~��)�j��)k�}���y3Ԫ�0�%�ǞS!��wX[8�a\G֋ǀA|A�*r�����}F+m�Е�Gr{r�
S�MV|��G"`%�J-)fo�bu�����][f�8>�_DG$ �r�3eZ���2l��G��aD*�f�Y��Y�"&���eH�?7�ss��h��J��v5�b�Z�O�F�:Z:o\�8p�ފ�����Ksĕw|�,����"�&� W�vo����)�)#��Q
����ш����sXU�ʖM IQ!¯R�Z7t��������Q!��P2Z��~���]=��ÀY��{�`��b��K[��R<���I����&MQ^_��j���0��kQ�RK�1>���
S�~*�� �[���0�=
ZƼLR����9*PY;�~����E`���<�����qV؃Y�~�_ n��z�>P�5
���Kѥ`1��-̸���|��
���#��OU$D7�L�+�d��9��N�^�B���d�i)l�d��p�����O���]���3�t��ġ���(io�N�E�#2R
�)uD[b�I�m'0	��]O1��u����~S}1>;���wR%X�`�C1�A�Z�\���vHFD���?y�)�J�!dkt�5nt󭋨�����w����0U���LqZ����df7Mw�?Ǖ�����^��ӫ0�Ӝ�����W$.G�v�4Z���A%y_�_��;h�.G��c�M�/����hJN�4�p����)��;{ h�s�@��K�����h��A=�J�|#?zib�رl��.�������~��6oƮ��r��ߣ�OD�0+fg����K`s���L1X���<Ĵlk�N��z�)ۢ�:8J��}��K�v +�;JXh&)3=��4�̂D�C�*�ЬCpgaK(�U()lW�X��hq�+:AN`-�]v����Ǯ�Iht�Q!��:ox5�/���,��ϴ�X�Z��Y� �_x�e�%w��O����oa�I+�e���G{�̶�:� #sR�>o��N���/����߹��F`4	ˉ�y���k���}��M��ypX�[<t�B�^�����0�!���p�B�ۤϋ8���ߍ���8q$J�3��DU��5��A��=u��ya;Һ�>�<�xإ���~v���ۖ<ԉN��6�ҏ�.F#
@]�d.�PB����p@uh��<���܏`k�2���SvV�� ��2�����&I	�=ϴ��t9Fݮj}K��D�|u$a�m����$λ�K�"�A����10���5���W��;{Q�LΒw6�Ѝ�h��u�Tc6���$�0�$�K8N�2��}�d�}��w�i�'S�^❩I�Ym���0d�)��Y�E y0�<ZjY��{;���$M��xX���{nU���<��@��4B�i�{��ߤVX�7]�4�_�:P����Ki��B�k���an�=�������8�K��\�1Pt��Ž��T��9��#��I�����K\�k��ʩfq��Q�K%��vv��q/���� � �@��v��t��ZE��d,@�0wZ�����<ge7��+\�F7|�E�3}y�����T�,���jn��٣�0���z�ɪ�~��dyW�k���m���(>�R:y��&8m�,Fq�&���_��@���U1��J�_�?�����	�9E�Ϯ����)��׳��`'�i/E�@n#�47s�Y;��.���R*�f��CXs���f$瓷 c�@M��YbS����7;�:���K`!a		J�ak��$T�u�>�ĉ0�d�޷r�����K��=��.���oL�>��@�������AU�	p�T��;��I,����G���x�.���%;1�5S�� -$:H�?�s'V������&&f�=k�$
��ֻL�4�:���*ҡ�F ��<���lS�sM���1���3Ӗ�l�����S';�_>������J���_(]�:ꜧ@W� 31c�q��v�M�Rn�]�ƚd��d<p|���SB�X�sL�<>la��-�p�;�b�� I��g9L�~��Ί%׹-��@�N�h�M�l��Q\g{�H�ߞgJ��5ƞ�1\��Ii�T;@�⌸���A��-e�Q�����_�&�Y%�N�˿^�,��?/>26�=w\�����1T��O��JV�����1��,���)��:T�����O	���</�l3��+���a`��`f�no<f� �	[`)P�n�iȻ�0��4K}��� �l���������0�n�m*$\����SJ��o�o	7-��\�J�.�+�6� G�-_h��Y9^��5G�Si��O$�*���u33�?X�@̧J,+~�{>P%J*l��H��K��(Nw���8��An~�y�|ՠ�dIr�XȦ�1�������4�~{V�~�QɕN�.ě��2��b�����l�.;��(�P6��%l��� t��Ϻ�jr#��wͧp@�� ��jDf�����t=�ٜ,�m��u�L��o�C�6�u�)�C"N�d\�i������JV�F:< DF��DZM6�^�9��}���Xb�m�ֽ*#��3t�a��������>:z�}�� -v,�x1��!8��3_��cǯ��.e��W�#�J�n�DxC�+��Jʍ��,����i��$eYU<u"^��ɳ�X�Ǒ��؏�r"/���D	
�vԈ�X7�Y.H4k�r���(`V��
�ʐԴ�	R��WSv-�S��{�z��/!��۫[�[2�e����X۶�/���(�Z\�z�繠h ��L��4��6N�-��D��J����;C���hټ�_�Y��|;\��
�������0ٲ�=���� �D�8��X��8C���8���7M�@�y�6Vb����4�Y���߈,WO.�'Ӫ_�eUb{3����[:�ҕ�y��.��oL[Þ�P�q�f�oݽZu���r#���ɞ�9)�!�v/D-�	�������yD tpf=�^����t��xC)�dO�Β�x�f㱆��v�e��e���	�~
���A��#/-�SB�Ɍ�^�x�{	�C$Gg"�_�t qR�O5����Q�)�Ug8��=<I��b|6h���b�Ԩ����	������'�n�r�ݶX���r�ۅ�%'�w�J
��9�H���1*2�/��''��ktDy�Z�~7��86��d/�^�!�P���Sǰ39v���s�H�	�� $�������C*����}G;���Zu��=��S��4�U?�̤����$vce�5�ȒG���L�����<�5?3t��A����TR<�숌T�g(�?�����;z�5���7�� &���a�-؆�pz�q=F�� o�=��s��aA�o
;��f#"��0�qd,+��Kw�5���G�1T���1$�~E�B̭�6M�
k�|������-�Q�E7)V���}���T�����Tٱ��&d���
S�V���G��U��
-�{�gz[%�&��)K�su�O�j>���<����	���$������$�����Vz ��<��Ǌ��>��}��쑅*։Jv�bc�~�4���^����g�2-ea�*�vzu�M��% �>\��V���
�Q��܇P:�lh^�=���_��*0�h�*�[�c�|�E0�#0}u��D_Q���Ye�"4���@��{�L@4d���*Aa�q�3>&��>άI�����2qr��=9�!�����g��������W`z���n��W���ܳ�T����PWfEtAP�2��y�ͺ`��F&�T-�*�?���������{iN*�w��⊲tÐ:���/�cNe��EB��N�,��K��8�cg�/U�ϣ��uk�4��%`e7|"ޭ��}����u5:��w/�>=�.P:WLN�N��`�>sJ�dD�Vi=XDvS(�Z]��|'9��\�,P�� ����Q&�л�(�5,������"tM��� ��Q�y�/v4��sy��lF��O��Ud �د峀5��@J��ڥ���8es@=_��ؘ	A@	���9�-!�U�U��DA1�o6S-?�h�M0(��n�-1��j3t�ތ�\���V������Ɔ������3��u\`	��#�������E����foI	,���M�/�m̟�#M0�%o�<�l}z*nR�њ2�\z�3m�ue�dX��6�K�E����| SaI���]F���3�Я N'y����9�
����Ǿ�p~�R�;��>953�;�I���dE�x_�P� �]N�T�������ʂ�M�X_�k�}���C����_�{0�h{6�R�%������4�(ᕜ��{�� ���}��%bh�$���ұg�_d����Gz}�xo�sq����(�{��f
�^�Ζm4(�I����������A�QI_}>�"��E�s�Y-�ǠI@6�[kwʻfaJ6����=�X%20!u�e�� ߑL��3I��5�D�-�X~:�n����Z*VT����j�@/�{0
Q ��3M�m~X�3�z��͍�E�_�� I6|������)�n��Č-B(��4����]���b��?��_����I����J�2쟲��}2n�A�>51&-��CP��p�����a`�K ��� n��"��?�`W�������x��_�G7e�	����<���x��n��)�OZ�ᶔ:��/1C���Z����*�k���/؈�d޺��R���X�[ʺ�Mh���%Α3�e*+Ǉ�<I>�0nz���:��[�0#I�[��?��7W��Z��(�w��P���b�tب���&���s*Dx0{�n|@�[U�V�Z�R���gvN�$%� ҙ�1$M��8���2]y셏K.qp8Z]�gMpPݵ^���89E�K�ZQ�h0�_)�:uJi�|�s�*ƈTc^��"�,}(K�^h#���ޭ�p+3my�I
��}�ZG�S���9?�Cx_��xE?��(y%�EoHe�R�P�BKA�o�yοO$�}�͝Buc8JK ���!ľ.Ҕ��֖	Ep߾r�%����[U�;A�yH�Z�{7�_󋾾��+��=��^���.^{1����b��{����R��tcH*��R�/Ѵ�'���|���opJ����3Gp�r�+�E&������� ���/�j`T�9��C�26<��Y=-gL�i����!�b�����C��DTɧ�`�8WW!%�P������,�/�X����$��%*c�m��W ����>=��1J��ij��y݌O��%���bTϚO�ô������Zأ����it���tq�������i�GhK�TU<sa�`~,�}��8����m�o���ā����\-��L�6$=W����)�0��V`��&��8��&�(�	�Ɲ+�����"���)��B�ϡ� �4�{�A�',u֔�qc�@զ@��:3��5�k�f�,��1�L_�5�DQ�ᪧ�f96� �w����uΈ�u\�'��ߴ�<�Q]܇ZX!ʤv~����Q����A^�aa�U;�MH=`��0ӻ�m�AI�&��T�AZͅЛZ6<s.U���=�1L�aaVZ����Lz�����9�B��H� mN�rnά�F.�sI��<E�� �Z����5��gR�oL������#B/⶯GT7b,l$c\?j����N3ov�y<���K�۱�ۛ��TX������n�:���ר"9)���t7�o��=�u��z��}4�_P{j�N,W�Sg�LL?!�C:� � IW�v�o��t��e^L���a��e���C����hp��SN%��PP��u͓�죄T�%�䯐~���p�`V�G�CJ������=ς�@�j�	����M9?~_�#k�G�>���H�w -H�G?O�[����?%�Y�笣��?k�5�~�d��]F�Т/ӽU/+������jk^�n	H[@ߛ��7����@ro�9S5ecJR �[�Vx��j����e���\�2��lTA��ߑ��S���p���>��cU��kw����P����eXf��6{	G�/Wd�SF���|�%�;'C��S�R�f6����x��,JA�~*^4�EVr�v�h�����������Q)�RjM5'���\�U�z�� ��$��iq`
f3w׈�m�n�]W`��,��.���~�(�?0�b�ы��Ø�l�
z,Sht.{�$�����f�	���|9��.5���F�ҖL�p«S-�����q���w|S齎���w�exL��J�Q`�� �[��l1@�pTr�"Z)�'{��_�X9��o���B>�q1At�?�,EݧF�%f�K{x����o�M�G��ӎDK���a<N�y�;����1<�^�3U���.�%9��=h��Ӥ�Z�]֩���R|�Y]������I!�`���"�E�-��Uw�=�5��F�	G,WD'[R�,A���|�ފd�f6][�^q������'����Y)-��ڂO�}�6���0����lG��n�b����6q+����*:j��+�CT�A�K�&G�hJn\�|k�%O��`k&��Y��]�/Sʺ2y��T/3!�L�����C�踩p@ν���J%���bpQ0�'W���[��,��A�H`�>c����p�9r(��{lM���"K-�6��+E�̙ݠ'q�R�ހ��wӲxV�0�&V�a�YŨzw5�g�8m~���On\����!bW+�:}q��]��흓Þ���?lI�l�|�PuG{�����h��7�,2���]dȾˍ�@�L��o�M��[�o�R�;���:�J�����}�2���3�Ȃ��]�v-�_��Hx�I?�ᾊ���Td[_�l7���H�1��d�nO�Px�j�ףqZ�����t�e����($"��-�>������Oqf,쿓�Ŀ����jَ�[�֬�͏	�Q��v]�⎼ne���M���M;�RQv$R�e�Ä�����Լ�2#�,�����M�cߵK�0���ͣ(���N�d�8%�Ԍ����.�$~M�Up��SHz��`7f��G�����9>��������f��-Ew^���ĉ7����.TT�_�Ҍa?�!ә�a"���9уs�G�m���yé�e�ձb��r/H���+��W��I'6$�0��i�_�9I�n'~�z�;}�է����~��^˻v������e�iN����c�����Bd*�T?���OA��aɡ�_�T&�ML��婸G���sv����r���̶��E��QD�Q�t��d��Z�z�^!,�1���e9Ξ��֯6ܧ ��~=@��Ph�#��3Q��F��N]�?i�<J��c;��ߩJ�@D4k=
`�|���F�(���|}��޼�^��<�m?���Q{����H�{Xx���I�	k��װ[W?�NUx�f�ȹ�g�ȃ��|t��|�yA�G����;���.�����L]g@SK�zp�WT�#]����H�%@�*R�HU��T��� ���*]BQB�Є�B�s�����_����g�yf��l�5�ʟU�����&IN�Ck�����~r�}EkĎ?/n�SU�����荗����X��7���[w"p���JzL;�^�"���ފ�j��`I�;��z���R����(S[Hș�Wӱv�xq��*K:k���#�1/ialU?���3����	���C\�d�򡶹>��\I5Ë:��Zx�bП�x-�#C�τE��:�E;A��A��!*��Rj��2��H%��/���,���%M�f&�:g?�,�B�F�CD�1Ĳ��oNm���h=Gm��f�Xv���S�0�Deݭ��P5��.�ZC���0�5���ӟW�pդ��E`���\�`�+����[�_L�/W��s4�u�p%�tj���ꃡ��<�aL�L�8m�����������<���Ǔ��,�¡չ=К>�(շ$�����F'�<CG����`ӛ��_�����|��%���ak0�X&6|�a��ҀxQc�𔲋�/d\�j�S�K#)h%�le��[-8��s;�^`%���9D���w�hzuJvP��UX���vJ���{j����w�{��?���,���w?�ΆPY���w�[ pgW/�F�à�&|��c�h��{�J�*N2q�JR}p��OwkON�S�����|%�c�_9�5�ܘ��-�㿙7q�H�L�G:���'U1i�C�x<�Y�����i��n���w� ��V�z�Q0j�����9�����C���Y�z"4D1Kv�x�8�b:�;Ow"o=�ey�ѬL����2���������v�,��q5W0G"��,�c�,H~���Y�=c��^������Z��Y�ŽmG�[�IX*�y+����N�k�2E�2C	R���b�������"BjI��+P��O��v�d��F[�����/�Q�N6�BO(���p�j�q����TNI�De{|��]�q�	����_dw��/����[��m����d.������d���W�G��
�� Ȼ�k��/��Rv��~�����p�1����PA��'O�Y���`�Ef��ӧ��^��3�^����ͲK�oM�@5��im%4�C��٫0��T?W!()	j,iF`:�dW��aQ/���k�S���R�����S�/�:Q��z�~��_ӘO��hN�B����w�臒/�3(��%�]���}������l�;S����6�#��OR�2���)Kfd$�[����Ǝ�M8��)Rᡄ?�*[L�$'�tL�-��d���$�oX  =��w��7���Y���jK��qP{�s��h�R�ehȍ�w�q 	ժ1ۅ���rL�.o:�դ)[*�P��QO%�`��O��HH �F�ͤe5�Q�p/���b3	���EHL�#n�{.��FD�do۹?�j�����<$2�CO���kE*�~�����Y��Crá���/M�k�gቢ��/:ܥ��82�I=q�ܨ�#���my��Q�~S�\2(��`:��p� �wH����UR��j�nOB�CO5��[K�\5}��6^�ýt��Gv2U�=��rM��mԺ��K��ˎ�rF_|��Jz��bה�,ڹI��ڷEY8s��˗]̤w>�b�@��r�H/j�iLY������&�r������l�ܝH1n�R�~;
״���KL�Qo]e�[TVx���Z�3�l�V�����2U�
��g����I���:�w�4ńN���;*��.1�>4��{�LLf�잦|��7�|8ו�*��X�qys����F<�n��@A�M�0g����p���j��c��֛�N��}�'
y!r��ñ�x�4a�RH���5�<���kQ�i��]a;�ұ�ר�zxv���G��\���0�J5�!��Gn1\[�{Wlne� �ֈ63力������:�j�A��,��nZ4��:B��!��~�s��E6��~���k9���q���)�uAuQ�Bߴ�w��s�}�'�'���1S\�����t�s×r���IGs�!?�o��n_Mk��l$<�YX#q��F,��V'�gT�O'3������홚S'��u�:�o[xڂ�֪�nb��+$3������G/��y_3�|a�[TS��^͕l�<m ګ�Ng݅�-��b��ܧ�aGX+B|�``��dm4��^p�.b�o��B��S5��B=��C�4�J~�_ۚ�",���th����]�$�v��c���n�P8d��?7���`��r	�R[�;E*f�M�F�R���e�M�����K�\j����/�����9 ��)h���r��T�����.$�4�nLn��¹�����*1��?����s��e��{eQ��S��l�����|����,!�:�{�~o!�J�e�Ulg�FV�>Io��0�W3��9Xp���ҽ�m����(�^&E]��-�*�{���4��nǔJ1S���
6����8΃�߇B|B��T~�@_D�a%o�������exa�����.D|�(�r��Q	�~���~�z��0������@�?T̀�t��i�.��x�2,)����q�6�~V��:�g�S�+�J`U����������B��I��Q�;/�wj	����*� ��̝�.�f�c���'����졧����K=��/���'~�͝:ع�͌������Oy��8�����H�!)|�{�uS���$�t;-�:����.�X?�=�,^Xmdˏ"�=���y���j<G���A0�<��d8����������#��MUbp� �irgP�Wv&���_�Ty{����Ub�a Csc�
�mK�F�"������lV�(���X?���f�e�j]#�c�}a�k`3� S��%��T{7��z{������j;)��&�[u@�ؘA���܏ˑu5R���<-}� l߻��(^�tW6�&,�*����{��R�ù��g�����&�k�Hy%y@v9S׹�+�X��]!�rݗ"�Dn�ٔ,尞��.�T�v�j���9f� R-{�폿F����"���h�rs��5��{�$��6{��🙏�<>z���i���&7g������z���$�2z�V�a\�i�_"����^�D��!�=p$#Ƽ#�Y�5�;�ʥu�DR���3��\y�Nuk"��J���ߔ�b]��	������� U�:�ͺ� �OR�FKLב�2�{(S��)���,�6��4�Epq2Q�����ґM��&yl]� �9�F�a�ȥ���8�d����>�:���=�9�5��R�nkF&�i竷?b(�4n�IM����FU&��'��Jz��E�{ y�6���7�L~��[d�0'��tXVb`���(���Q8/�����K�Y���b��6J��6a�C�в.aN0l(����0��F$%��)w��4A�C!"
��g�ٱQ]�j��O:ʮR��SZ���(��j��<�����M9�]m94�!rlA��U����M�YC�Ő�N�ڊR�d)�j����BOdꩄ�����y�wI�/�A?0�暆x��j)�~�F��K��r׍���w.,�P<靬��������� ���l}����#�2�u�x��;t�T�@پS�q�q����A�܁Ef��|���l�׀Ph.��h�\��F�g�۫.�r&a������-r�\X����t�0M�iD�v�@�*�|y	��]�MO8?^�H辐�6&(.\OpM��e&���0}��L9n�F�j�����Zy��(?��!iy�g*��u��]��A�H!�{�d�};L����'��_��6�|�z�#�R#�C'�ö��F��&"�+Q�&^��@�I��1P>��N���2n`0�Nh�q�8�A[Š��9,*rf#��3,C� Ȟ]UW<~������j��hZ�����)�)Z��+ǜ�����閕�����
�J- ����m�a]&&�*)��^��g.�5�S�(�uR��y=�3����Wz��Op��LR*]
�F4X	8�᡽[�Cjʳ.#�A����Jg�f�|8���m���`$���\����Մ��/@(��髊��B{�81��,eg:ږ��^ؓk�����)>½qw_qcLy�7ִ�����*�F+�_�Nz$���%P�bܡ�mQh�{�QH1L�Kr��G.;JVPP�ӻ7�d?nw����)���G쎢��:��8q[ա��@���##t�~((5��Zb���g�=�]
���:!T.ܨf|~����["e����L3_��s�=�$=E7&��m��w������4]�wvDu�Q�Qo����(wJg�a�'MS��rW|h��?���ri>!���#���U��j�k�.���x��ZW1`�9y�x?��Iʩ����yR��g���P� 
̋��5����/ov��+X�Fp���^��؀��=�T]נ����)��T��.0
v�����L�)�Jn_S�hn:S�(}���eV7�J�F�uj��;����kzG���nρ�����g#��{�pW���������("��S�n�O��r#��0�� mM��
����<g*\2�Cʪ��t���1̸RQt|p�DT�����9�.����l���2�m�{�4"C^^uN�j��� z-�mexlnC�,Ě�mM�	�2~%t@}�#T���1ԕ�� ��2%��v�>hD{��m���9����0})*���ٸEr�ۯ�_w���lqj��L`�2�#���7�����8�Zbo��!�"�lI�Q������p9�f���z�h�:�3T:^�%i���CL���V��I�f �����
 ?�V� ���ٯ��������"j�J�j�1`�+OU]�	���&��$���o� �>�r��ӫ��:T0����{�q�[!A����P�S��B_5��	�.\.x-�,��&�cQA�۩<ˏ�D�t�����x�}�;Y,��s��,�&y�_���2��`_���������0ec@����U���)��az��ś��DG����z�@?��n�ݬ� �*1c`����|���U=]����>�z$ʏ8D�O����1�L�Y��pTh�s�؞vL�z��2���Ӳ�,8������ah��z;���������rz���e�$ߧD?�z�qAXJU2�4�xSx����ԣZ[,v_�E<���A|�T �*m:^�p��B�+<�]NԵ$�E%����1fU�1!�8ꦵ RWQF�P@���['�z�{����L\�g�Pu��r�MExkOB����aJ�xi35˒�D��&%�Q>o��]����j��r�vmI���-{�tN��_i��.p�c�*IN�(v��=�K��4���{1�� ~� ���N�MNޱ��֡��,yv�o�%�<땘eQ�n��Aj���E%���:_�t[�|l������ش&�m=KrI]"�J2���v.����/B5�>�����D:�*�ѵ����cB�3��j��
-�md���F�w��SAv/�D��y`�X�BST����H{���y���G.�:z�r�Ʒ{�[q
�g<7�N8�r��V�����?_��=	��aJϺ*C_�k�J���2�O�	������N��w ������_V�ߌ3z��#Ǥ&��T{����[;�q��do��M��nRC�@���i�U���&����>k7�\pB�>���	?r#3͇'N��!�g8�S�2�+�;�h޵�M�.�1㹕z����% F���V���F��Kn��H�<�*�����.{K/jq;Jͤ�Zp��I�`�}��3�/�veZx��g�� ��XL(��	g�P}�/�?$u�KWn�x�neMyG�6���j7<��C��i�n�:TmE�y�
�"�����Y�DR~/����	쓜�7ZN���ݪ�u�_�A�+<m#	.W�*��[U���k�/#?����|E n�������P&8}ڴ���١^�T-��_�CC�'5�(�������8r.����p���0h=���"W?��九92j�Q	�`#8��j��:&4J�^]�Lv�ڮ"�^`2�}YnKy�`����j�����,3�f{�+���\�"2n�^(��}M���΢�}�ۀ��8��p����
�Qe`5m�������M�򑬲�	�K+�����%H��q�É�����,�X�K�7�lPsç�څY�
%K���K7�����r���k�5�|���������X�>s�V��m�&2i��Y�>f���j�[M�QS�����ޠ.H�ʻ��[ėԺ�c�D�2�[��F�MI�4[��G�ؤ�
e^k���'�H�)M�1h3��YL!�J~d��#���i�hu���l��GF$��|��]U�(�4h�2��ת�:����P]cW����9��3���N�QI�G�L�dW'����˛�C#���N�\v��O\�?9���_���¸FX���Ϭ%�]��g���eO�a���	YJC�Т8ز!@�Zʟ�,�HK�	>�nJ<��$������y�W�`M�HSf<���a#���gx��P�^$�~6�-(74��FI1y3Ћ�gc9������+]�-�0W0�F$wΠJ��� ����e�N���|Q��m�]�jS��$
���C����j�2����/9�G���i�z77�J3�|I��̘��KD�����*����#��d����1�c��M�6nfk��y:|�f�慽���{G���lYa¼�9����痍��e����A�nGnj���G�\YS
����r�˸���������z�|���PY��~L�,[�u�Ӎ��z��2)4���}�c�7���"#u��4(XD����W�gs��Ն��Y�渽_���T�1�(�,�M�u��n������9 #���,�����Z�3���FB���o��IĬ8�dx��e�]�ɗ�.����Ӹqw�:�j��DͷM�gHс!^rݠj��W*���RTf�G_.k�qs�P�rØ�5���W*��,�}߷��%~ ����;��u3�9yJ~^}�ߨP����1��*�%[�6d�q�ɼ88�}���l�@,p�qP��l�;L�C�Y6���������C�{9�����oR3)���v�������l�_Բ�z�6����>�Qg��;0�6*R��P$q�CTJ(�W�iŐ�>n	�#T�O�0}3ں����0�=������5:�y@�d�&P� �ƻT��)�R5䗖�r���X������U�Z�o�p�e-��z�ㄇ��J,�����N�Z$���a>�G>��?M+_a9��Ѥ��\ڼnĂ�-	�M���Ɨ�3��8��^,������v�R��f�/�W���C�F7��}Ɨ���Mi�
)�ZZC�}��(�C��eٵ*_��~�oOIs?�Q�k:��f�!��b��^�d�Y�x�AQd�2�\�	�K�1|�,<'&�IPG��{���c9�o�Nyp���pA6��國�rp}o�ދA��ܢ�-��z�;�d�*�� 8)�Ƃ\
I��[&��ܬ:3D�E�lne�i�ť�]5�18۵��L#?��6��f��t+ �E����*���"���b����?�e�!��3��v0������0���nￛ"U��X���6���l���E�h� �b��4�c�>q�R�#ұ�g��Mr�:,9K� W�(n%,P�U�ۭkO[6C��vEwx�����K�)�k�^��:�fB�D��[$hKM��m���L�d	���\��u�gX�(�Pi!�d�������T�3BnrM��4n0�n�.w�[e��c�G�긆_�Ҿ���I|�;w3��rQwb��ln��0_��@��Y�Qu�o�x����<3�����R2�aBh��X��ݖEn2���(�epdT0��(�.:�A�˲�_�}�4-��P�	[��"�R�@Y�=?ˇ���L����d��G�tϘ��B�kD�|�J�1)�]?�k���T(1�8r���͘�[_�姧Y�J��o�w��� )ȕkn����+��)Ϳ���+DV.2Ⱥ��od����I���G�o��MQ�oˢ��8��1�JJ@���==fQ�����+�\	�x��gW$}M�V�'+n��2 ��ضi_�?�j@��1;Q�e~�,�=�vX����Dc��+�!@�W�7́����]��GG�� o*�\�E��4 ^-�p��`�j��綛���g���Ik�kqN"!y*�۫������M�hXq3�������LU/y4ÂWsbb��3���""\�jo��T����<�?03�0�|�ċ޺L�q���ejw[�bej�0�f�|���mI�$s&���l-<x��Q����Q���f��\�ࢥ��^rrm�H����n�@�٣R0���U���I�?�S`Zn\/�vhls����xteed�3S�|ߺ�ұi��@,|1'\�2h�b����!n7�������O�P�ݫ�XZ�����Ր�Q�Uh��8 �[K�����WVG��ip��Y��ay˽
R�h�oX�� �Z�f��Hi�\,9� �"�Qt��9S �"�����BYt'c�ٴL"�DR<�J=�9z��P
]�/$mT��h�����w�7|=IN;�MXk�T�)ﺆ݃�f��.����7e�V���>�Z*A�l�=;ԩ�:|�=�����J�M^d��J��Zښ̴�s:=�5��p`���Ȱ�T�3�����%�O:�ԭ�o=2�o[�p��d�x�`�)]L�<G��	(R���v���)p];��4�4j)L�&ni�~I�5b��j�M�`����}���鞞^77�@-���Z��XN�u�Sƀ޵�=}�1�<��'�X��ĳ�~�D�1�-Z*C�$I^8��UT�^Z�?�eb�|�%�?}�4koi(h�K�pZ��ucHYz&�Z�ɮ�h
�"d[��=����'�@p��-���VA����ժ�����IC�����:6�g� ����v�*�i͚O�OK/�?@�Ȍ6s�jR�念\cֈ�si>�,m��ѓ�)5�����Y������Eù�=����{k��a�j(t�	���R��j��K6HWٴhZ�����9����}
�G>M�=Q�ӳ�q���y<�⡱�Yx��EFOq�N��	��n<�:��r��K>�Q=uܲ�(�Nr��I# �rD��R�i%���կ���UC��Eg<�
��@��H��"��Va�J���}᭐ІM�����<�&��2�H�ť-��n'��s��嗇�t��-�H�\:�1�(\7����ď�V�^|�%ZǑvN`�ʥ}��Y��Jwu`$�M��GH[�/5[hu�ʹ5��0P��m�� 0��t���e�ǐS휜�˸)\]��`˸�]Q�������/��h��i<b�'��vdAG���+��h�í���q���e�%��l^I?��H��r#N�+�`�w�W�TJ�T(�t ox�S|(��*���H	G�f<�蛉�ͣ@�6U�S�#��!�tX�q�B��S{E��mu�l��˧�&d��?V\���՜�_)�S>vr4=�'3���H�MԆ������j������z�M~��OSx�jy�֣�G��m��0��cy�XB��Ǹ^,>�l��I���E:y��rǙw�<����s��%�o�s<���ETiD^R�o/��Z��WF�7�	<�t{-2@��:�V��Ώ�5�["��a���6M�]����W;����}�rC��=��<���B����T�~뾢��+Ktg����³h�9����+$��\��!�2�S�w"�D��u�m�=�Ğ]��V�ĵ���cl�6t\2��A&+���< �[��f����6�@�����q3��q���!��߇��τ�.
B,���NdJx5�>�����s�9�i��C���v��l�0��3�۲rV�����!�l<x���隥�쐊6���=I�6��~Z�#�
OZ�'��2C˹���W$+���z:.ӮJ��!�>�W��𦸵ȟ��]�7;�r3v�9�f�ˬH��\�P�^��䰾�#�;�w��B���&n�������i=�q�V�}��"$Y͑O3�M��c;2<��\.�Q�3@J޻�:��m�.�:Bg���E��b����n�'���)�Ma}�Y_z+��:gW�~O	�����ًɿt� A�7ɘ͸:GH�L0�8�,�4���"�tzYr���V,\n���+ �D� -^J�4-�:�ݯj�*/̥��3��a��L���c8Mw�"�0����n0*��/�=3[��`����m�Q�@RL�����5���w�`jøn� ˓���t����t�뷘_Ѿ����ʼ�r��{���j+�٠��m�0g�2��|�w|xhP���FS��>�ҵ���i�["K yzP�&��q�=�����G?��yK�Y���)n����0C8����J��/{�� 'Ɍ:-\Y8�O ���N�B�
���sz����c3-�F���Ua\;oh���YeUO�f{�	&�O��ٶ��"��Sސ�ָ�{&�x�Ǜ�׽������9:-x&�;�V�k� ӓ���4QS4�rP�$�*ll(��IK��]?�R���ȓ��*�W�G=+�Wl6P]n[zl��J̔C]�=���*X{r��FjLaC�<�K��v�0�j�|4��|�K�����>�����m����J~�Di��f�!�P�q��3��5�T�
>��bJ
����W=�	��=q�8�7���6��K`��U�m�T�0�B��x�m���>V���@�CZ��2���f��+�)\˯n���|�f�_s����̳����@h`.�k�X����~j�/Q�5��&��c�������A?�4���e�|\���M߱�0�vN���2d$K\2#Xks}Jz�n(�$���d=p#=�I�i~.�yb#��v�w4��{`�3�tI"N*˒*5&��U�9��h�n��_�0	���� Pzu\�lWn/h�-�,����14�R^u�����q�h4��6mR{6�/ņa
�qkc���ר�r�(��y ��-%1˯4'];�4S��wJ���2K�l��@P���Az4f���H�)�  ��c��UP�c�%�V|fy�j��nn�^,n��bR����u�ྼ�*N�}4dEyU�_7�.��{O]�>݃�8��*>��Mw��?�J��kb�{�t9����� 5e�(i?(��:ވ���TmuB��Ƅ�����YՊ�6�_��tF��̯c��R,Ym9���{��O 6����t�	y\�ԧ!n���	��8�4����(�NA�\���y13�S"\�Rk�b�����Xu�:�e��k���Mײ+BQx�<�4Ģ����z��Ew>��?�����)�F��
Q��k��e\��$��d����F�ǢK�����v߳_�i�c�~o�.f�U�œ�Nf.����_���P
�%��v�<�v����4+&��V�v珙��̳츝��E)��@����r�c�V�*�7�p9�~���^�w��;x��6jH>��{���m�R.H�+����V`w &��2���7�u�o����1}�u/8K�4���۩�z�B���ӂ������6Q�<��u�#�M<(~,`�C1 �����T�c(�C|��2Tx�*�$~�:���؈|�R�~����^�{P�y �W�W���8OK���Z��v~9����^=�k�qmJ��,�_�
x�+@��X�zpSN�h�����N���v%�~�S_Z����l[07����	�ҹ�3��0�@�Х�zG���ZG^�s8H��s %�����G�Cr&�V�&-��9uvQ���.�w���e� ���5��-.٠u�+�)yx
��NC���c��FD�Ip����@4�����[�:\�-��� j������,S�c���"��Q��THK��{�2�[,ݾ6$��e�Oy�*�8>��5�a���V��S0��8q<��L<���"�3���Ȏ�=�����a;��ɷl0�@�!��1W=�nB�|�����y$�o�e�[�*��9
�ۓ���v�����D\��1A�(T���_C8��ǣnk�Q�����z�6 �n��%����c���E �f��o��[)�;�<ƠX�%�j�}�x��
�mWc��w����-��S[��Ϙp�H�.Xe��3�@�.��F�����HCc���*�n�Z�t�%.��᭣�Zya��ae��q�5]�$l�F��&��⨛�I,�E-��\�cbX����o���S���?�QN���Ժ�ks�FHRl�j���Y��a���+��<�z`�-�3j�ghy_��Q>+�PgQ��vI_��b�G�u>:�����W�9S'}��L;���u~��,t&:�Czh��A��?����龜����옸��EM��>P�U����	���%��6x�uN�c;@=�
F[��1��l����2��m,�����Zz��ޞ_n��J������߂���	j���NC�b:%3>��nH'<�z��_a�����n�J�������3��z�����NJ������v���a�V��!��(����N.�ܧR_@����ur�]K�Հ�N,��N/�i����C#�ZgL($)9RWH�le���z������'�����J�B���z�ݍ1p�N�c�����Y}ݣ���K+�xj-Q���� �)`3d^���LD���^{Ę�
Ÿ6�!~m������Pl����D��聕8$���<ӳ뒝�P�����C� -wo�p��� 1P��waq@PS��ߺǪ�-Z�e�{���:��=��ۀև���+\�1 R;i ���"6������"�/�!�WAB��؂û�����pk��<+��x����h�mI�+a_�6KG���͓����]m�bd��҃wL�4�
P�v�ߎ�M\?I۬�ߥ�����)��K�k&^c�om��$8���x��L���5$.P٬	�0����H���	_��/f3ҼU�+���	��	��ՖM��񣅹x.������Ā˩<Q�7�6�k�,��-m*������C�!Է�~�0��AsKDJ����!���֝�)��_�P?��_�����g7FH����}m�2�)�I,w���v��݇+^�˱C��9Zq^1zQ,-����)B�>��U����"D3�x��C����_�������m�S��K�������h�aQ���ߝ.�����s`wu��aٔI^V��r@��P�{hDw��ni��7C%��Vϵ7���f\z��� #}���&�*h�k%�o���kR�\��i�
c�i��)��Wzw>��2�AuXg����i)�B3�(���~��a���Dǳs�]��"�跎U<p$g��˃!��Ѿܳ�G�.�=Ui��@|�̜>i�tB�s���5J��l
_}���rE�&�Zh��'��	'o�E�I#C�;��;$��|wY��V�?��c�8=���My-ˋ��Ňb��r(�������
�2��2�����r����wg"�d��D�Z�<x^�W5����i�^�'�~��]�ܯ�a�-4gVn�k䪧)���4��[�4���
�m}:��O+��6N I�꒸zǑ����A:� ӕ���A�]��#{5��AU��������mA0q�ˑ"�Db[7f������L���gMĨ6� ��	>�&����	d�'j�G�P�Y�uŞ9�X0���LjP��O�`F�#-��9���ZOB��]��qχQW�a�h�>%�w�x����0�?]��B��NB׳2�jeo|fWج��$m�zL8�8���傹�]��'�ý��|���{��~	�3��9q�sH^��1D)�	�b_V/�5��{�L/�B��O���u�����	�a��D|�ޱǉ�[UW����.=3������YY�֨��D
r7��߁�__a%cup�(�?Q���v����%�5�v�[5�VR�%���w���]�����������g�Z��r������B����Qz'�g�gәF����&k������[��+������+�NV8�%�+8;R��h�>�ޢ=m�KK����Jĸ��Z�.BJ%��U�vj/��^�Ul���s8G����ܦ3�c��@�^/:-\��k5�{.��C��rʩ�֬�/���ؓ�������(��{�����L#�WLe��o��#��3�Qc��Ӕ�$|3����Ck�ˏ�z��woGu/�{�͉@XB���חS��d�lr{u2�0.݀� ����#�=e���6�u��t�?��^r��ׅ.hOJ*��v�Q�a��!������\���Z���zr�=C�ϋ�8��J���L��$mK�	�M��u�Kq�
���r��?�/١+��V5��BOW!����u�!��=�j	"lҁ���`�/����)���Wf+�j}4��(,)怤zQ�;�a��� 6a��7R�"7�����z]`��gϦڥ2��#�K2��R8�,Hb�b~ 8�,��2k�+�ئ�ү����x}˒�����j���oy�h�j��\z�i���*�����+��I�<Qh�l�n,�q"�)�h�y�b+�~-v)X�v��(+&���U�މ$,z��˖�rM3gֲw�I/�
��NN����n��-%h]jah��L�.�rl�5�@\[��B�0���޳�?YvӘ3@��ϛ�1�=^c�w��O�~��Z6��H��	�]5�T ^�J�b9��o�0p��/{�!��R���Æ�:��9�����r%�h�_�2!C����.��aNw�o�8|P�,Q�-�W�����`�e��OU<��<zE �.����1�D��N������� N �:K�d-J���s�X�ǩY�R���<7�>>`~jݬ �;<C����߳��������@V�Cw�D�� �i�ɉuA���>�_pY����n0ѱ��dK���zg��|�G�gg�%������瀢:����C�h46��wPa�sML���.C��oQy�ޤ�lmBF�X��o�+��D���y���G�2Y |�k����w����"/8���`#z�1��E:?�.��]v-���ߔ���s��v���w4�<�eWg�?�OG����M�*D��	�	�X��n<uL�E7�eJ�0���L��̣E��]!7bQ{��D�@��k��)����u� ^!�J ��{`e�&�צjPHƄ`�� ���ek�Tr"c�Z:Y9p�������ο�D�|	BC���[mת�%�Q<l�.1�	���	��=jZ����� !����������p%V��Ȃ{2L�W� ����w @�e�0�Ճ'�  !����Hl� }%��V-Μ�K�dM��r�jxj]�Y��!�� ��a�y��}���<���{G�8�gN�����㗘��mA�oN���W�R>^V���c��Nʊ�v�Ʃ�W�� [��p�o[�9Xԝ�4d�$ߗ2;���K?�#U"?��É�h�& �!�3yh�t��'Jb�3�����r�3�]��� ƽW	?W���F�/���Dw���y�f����7�R��W�X�����V�i˦p��4�)5Z_\��O;`�n?��M8�2�#C��j�|'2�$�L�$A��/�\���hMkܛKe����9�>w���t:���PQ���Ć�9t�5�c��8��x4D��]���>Ϛ�SnepK�n� c�T2q�&RA�au����;㟚�wm�#냸��5�Q'D��/L����h�����G��c���j��<H^�����ۛ�D�,ub���v#PE�\�IN�� �C�?ﲨ�M��2���������Mg�z�j�'Qv�X�C�$��b2f�r�voX�P�q�x #:Y>����7*Ȝ�k��9�Z(g�k�,*��n�I�ټ�cT%+�8��$SߖbX{*�'n޽�p�, O��������W�h��I
5��cH�	�leo�Ff�>�����'� �M���e~P��G�2��1�I6���N���]6.5�s�Er���W�I�t�B�+�?�}�N�'�	R�<���go���;A���q&N��t�p�	.ţKHjhV6����S5��6Q6{=4� p.O��U�H�����J�>ݡ+���/�p�W��8_�žl������`�'�f���ζ�)�u]��A@]��Y� .+@�����q�Չˊ8F�V(��$��
P��=?�&��N�|��
=����ey��*��3��|��mrl�<ɝ�����9���N��J?����X�H�m�L�̬��l�/�)ܖ�nTÑ��+���ly��ﶤ��o4����oe}s��]O�9�ԧ��M��L���A�{jм87`v�U;qY�V�S��B��wN�
p�2��]-oD5}eUߺ�[��~W~H+�:A�i.����N�b5˺��Vf� ��X5�+?�U~�x�4Nw��[��Åμ���n^�I��0��-��^Sצ��?5�R���9@HH���2ܠ/:����K�=u߲�����ŰgZm�d؞��@Q\�@���
�v�I��[(F���@L�AC����z�J&�z�#-�f�<�U$���C���u]�������M|<O�@jLH��J�'��>S������U�$��N�?K�L��Y?�-�:x�<�^�` ���sb�H86$�`�=o�D��D,�����=t��S��[�3�x{1I�s^�.����Q��=QI�q���0=Π2O~ȃ�v;[2Yҳ�b׎ȀF�?'x&�EH:�<j<�:�u����0�8�L�G�ηؘ0V�=M��<�c�5^�C~S�G���v�_���+Z�����h�p�Ŗxg4\�r��~4%G؛�g��{���ng����m�I����i	h=�T��m�=ώCR�5�3q��!On��v衤l���]����W"�WC�E ̾��Z�=:������g��V�m��x��]��!���M��"�z$�!�qג�3u-����}�kC�va�=V�泽�Ь�,�����S/>�9zj��\��nGTd��4�?^������	�;�=�nri�ə��I㧐�S�Bu��(��[�?[WW0"��2A����I`��sһ'��H� ��svt=*[�W�V�)��(�[i���@E������~U�H�Ʀ���4���Q	Zƃ_�2(uّ�}����Zٶ�ƇP,�*���}-�-H��g�6��oL��DG;�W y3z]}X�Q�Au@��+[�E��Պ�'����.|`\F�ߧ<���gHI,]`�_5�&5T*	y.�`�@�pk�QC`�'���g��%`��	���y��*��Q5�Ŭ�O��"��\5�}�O�LZ���/��R�<Ǚ�����Y���&�����3S���QK�R.e#�u�ǽ��Dq���T,x�s���q11����f�]�K��Z4���}$��ɋdPd�	�}�`}�b-K�tW�o�w����H ��ߌw�֨`�(�9k�R�^N�����F�KRj�T�>�L���rn��F�g�q���ގD�O=j�TZ~3�3�="/����N�x5��������jj�@��("�T�"�;bA�Ҥ�*���(���B�J tE��4�I �5@���;��{o�;��u֚kι��guA���:
���[9ILay����Y�e��~�x���� �݀�B��lxE��
;\�tV0��|d����JF;,N#���#�k���?I<�\�72�5�+,�UX����lW�LKvҩ���*�eC��g���Tf ��Z���|����5�z����l8\Y$o��D��C7:��P����V�b�d.}�,�	/�啿�t8�����3` kTR��|>8�տ5��ok���~^@*-����{��P�n�km�}��*TM���>m��>��r�B����V��E]�\Q�����E@DX�
@ح�����U��^�sBo���� ��Ҥ�b��[F�L���0Li�9}�T�#�,Y�0��T*1�ߪ���S*����7G��Qe��*<�*�b8�� �7�4n+��dOU��	�QȾ�K��#�����초�J¢��t�����#3�K�b�j"R*/d�����<�_y{��%\K�`.&�*� �4c/VUA��B��U%����;�f�=g��1��fթ�ˠRl�␆�V�VG���v�� Iqm�r���y���W!"c�3��6����}V5����H�E��&�bbc��~�{���Mfz��3S2��qo�Y��rNf3Kvro�	�����em�!,;����f&н�>A���aM����(���}%ܨK^�hL8��'r�������i��
�m*��#�ި�xs
J>�b��џC�@�(`���*0C$���M�c�N��d�72櫵�o�/�ha�d$�������R��VX�*˜a�S�m1���i�%r�aV:����]y�f��op%��P����"�<P�͸�?P�>����kl��[7�&f�O����4c�����O�,r��wk�%.��$�eB�ŀ�'����O���7�{,��t7��fÝ�����Oob�|%p7��%���=[5�~��1&�i������A�?�X��!_+�'���Co��6̖ȷ6���o�B���^�6
��>�_��48L�`]u6j�4����>91M�D�I��M<�It�w]0k�j9rf�D��v*¥�DSlM��T9�E�}�I��(OY	�n�J�N5����q�7�'N%����0�Z���:�9r���+b�3x�D.��<����G��:7=t{���.ѹ��	��,���h��YҺ��,��&l���J�����r0��̮�N���"�>���Y6�x���i�ƙPAl���g�jA~�ĄK(�z5��'S,~a�ɢ��/[?Sizf"���ֺ\�<U�:�I<�cP��6:"����+�x^7�[�TafM���V��)����g��R6��#v2;�m1f�E����9������2�r�Na���?N_?�q�����݀V`�o�E�W�943�(���s�ns�Z��z>FB#/�efg�7���A(���Pb�X��.���K�÷�N�??H�"�����9�k����+Z�������ŘE:ঌ�y���G�$ۤ�ڋ]<Y�c���T�4��vP#��!�Ib{��Q۱�	�7��u7x�-u_i���q��9�4N���$`�E�ǟ��wZ�M�L�� ��1� #Py���b�М��Li�z���у�-j������[���5d[탵���ӥ5 ���w 3:�%?s��O��C�x�j�E����'~"�^Ti��H��7]<5����Җm'}m�=��N�,HU�2��*`o�Ԧ��:��Ur��hgw}��͍�!'F4qrnI2`��,���{CS,+W1!b�8��(*�	 �r�����6�x,c)sz�Q����>�,8X����f����Rk <�]po�����u;V�X?��S;���߯��� -t�g�?D�#pyIm*�14�W=�%����:��B�
�fꧢ�B�WO~��d�_1��:�CDe�$X�F(*�c	�)ڃ�,A�]�����RR^�6��䈟BO.�t�=)���'��H�Dj�eK}Ǧ!}\�YX�qq�K��̢:��30����x�
�䇻)/��$[o%��YV�w96�g����ES�os&~a���2�.9&�f���u��I����o���/�E���o��;�n0��D]�v��"G�'�ceKp����g� �\��Ԭ��}O�$����R�ud�Bo��m'��@Z��p>m�tI��:�/k\@����~����,�`��i��l�%�q&ދ�87黊>�)�5��G�!i�S��1h%��Ƴ�/�� ��dY��v�|�d7;\Us��l�����f%F>Ӕ1{	1���9�C]��mh��BqӲ�����7ַ�������(��@B��U�|���{�ؠ"뫺�TBj������WS#���3��Df���E'���O�f�N
1t�K�RG���G�t��6�O�V�L�o" q��q���0�Woѭ�{�D��k
W��Ơ��?RY��*�
;����>M�e��s�-�lc���s�1V��3~�̫��o�����r�"���N�i��q�����NoB�P+�Qof.�
`"Zش�?�w]X�eE���`D`��r)`������j��)V�/+���>t�>Qi��L���P���J4������)������12�[Z{n�	�B����;�K��"�<kۺ���\o	�f���� ��4=���q����o�=��<����j�S��	��}���̡M;��q�����]ٖX��Jgk��05I`ZykH�[�=��������ɭW��g�vb�	=K=�aq#����zY��G+�sù�1C���O#��t^b��j�	�����rBw��5��/�}:�X�Wl��E����J��\��Y��F4��Z�'V\%���y�J�L��W$�-���y����ܝL/2/g�5[�;���¥f;g�43�'�Y�̵�����ɎN�#�jR-|�-)o]��!�E�'��D��D�0���1��UҫR�XD�}e��68�����Hm�O �}��o�~{�L��l��✢�����-��i�T���cei)���[���?�1�{�4v���ӫ��Z�|� 8���絻�mC��|}f����g/D7{��H��۟O^^��E|Oemym��D�A&�A�oy}-N]�?͛OZ��jZ�n޺EF�!�|�9�X_�~Z]���MzEq�}~ƭr�Lb���㇯����=��H��UI�a�8�S��p�E��e5�g,YǮ�Ȧu� ���~�?��{'d�f]�ik�%����Y	��W���ZՉ(�{��0OCYD��8 �y��Y��9n]��L�
3��+�6�)���	a�m����>y>^`��qKͳ�q���`��䐩���<��Dh���;��n�e�ن�òY}7Eo��e�Y��VG�|=b<��:��g �0t�"��E��E��F�X�8�f�~�d/FN��4au��.ax���}�+W1�vO�@ȵ����q�h�4��;�o��锪H�0�2%ɒ��$4�	�y�fG\:7�U�����r6����t�i���w�*~�H	�V�/r ��w�p������P�d�ݾ���p������r�O��dפ��uӖߊ�O�������5e��fB�p��	���"�m"�F�y��*�/m<��fI*0"�Ts�寑��B�`�1�P�KXy�}���P�0�O#E0�/�ˡ.��g� �q�P�'�9�+����/��侱q��5�.���%
�1�� cQ�^�����+m�����!!Bh���Vl��6ǁ�,w�����Ŭ�,�m�nc�-0i�3|bZ.��n�&^S�'=������2*�bF�ҙ�S��X'�Y��[�,��h�f�cf����Yz�%��ys[�W��B2�6�0*��-�_<�8e�̢!D�M� Mq�H�i&�d�Z���]�pF�O�E�
�:��EN�����%ͩ^�Q� ���N��;};�U�D@�2���9�;�8%ɼ>i�.����*v��X+l�r�-7^n���1�V��֯d%J�59��WN�j$N	��+%R��oz�%6b�_�O����o(��L��^oKB��[������&@�o��T�֒P��%���B0���d|w
��
�Sl��$�������};t�f�jS֨b?�A�c�ڲJvV�D?�F	Ȕ�<H��m��&=�]~�v�ݽ ?�Ǵ������Ȇu��<ƺLB;��>�Q��I�S࿸rҩ��e2�=��B�0![#�͘/���WY1���r�C�[iD�$��Q?�B�ڹ�j�P>d�Џm���B�O+y�w%�.���K��馮��$s�G	�l�{��� g׾�V�^�i��d/5g��|T�w~�b��W7S�� ��	7���c�}�2����/�X�G系t��1;x'7�
r=�N���U}�����G��l��#��uC#7r��㱳�U�6:��s��|�2��ou넺 |��[��-W-�)�&�\�N	~ba�/"V(T�jQ)r_�*�s�T�QXE�J�v�DdJ�E9oy&��)�� �����l��H!1#M�P��tr>Њ�295�T2���ϯ��r\�����(���u�o���ټRhrT�Ќ������ �YF���"5L�ɵi�1�uH2tB���aL4��5����tk
'�q��w n�%���?��}�t��˶y��8I�H���_��ۼcip���~d�li�M�����'' �CD#)%{��
��>*?O�	H0��v;�Te1L"È�.ek�P�y��_j�Pv�`]ϒ���WM1�?\	�ufgb �`J臇d��q���vqP�K�P�hOF综�!}�K�(�m,�M��k�Mgڨ|��m�(i���Ϸ����R_����j����	޾�,�^J}�������5���U�:�+�M�k��A�5��~����@j6rß�L$�16�o��E˾���k�	Q]���E3l��닐�N�Sm�O���U?Y=1�-��Kt�V��c�4KX}�护��J1��sPg7�j����n�g�1?��N<����ֶiM��}0&1�q�6(~Jd����ط����9��)��8Ó�g8n\�N�#3�nqa��[K�V��vXhA��%��FK'u�ej_�
گ"k��+@�-ق]0��;�.��*NLB���SR�T#�WÃ<8�n���/��_�5]t���;�4
9�r���<�fV�#�����aH���ǔv��i�}ָ��0nM��U^�rVf�"DT��ĂqpV�_z��^��%���ʕ���ɽ;��	'��1ϗ�6@��F����ń>���GnѤ�p�!:\�d7��rT�/���ҤϨֵ�z��ࢄ#�دԓa�j�[�yfgW�xV�|N7��� ���h�a�a�$4)i<����}gj>��Z�&�՜Se?A�h!}X}�=�0��Y��(,.V%ǒ��R�[^�՛7p��%��r�������,���w�e?�ce�e��&�p��j�̰g�y�#vW�u"3�X�/r�pc�z}������Svsd c����U�ԫ����9_%Ϛ��|��RkQ�����( �72��Ez�|�_U���������F�M�}8��Ԍ��8�'���}mb�?4k���	hf��3ϣ���b�
uI���x�G���=��.�d����uAw�ȑ	n2��������O�r��0�oago��Z�u�*޼�K=�G�@���k�a1'}�'�<��E�w�z"`m�ˀp�V��Dq�ʝK��3��b*Y��)����,~*�o �O���In�f9�e��#䈓zݚ�~fw2E��x<��������g��_ݯ�F���U/+�RQ~S��hB�F2�W�K�#r�������S <�Ub�$d���l�Ve;��a��+���M��l�;�｡O�8�����������������ϧ;7�He��=gdv������C[�DDv1k_P��
d`�W0�����$8<,H���i��[{��b�M�k��j��4c�u��2�ך�̐7��?^Hª��<�w�,���Cf׏����(�m�\Č튂L~����\L�W��X�@G��hx�[|3(Y_����z�ȌNd�*��ܐ��.S�4R�8�q�}��ܸ���3�,w�T��?����� %g�%6����X/�v����%&7����K�g|��EN9D�H��i���9
�N����~+��
�0��J�Ӟ+�+���.i���NG§SQu#ē���2ua[Ȳ��yʐa%\���xiI`�1~P4:���̓J�F��Ϛׅ�٫M�m�n:��/N>�>ўJ�?a�t�؆�Ψ(@}�	�a�i���}d��;�U��O<�V���9W��䶊��LJ�i�1je��˓G��QE�ޱ"c|w��W����b���>"]h=��q�\��j����?�5k�Y�=>�ɶܳ8�����S��e����w�2����X�S*2��_��+4E_���w �p�\�t*��GP�V`<�и�$D
�p�i/�&��a$��BP�K���W۳U��ޓ䈚Q[��9�߮�L���f���rB�ēq��<��8[�MG����@�!r�W���pV}dn����D�yS���s�T,�d���N�§ᨀ>�O���ra�|����11�e��=��k��*˱�{2�`qC�vgP�� ��sw���X�ɾe�B
�nX���b��nv�¬}����[1K����>g�[Q�쇯y�z%�#��.�?bb���P��C��E~���br��cE��di��*ٛ�Ќ�i Z=7WY��]Ɲ��j�0��5 M�Jq�t.)%�H�;O��y9>Vh	5[v�U3J�b!\Mމ8k/6��ء[1��%�B��ֶ|x��8�\_�T���mx�����|Cv�D�c.\Y�H�^īkW�2��T�sI�tr�O&Ja2ή���7���鏉��y��$/׌��{�s�}\�W��-p�	��v?W�W���Ͱ_�j0�+5{X;��X�UG��� ��-p"%B%]����-̋w|�2�`��<j�pF�+�֕s_����Ņ ���ľ�D?�؀X����y�2�*w4y��`S���!�fߨ��bb��	�Թ��݁j&��yj�2TZ�s>�E%̨��Փn-ċa����*�B�=��=��P\�1�orP�è�m!�9A�	ΰY .���㯉�X�*:�̛�����Q�DE����/�[��-�WȓW�$��c)@ �a�T�Rp+�CLˎa�O0o^\T)#����CF��X���+E5G�����SS�I&*���Cw��;W #�i¥��6!\0ܹZ�N���$���Ơ��*�|�3���5�R�r��t�@(���}��ɠ?������}Bش��FE *N��m�5ZF���Ci�6�*���� �M�P�O6�-W%W2�"fb�\u�| ��;w�u��g�2�]��Y�
P�T�Ҙ�֒����n��jb넴[~�ޞ�x<J7�T{�RHq7
C�y<D<���"������ç�N�����أl�D��QLB����%ꂪ���n�0�6�j��_l*ԇ0�*��e��I=����M,V�:����U�\8Q��kL��_�����F^��{����7�L�p��b�q�$o_E�"���y�Z��E��x�yb#7_��mn�W�]�����9���b��~���,п=�L]2ޱ�����%��',���J�V�F�r�%1L5|C��g�,�v��o��G��bCjfJ�x��}n�tkH�Z�p��u<e"�#�E_SɭA�ܓ։�N)���,pz�;�h���]�(�?������0�����B�te�
1���s�豓��"�*�z@֖|UTҵL�0_��)���əqI#��_P�S��N[��ҩ�fG���|9�^M�����P2g��V�e�tw�dn�I�2��M��9��/Sw��G<�>�X�"|��7���wVleW��cx�*f���r¶yf��$��=���;5��:�4����A������_��%2/Y�I!/k���g/4���?i9�8���jSA��<��NxAU�����\v���o|)�j���`/^��e�k���_�;|;ґ�h�0ߪ
���z��^�y~��� �J0xqQ�W�380���B��@��<R�2�8N���2R
5 0��uab��zz�5S�8Z�I5P����CnUǈ`��b�]<��@~�Z�ŷ[z��p�N���˾�$�O�E�/��|�?���I��ɹ�P�7�A^Mp��y��9��d�P6��4�9���.��įx���ǻ]C�Q�q[{��!���IR��)�P��K�x~�%�oę[,c�����T3hWa}�;����#�Igڹl|���H�ߏ�ɵ�
y���Ќх{�ฌ��F��kB+3l���>�#J��~��<�j�8BhA6<mKHˣr����S��	��Ҭ[�s�p�HB��iN�@�3~ь^h���k�+�l�[ڡ?y�q��EK%��_a�a@	�`C)�}4�P�W@sP6�@���.����0!�4�ui�@�r��m�j?���>oaaЭ���
P�K��H�]�*����$Nb<��ל;���S)fM;�l�YDCʢEޚ�F�y��T3{O�|5
���]�x�Y���e�奇t��;#q0yO4W� �t�ldkO@����+g�����ch���xa���� ���7;J�sl�x���_�m�
�Ҭ�d�:��)7�a\bO��F�2�w�:yX��H���r�������$�U�u��Do���d���ñؽ�z�F��64���6^G%U��6I��0�~���t$~��#m�݌�*�3�0ް�B!G���~��z���%.`5n9S����lQ[Z�F.�{��^�{#G�/t�c��҃o@���|-�ݚ��l" ��O�5L� ���0�QS�HQ�I�p��Ϫ�خ�Fp!�D!ZNŰ����{cR�=�]cvv�w�n{��);>��<V�3f��
h��w�}��s;�;��6&�2�\�J^Q�Avr�\m�y��{�N��g[?l��ʎ�x�:�7�_���ۥ�Ќq�k��K�Ϯ�?|���ɷ`��#l��ù��"��n[�T��'�`xy�r���,������W���ssv?:g��E�A+���I��������Z������r�Xw��f�1.I�؄Hμ�u����p4Ai!Yi!�1��]���Z��������u�������9� ���1s�ʿ��-rv��S���*껅����%�3ܺf����d������w�n��ùӥ�6v����иפ��v(+WJ���8�-x��B�6�RG�X���Ќ=4&Ո�pv�]�򗻊����R0���.U��01s�XG�������py��/A �t�.�k0=���5MI:H��0�~i�Њ���y��x/n6�ܰ\���W/˝aͿ��x�g��Wz���% ����z�)�@�ӿmg5�j$�٦� W����G�Pʚ<�P���.˲:nq7AX5c�,��ks�	32J��m�Dp|���[reEo|~�h����Ѹ��C��0��{@r�3�us�ސ"�6���G��R�k��C�ΰ�'>�j῏���6��Mx�v����ȟ!�1��@K����RHЦN��]�/7ļЅ�k�2�bgWU^���ԡ�o�+��t|�0�!���[@U��d��I�X�[�s���A�7ee��݈�9�gOU<��;����Ƃ����c��[��2��x-���K�J�zt���e���m dF�8v�O�TR6�đ:��;�1�ϔU/7�B�o�9X0�E������n��lL��B�(-{2�c���%��@�W��10Ψ���^kvy�q�E�.|���ؤoRh�Y�e)ww1Ŕ�˜�S�J�f�kRY�@^��)�MSZ����H�+���$����:*���d1�R�Do��q,��kE�����@I�o��D:����!: w4У�� �E3G�ۮ�1�.e��Kh��`���a��S��\�4�8T��;��<����<����>��T��ާI3X��Q{Q�xT�#}#��\�!��w�C��/y���Y�E�u�U~ä����n�6��ֹW{==�c��pBQ0���1xo�+g����P��L�����}�+�^�.��taey}�;����-�7^�{ߌ$�Vi`0�z�ˇ���[H�m�7�>�I�D�I��ҷ��%r�6-�w+����!f
��2���1<+������e�Y��� �][����K�Wjb�� �Z�Z6x�9����/����2��K��6mM����Fș{<E��̂���K����vЩª��B�.T���TU�m�o����@�s��t9{l�EJH}�݇���n�&f#PP^��F�����ݓ���m~ ױ�@X-?�8u�<j:h�7ӡ���=#1!ִ������r���ϰ �[�ʩ���L��e��KP�E��:����uvЫtb��q���:��'�hYL�!-�X�({Z� /��y8S)�����8jVwB١v/��j5����b�(��tD~	��e\�z����B����jYF����j9����<����#�!%d�İ���+�r�:V���ހlf3
F̥�j����� #��@{�9����lj�fŒRf9�Z����q�!��!��6!]�wb@�vA��4��Q�@�G�!��z�@�g�P(��gK�v"�<V�������˅�̍���R7_��X�;>��L�D�
*�S������.	p9o�+V5��{�&Y�@�|�.��V�`-��#����B��0x��AH0w[I���?��%/,t߫��>�o��Jf���,�Y��	��!�gH�d1{@%j ~�'� ��N=J��,��]}���Q�hzupo��mGJ�֚6.���e!J�&5YS�����4�,c�tSK�Z��^m��%Ԍ:�-c&���|���N	�S�O�~���Wv�^�(R���y�3���l`���y.wNy��ϥ��*��s�G��I+��>2��ܝ���},�?���_oX_P�Sq��(/���	���J;�i22�h.���FMR�]&���*U�T�T�J�퀴-W��W�����e|m�̤7t���mE6(�SRd+lb�3NRk�\E�j/V`4}���yulp�|���WA�mK�;k)�����"&� �l��,�f�t����� ^�s�PDp�D	��T`hM�&mp���n�F��#����!s�j%%�����Eڪ1��%���ֆT#����Ȇ>�X.�S,6�lI�q<�o�2Xz�(���
�g�`���<�
��/5�[y�B�8o9c�w�˝�\�\"�;�Kr�-�ՙ+5d�ac���{�U`���jþ)g��x���J�&�<Pe��8�Uցݿ�?�G���,�/��^��J�O��n:�/r�]jd!��_���9��
�H���W[�!+��E�/�g:΄������C��m?���ؗ�ˌ�l�W�6�j�q5|�����Zu���P�هe&�j���dk�K�O9f�W�������!KX�J��4��{9&w~�,��*����H�[Xz�����)��@ޗ��-��65E���L�ӛi8c�iA�~@�����;jl��|f%_t	�+8�����w��s�WF ��kw0�.�Y�߻1!�m6��7fS�Ў"�>����:E�[\���|��-ēf�f6R�R}���ͷ�F�QE��A|�Y"w��O-pN>�gHm�;��40��x�Ӆ�G6'���	٭�c���6G�fv#ͮ,�_�Ϻ�M���0����/� h�ΙJU7�,���Ak�������<�Ut!u�P5�v|M���w�hϽ�ߓ�E�܀ ���{�>����'�]��G;鬲�]_)*�E\;�5��9|@�=sѰ�m<�ou���;�j��#���Z�>�]��2��`:z�ײ�W�����:�d��T�n 8�EE^F��^�j��� ' �p���|�3����>z���?�g�{vr��g�����}$Zη�N��~��oy�}�-{��QC�_�;Ě�Bhso	�Kz򊘦������]2`Z�g��Ϊ�:����ɐ断,��;���yoDZN�h��>�X��ԐHYz)�zBҸ�0��m1�.Tŵ�O}D�dK�������^4��NC��X�1��[4��ˀ�y��m�憌޺xG�?���*�l�?PCC& �i�Q�c��栙Z����*��V�x��%T^�hs���b��پ������,�׀*ѵ���|5 z�� Mz���d�u�Q�,�r��b�ю�
�����i2ސ~n��d�F��_��Fq�=4�U%�xAUf&�#�'��TV�[y[��ˋ_`宜!]�F�?گ�W��j��Id�&Ot��}��ꂈjM�<ŖGC[@����K �A@?v��r�bYh��Ddo�m�ktOet�m+W'j��$y��uSh[~���_���9����𰢱���U�^D�8�T�MbdJuY͍��eK@\\p�anN��x"�y�HJ�Q���5�SS���Z�?�ɗ��^y�<����29���!��Aࢋ�M��C�J�3��)"��>�8���*j��oI.�q�uβMs�3�F ��3��[OZ�5	5b�Wɾ12�
CC{ �a�bK�{a"yo3���/����?[��o�[���c<E�~��)�QΡ}��w��>2��@���0�+����s��e"
)������8N��FC�,,��]:~�l(Y|�����/|5Nf��Z��Î<��gR����z[e�k��0I�Ղ��X�بʇ�, +�q2��������R��kB9������Ϊ\b���Dʺh���E�A�Ke�{'אw�Y�Wߝ������׋��cs�����22uaZ���ں�З~	���v�5|�T#~�M�+���F�M��^����[[����A�f�����֝Ҙ�¹�G��֝���
���0ghxJbڏ"�n�u
�� g�eV��&>}a☛�k=(B��z���#}�r��p]�9����nm��d��A��q��V�<=B0���	mA�����b���T���XhŦ����P�Q��g���d;�e�+tm]M㠑'V�I��V�g�.R@$�˯	�$���V��,�/�d/,���p���ھͷ^-����=$��Ok���XH�H��O֓X0'Sm�֟|��O�Ξ�81�
�.�Ӟ>i(F-�V,Nn����?�c�"�byN(6���2�s`�v��:`�K���Fuӟe�m�A묚E�a��X@GJ�����B��e�E7,��t�T�Ƙ��>�?��d��W�l腫�����=�z�����yEt!�o�GJ���l 	2&~M��c� c0ѩsk9�E��J��M�o���U'ځ��П��J5	�c]C4������
�^�ϩ�����~���v�/�d�4qn�E��O�X�+~E�z	0�3ߋ1l<�7�LI"�:��S+ڟ�!��4��jӽR=Y|�Ӳ,��/�^�o���H�-k�~�y��a�����zZ6�?;��9��ůt��Yfy=���V]�;����>�`�<�U��;�{3�!��w�B�<wu؛�8W��~�����?dεSa(�p2N�4�x�d��������"�� ��Q[��T�}����gH�� �pu�c�aQ\��	τg_=����5�����	̍���h@"�3�F�3�Ը�L+yDrڇ����P��n��9}���EΫ$�(u�����j�{� ��E�}��?s�C_� b��@��7���J����O��R��1#sH>3��=��0�(���>�fq,��13�T �N������� #�'�CJ��&���.���0z��F~��}7ͼ��HE�ײ�Q��i�X`ܙF=�M�vw���B:?���W�P�ذOä�lx��<{�]x%I��H?����z�q�#I��q��U�ш{i�m����#�fC�Uh�W-��~YZ1��ף� �r�I�uDm�����5ts���MfH��ä��/�D�]�N��G��,��>t>&�GiF��D�i��2���p�5��t0ێ)���τn�;�&���#a���0��=a��Y�F�6���(���	��.Ҷ\�\���1��������dc���7諢ǣ����1"��8�̇��v0������!�T
L����-�Qj��o�4�r�F>1��(>���d��`�;��A���2�h9 �8/�s���ڐ�@�-�� ݚ��nj��m���_Q�[R �F'zʹd�U��L�hl4�]��3@(�xܬ���w[~6�/�f@�62B���-:Hi=�XhY���A���WH��>'%�`�Ow���H��ڹ;���yj��ޤ�6��V4ز�Bgo�r�GՉ��
ÀѴB���M��Y(y/{V�:��B������@�J7�-��� [~��G�������Q�i�>a�(�޿��sٙ�����
���A�qb��	�$%�]9�5��R�R�T8�,��	Zđ�����˙R��x�ӯ/��|樳�.we(�,~�<\�ٛ��/~d��$�uF,�I������2��w}gA���f[���Y5��;�|��A{���@�y��"?�^����S�*�	�� �'���L~�[��H�@M�WX���~��Y<7��N]'�Ҷd�	�w���jD�ޘ�)���j_��J�i�ٚ[Gkn4�z"��[X�@~@&�j��i�^~���줕�'��\FBc	�nƈGۂ�1C��N�[1�U�����^h�yf��1��R��e��$�r�+�����LQ�&ѹ��2}�/����*�f[�i"d�M��n�ŭ�d�*t�=��	ԋ�R�/�#��� z+�ӎ�D��ֱ��7	��m�0������� $'�d�=M4�b2��EB��۫����c�	�*�)�E��JE(pA,/�	a����WBb�6Y9��m_��K����U^6GK��u�����ӌ̡�t�#o��˙���SXu�l�WTM�ȭ������ݥ�.>ٹv�n[b?��t��n�xr�K��3������ʽ��K�t��3��ќ5y�Q~��J<�R�����&�#> �^*g�)�R_|v:�W��&1&���K��D�s$9e�}��Gd6�/��R%�cË.,��:!��	����z�������Z���66�b/�8����:�/��SqŻj4��5�`��
��J�@�D��(�(��x�	���m�\�fk��_��a��	��w<����G뼈IG�B��=>?`��̕/�	~~[������Ҕ��/�I�P�q�� �"��$�a�EW$l�s~gh���K��<���e�ئ^Y����[x/���eM;����V�΀8�寧�<w�G�Y$����1{nDL��n���r���b�r��<��kJ�����������6�2�)����*�yT$J^�/��?H8���lH����"��G�����Aѕi��w�����p��ٛ����/ZX�f&J�k�s�yH ���vdc�*�%_�t&�|u���v�Е��eK�tO���J��B�M�hHL:���6�ѡW$��CIF�:q(��]ٹpF�X����G��$˨̀��Fɔ���X�^�ڷ�O���w���|�cl_��u\���M�Zi+�0��9�5�����X�����o;e����`ϐW�w�X`!��8�N�֦.����[9�Vg5�/Sr�����U>=��p�+L��~ӗD�D��������q�ڛfYm�L��3��tBg]دF�N2Ç/o��Yt�'�K��6�+�~aۍA-	��#vQ��G#d"����k~��˳�+[#T>aa�^m̈́�Xh�v���������ѻ���h�Y���oGJ�o�>�8\<�����E���z���:}���y��J��b]]�7t�~j�uGd��j�f"�>����O���S�-���c���7!6W�/�M�M��.{.�Q�b��G���g��� �#��l�0�'o�l`�|Z>�Pz���|��s��T�6����#�u�i��t��9�4��m׌��c'� "z�c=�)�[hQ��M-S���Dӝ��go���5-K �Q�"#3(j���Ȇ��`�O��~bz�z!� ���T)�f�ӄ~��[x|���3�q�x��$а^_����N���o�J0^�V[�������}����8W''M5�g0�'�����1쏞)���I��q���<�w	�0P�SzY��2ޕ�([4�׸�^��n)vᓽ�Z�7�}p�ܶ�ïh�o��Ë�A������w�StfI	�Of�2W��G�j�E[cVsPG�����[J��3�{_�����R>s��ɋ:��eD���sg�)U���s�!˰�#ky����Y��<��~wۦ����y-�s4��s赤�_[�_M�~292>�7��0&��9��f�{�"�듳��L��[�p~n�����ǽ�x�[�W��)J�F�g��m��&�@���R����)�������6��^����ɷ$0{���"��- �/bk��lN����b��X�,�q�SZ{����]�Ǯ��WF�)I�u+�-q4�5ץo٧VF��s��Q���04����D���뇱X*�#9l���i�O���ܚ-<��Z��z4�����s�?ʀFb�8���//��3�,�g���
���.>Y�`�^ a�I��:C[�{��^#�h3O��ŧ�ج��O&�[z�<깾�]#=��l����u�/��[��X���!���!�}�>�)��)�8�Tc�b�����b�(�����A.d{$��|���JaDCf��Ë��3&9k}��\��t���f�}y,42"O&0yC��B�[F���&���K��[I�gYL��_����_�֙�W�9�6�^�s#���<����R7%QD��T���t��Pd�I�����f+�)R1D$;ٷ�dϖ쳐}��3f��<�������_�y�s^�9�y�\!B�v(�Ζ�6�vWK��ԁɞ�
�1�O�wMk\ׅ��4O�Z�/,_(�в��,VR��ϧ��^���O��~����B����#�� k���ɳ��XD>�=�?�rsJ{.)=a7�R���8�X���j�l QC����R)�R ��u�iT�����DXYRT���;�_��F�ޅ�;�������7���\j����U�r|�-�f�#�_w�h	<�f%mRa�+c��SJ�/�����I��}�`��/Q �^���b����J�T�" X֕`^�ew���)[s��:ߖ���/�ǃ�<�vrO����:�� �'����3^Z�1
�E�����mmǂV_6����\��j|���yU���PoC���:�)A�� ����V��)!����$>���5�yWfϾ�c�,>�x]�t��@O���3 �� !��\��2��7S�j�d�Y>��S�D_Es���	���=%u�G��Yo�:������M♜�֖s{���%=?��R��E ĉ]���'���s7�x2`����&Dc�����a�"�$A+�m�]��<Z�}�as�6[h6)\�+�NM'�����\�@ᦕ<��^�T����Pgq��H�Y���/�3me�9��ub����;t1RY�4�{7�����bE,��n/~���!���!�9�#�4�h�����V�#��!\ߡ�ǲ\�&0of:6+�Q���J	b6����U��v�i�������+�)UN�i�\1�vR(��O�.`[E�/�$���s���jȲS{u��ԿQ�Β1���n�CA����|z�O��Ȅ�r�Nq<�L������P� �ݺ��(��u�y%, ij(��g��H�}��0N�l;��3���b�2nh:+� ���W���f~y˅�}�kr;�d�
�� C�ꌸ��f��8�L�~��ވ#��5�zՎk|�9 �Y��4��G�	�-I��BÒ�J�ф�3PU��c����'�$f_�=�.zD�B��a'W^�������v��̔�d���3r��uG&��Bֳh�D8AŒv�7��b�B�Xc��Oh(� �q�zz�_�X�� ��O*80�~4�ҮV[���D2�n�#�gD�|q�< G������.�\>03�Ȩԉp�ǲ�s@'q��Q�3h�����G�6�=�Z*��ʚ8��B��&�4T�;�[�8�м��ͧ���ȱ�c3{�UX�O�m�x�R��/@��{�[4���S������;�摪��G)�/�$�5��J�l⏠T�k�&o���c74���V��罹��U��t
���ૻ��5�IT���d+�ѫ	=�jn]�U�e.�r�2�����%����i�O�����ms� l����?�7ڲ�X�'K�>��W�{)�Dv��)u3P���^�A��Dh �c�����?Z��;����}���r�@y��X�&?ي�
WE��7hrİx����%��S���n����i],0�4X�t��re�i嚫��ָD��ʕX{��95�*�H�Ɛ�h�dO{���^��5�ĳ�����;9Q?�W>��*Ί�l��2��IE�8y:�M��Q�jU��������I�y�<���zX\�b;)�]^�;��b:�|V�%h���@�g={z�}�/�C�c,�����g��Qaw�" e��5{��͛�I��S���B����HɛN%UK4�@�����AO/ru9f"2�ψ2�}g�
��h�n�<l��N<�>�K�I_2X2�J�F�T���@�W�:U�$9ܪ�M��4���y�����U2��	��H�}d[�A�蟾�͹2b�%�.�������!���!�=�P���P��2}>(�ZM�\4@�����}��k�Ϩ���&t�o[����SL�h�%��Q��W)	41���ݳD��%	[〉1�I&:+�O�	�{(��X�33<��`�I8�Yx���R���0
!��pQURĐ��f6%s�h��@R<��b�P���_����;<�1��|��o��^��z�w�F+B����~^�f�'�Qi�����(���o��Wt�"��N�
p�e�\��������u]�v����ɋ;�r��t�{�#��r
b���a<�.ݩƹ&��<LDl���3#�Q�����e�I@veʒb*ǁƏOF��Z�t=�ƥL�_GEs4�k��]H��Ǵ���9ݯ�1	)���}P��9�V�|�`�Pm��vS�#����@�N�!�yH��Oם��7��/� +���㶬|�}p��
�5�WF���mg�J��R6hIH�����8֓����yqu]`D쇚xgD�z�64.AE��,8����3P2�;IX�����;[��:�	̦�@��v?&�~>�vKxD�8����=aA��Cm�� �'����]-ڸE�q���"sA�Z���g��V�cv���O���s{��I?H���'��82�2��~o牍Ev��VwmҥA"�)ԣVJk���Q���g��c�ܐ�B������I��=S�C���@��c������q|��J���z��n��zG�'ڻi=�q{� !^�B�j����՝x�u��ߴϔLp?Q���r���d��;7��n����s����:	�1�	(2�'�E�O�?����7�:��uQG�y&Y@���]��F��+�ю��t'~��f6��SR �[� x���;��x�$[ڝ.��͙��!Y�(ǔؼ��;�,)@V`7�O|�]m�ub�'f�)������'ߙ����� ]�����U�X�����
k�M5�wz�xh8��v(�r�=�p3��W����`]�@��:���KxW�zu����q�@�2����Fj��}���GP�
i#ϴF}l�t�:d�{��� ��PR��/@��ˑC�I˄$w>��"�
��&���xu�������<T���6�~�l\j�����v���������7<�.5f�)��c���/�͸O5��	\y�V����4��5_E@h�W�G��=�ȯ��gc�AP׈��"?��Z2}ZΏ#��4e�td�С@�f3@˒���*в٤?L���?U���s[%���l��\)�˨M��g�&7��*)���t���o:J|����A�D���qj���`L���4&���J+/�9A���`�%�e'`e9*�i���։��NH�\�\�W"�iӬ+΁[@��[�iY}}
;����� ~>����W]z�4�p�2�؄��C�:�����=�W��Zn���,J�]��W�������Tt�v6�#$�.a���/��r:���jպ?"l>{/EL
�AK��\АR���%@��k� PC ?��`e�n�PE�.B;���>*i�G��7����P�@�6�j�A}��;\�xq�r�_*MW]v�j�ȟ�g	fF��?��|L����ߠ �.���5���V4�^��u$N�MM(I@>q(�x�d�P<Ю�ϛ�so�U�ۖM���l�qM_e	�g�XL��q�*H,���=��ϣ.���B���:T-���<�pj�*D x^�79�χ�ε��W7�k_Z��n�1$�pRjS$�� ��oau�w��P�|����n���*��ó�8����B�4��i1�{���o�B��}~�Wܥ���������**�6�	�o�a�9,�zZu8�:F�u:���>h����]�\��O�Yih�4RZ���S���S��,ޘ�/���>,|�6@��ɋ�c�p����=�x=�;@�����3�|�=3��랠V��{���������0
n�x�
��
�e�"[_�������%���ߢ*-l,��@u�������(�=�2�a����[��6vhxh�P��p�q��CRC�2��#7DN���E�QV��o�����x����l�C�W���"d���@�9�ㆁA3�2��4���y^��@tG��H��'���C��@#}6�T2jt�mh�МS�O!C��޷�,��ing[`k��Gj~/�	�[�$Xs�|��x)��c=�GB$*�hX��ѱ������lE�����q�@�b�wVs�^O����"P�}A�)��3��;Ra9���w��1ͷ�T=��A����n�j����\e���Es�
�ҽ>��6���?�0�p�?�6�>�j¸�r�H���S��j��rF���@`�77���V�l�-�+h�إWdj���6� ���a�%� �%�i1�$��nJ�',OO ۺv�� 6� ��#�_�{F���ފ��y`��fOA�ٔ���Cf����fx�,�Xu��)���v� ֍��z�x��̙�[��[��VwS�_"�i/$5PG����7�Ҋ�P����f@ӀŦ�C�P�����T�҇����Y��)%��-�˵���v��R.�O�a�ˆg�tj��DJ}H0Nk</NI9�a���'�h�6@�a��xQ���)�$^���
��:�?��[�!0�����\Qg4�CX�
���x���
��y
����p�o�$ӻ��0�ة��p{/3A��������.����--��w��u'Bu*��5Җ�m�� }��kio�]��ʺ~��0U/r��(2\pPzA|������){������<��d/!S�tС�Cm���$
���ܣ���!v��f�#Ûo����M�����e�4�\{ �A�)�����}�P���T! �9��J���OEG�ʭv�;ϳ��k'5�9�1�+�D�a��C���&�	4j$|b\IK�8���y�Ԅ���)t׭��!R�7t�c��O51o�l ����3߻�P����G�42|�ye3��@�1ʽb���(vK5	m~[Oc�"٨���[#��D*J �"�h$��Q��l� �U
��Khxp�'��4��T�{�v�o�X@��Z1�F5��l{���	�g�3a���k��C>��5�Ng���&��i����ģ����+�@�GH�Ym��jt�$��*u'��t�> ��h��m^|JשCٽ n�*#G�\_X���ɝ�(�8O�Q���`�Q�X�a���|�-q:�ku(��������~���/,��=j����Q��Ts�L�aef��d�;Xל�g��yE��+�SE�sV���do`=#u[l{��r�~6?�u��`�8L�>}M;��7��_�Q��y51�?qX���*��A�B����!�S܁�v!�jx�h�m�2�;�l��x ^ �6| 9����x6�p�����@�R�٢�w�:Ō{�pK���4�ԂO����R��ii?o�;�L��CxO���o(��S��H��&AǱg�3�w��eMI�O	�k��$���O�I#���f�	�s3�NU���3a�"
�sr�qU�oKܴZ4s����_��6��n�c!����������4�V�}�k�F	6Rq��Q�8���J����~��O6��� �~EF螸��>�D��+�吐AeTq0��FX��
5g>֞b��i�f�ii�5�II�E����.����9]��&�0�;���(�G�oB.���C��\�+z��w�tL�G雧%?w��}�7�E�n��Z�fc�������CQ<b�Źs��5�;Q���)���-��J68�O�]�f�E.�U�ᛣa�a�}����R��\��I��YS�U��߆��ޔ�U �䴒2�\���VٟQ���
����Bl&��Il�w�݅
���JI����}O�O�jQ��G�%������=g��~�JpRA�L�i3�N�M,U�Q��/�\�ov�t�hfS�C,�����[%�TnUE���p�u�m�O.��s�]Y^�ڼZg�)����V�>I�]�7G4�F��P�����A��oÆ�p�����C;�.���T��x�|I��ν6p4pA` �>8`�m����!�.�,ՊE��9<�� �Q�M ��\�I�W�q�$}��;n/��	�"�|�e��2c/�CYo�����uN�,TO[�^\�S�\�}E
�u\%���^�.ª�M껨�Φ_.�*jF�P��/� ���C����$W�N����YH���>�\Kc��a�V;5���\�5��0�����X����������chj��E�6�N܋ E���Wp<��%�K8�3]��OKr�M�g��T�����"FK�w���Iqmsu���n�8�\Qš�-<b7ƃ`�K`�̙����Z�Z=�����U��u�F� Θ�#b}�KLY��±�/J�nH�և��}��[&�w�+G:q�%-j��B�	.�1_����6U��s�}X��ϟ��ș�Z�������sm��#�J��iH�֖2�4�<ɫ��ˋT��ZG�PӆO�����A�t�:����� R��s�}�(�z��<ϗ� �y���%��@�7=��6$&�B�^C�2���������mJ��yLb�DQ��|���5r�?5��VT��}ec�)��,
�S��Q3?W?���͘��Ӕ�Ǌ�Fj�𲡋��l�����)r���b������5M��o����z��7H��ٝ:�AB�C���a���g��O��N��~����pY--��~K��G V�<4�j���7g�F�eZ�,z�� .��:\\�g����P���X�Gi�1^ЍƗW�L�������:P��]��!���2�����ȡ�<��=o�������5G��ҁ� �
y{�~��ҿ@讥����#,q��Q���4_T�!j�G:f[�/{�)��v�}Dc��1
G�����w�_�;����j
VB�5��HT�Q��1����^,-t4}���=�^�i'Xly[���ף�S�:��^P��������i��Tv g#ⅢNq��N�x�{n�!�d�;��?�c_��3��(�Vޅ�}ӊ�]I� }��M����`�+��2F1U�#Ԓ��5]M���~iE�K�p�J��<y1&<<q���!����O*\~n<3��~n-�m�3�,k�@�e���8��%�B�n���8��p���an�V��d�pš��c����q6q�4��	}��,殺�-�)�/�� ������߅�מ�M]��n7���W �i�4�:��RB�q�lK�·�Sb�}*�n]�Ib��0T輁a=[L9����h��fF�o��5���۾$L�=���S��<g��ؿ|W
1��΀3�%0�F�������G��V6:R]�w��\r��޿$����_���
3�A?&��EQ5�����>օt��ofF(�;؊�JԞ׊�sS[y�/���ˡ[�x`�~j�7T8xB�\���C��잜�0w�t�`��p7�]��*��O���&��O�u0�\7������PY��B�r>푁Q{}c7wA�.�4��!�������y����j+�h�۟x�s��|t�;+9pxc�,��T���� ���\�m�	��G8~'@2f���F�A^���4}�{���m�X�L\)��l�S�k־|
b~{;���/�c]8i�4���-�/�<�9��W���~A\X��ߎ�}��������6}�uzz��I>
em�L|�w'7P��;U�EV�-|�m��?`��A%��v����I�?H\`h��o�{�ݔ�V������{��|9�2���_�l�ՌT/g�-��6�o0@njC������F�`��No�kSU �������P�,���l�%jG,��[+����RkĒ,ga���!�������1���z�Kd�� �i��#�vS��P(������}N����Z |!�E��\���SI�k��|���?�)>H�4�"q�>/\����(��9(rthw�p��%Ay��y�W���ny?��&p(������+�׍�1�Ν�!Uf���g<R�h��	v����<"&M���?31�{��~I;�}�ѡ⧨��Kr�6I�0��q/����2�d�[]1YY��3�؁]ZDP�d~�6Ū�hN)K'�a[����
����V	��3n�JouTo�$::����N����5L'r��-�`�ڝsm:@ld��h�{I�"vJ?Z���m�DT�.,?
���_���/`�씦���o���, f�gg�y7���SF�j���*�l�r�66Phyf��5���<���@ø%�h�u~p���z�f�4P��?�c7X�e�|��CVw��G��O���+�y�?WȾޔ�]]��f��� ���F
0�1���z�:-j�����S�~�U�҆��/劃{� ֖X[�Lc�<�jb�s��FH��̿�/5�?��( Z��p��4���-���L�o��� ��"�?-Q�(y�����{�NXcunc��8������b�t��D
BHY'�PJ����߫9!k �m�Ԝs�%�q_�Wm*\�o�i'���7���
1��Loi��-M�����Z�t�Ȯ�2%t�J_ �%kذ���΋���G�.7��S�FV�\�`��׺�R��qM	�zI�қ���~�Mu\��~K&)Z�m�,-ψB�Ґ��R��_s�%���v���_�c�wX���q�i|J�r3�~f����D�r����l3	<�}�]u]MZV��h�����?�>#2��n)���$����5���į�{ye8�:/̳�3���t��ܻ�(�.T4�>2,�$�6�ͬ�w�#ߔ4��Υ���z���d������>�]��_s�3��� ��(Y}kJb�]�ߪ��N���L8���U�d�K��q^+�C7v�=\����^+l�X(n:�Ͷfw���+C3��\���]���߸,`������,Ҋ�!��WQ��B���G��c��=���Ш���ŷO.'/c�J7��Ԭ�������j��ԭ��R5m7A�>�@��M9����цjk]���N���W*aP��% S� �Nx ;�G�gw>�>����y�p{[�!���!��ပ�WOz,�(�T;
���vv���dI�V&"q9�86Um�թ�9�ϣ�O��y��j�R�w�A����_�w`�a��:���g�� �s�nx6����9���jF��l`�_)��
���\>�ߠݯzu���+
���=��j=��8jg@�Z�ۀ1��;����f=xD�CV�G��R}�1��oK����A^�ܷݔ������5f�f�~n(�`�kT�3ս�4l���vR�sX��/�i����<����Ԁ{����	6/�o�����2���,�țwhM�?��<�,�}��=�*�B�Nds����È��5� ?�N�l��ǑO���)l@1���/@�>/�E5��+�Q�ʬP]XO^��?�#�V�d���Ke��:�,@`�0b~Iخ7�[UrA{d~/Z�㋟��s�	�%��
�0� ���S���x;�����_��$���{&���r�|������z@�����^ؔ�{T�Ko���ʦ7�`�{{�}ox��ϡ��=�0�|���2�z��9�;q�_C��.��HZ�RU�X�v�IgU�؉_��	��i��������+=�?���Ud/΁G<�F�6��FJ�-��WR����?\�<�:A׷���6{�I��h��nOߺ�y�9�N�k��uv0����-C��^�2NXy���P�ls~�r���Oxx3���^p�����cl�d��<ĬeH|�V��0���=��	yX���!v�p*[]<��u(�=�����u�'p��%�o�Xko�q~N4����oI�)�u��>o�����w��7/$毓j����!5-�+hP9�8���<�� 	�<����@�Ojy!��գ�Z�Fվ�ZZ{��0��]��YH�L4�K�+����)k�o9��Ԛ�h�;b	Ɏ9X��;8/4~5�����i����&�`9C��������YW>ffda�M���V�7I�`1�H	�x��	c��� �!����	��?g�֮.��h����h�,��z��{&�͌/8	�y:]�3W�`��GwR��)gؼ��:�b���GdG6�$��1u��jR�7�-�X� �rk�iŀo�kt Ӳ@��OS�-~Ҥ����rZ�2�]w�f^@�E�!�^q@@>��}.�It����ԝPT������@�M��/K�V�2J��s݇=�cN|�́t�7]�U��n���:��إ�}�rn����0�qm����=@�i���z�QV�� ,�i���R��r�d"�8J�*�x�.sDR�hŤ�a��;8x\�'���8��>wWm�Dy�R�&��|c?!�,�Mn������E�ض�`����b�-L�
uq�z����g��)a3���UZ�=(x�g-���u�x�)n��D�I2���}�4�[������y�?�ȋC�>\
C��g8����,W
>�t� ݩϬ���~2@�<�&vX�Tf�^��N�`�@�d�
$[�����s�X� ��;v�=�s^�#�+$��G��\�U@M[�B��1��� ƅL���&�%ʐ�g���d��c�o��P�2;k��'8�G�+���]��T��)��n9��ڐ����[3Q��,����0l*\Adb����h���5��[N��|��SC!�8���V�/��Xx�����'ކ��/�U�2'���2����~��AeL�R���/��}վ2�����@!��z�૩���9P.��j�#���*��������j��lۍ'�Ȟ^���ʃ������d5ۅ�/��̦mg�+:��~�y�S|��=*.�FM묖����,��!��������M�Z�唭�ޱ��g�J�~eۅ��̥x`R�J̡����:%��s��1w��؅p�e�}[����p��{���@MM���D_cM����#�$�M%��ʲo�m�L�uA0p��m������c|7��<�\���r򞩮]�b��$6��ۢ
�����ZuSqzr�Y��	�A��W{K ����լ���sx�1 z�ǫ�������I!��7�/0�*�ت��mguϻ8[}K�L����O
�<ɟ��I�n�aU.�s�$����m�z���ک�����:�q_J��̗��8�����<�?l��g�a6��Wj	��7�'���z�謵�V܅��>�;��n�Ĕ�����{e�$��c�K'((�ɢ������m�*�և�c�2G8�}:���H2-�H���.nj����ܙ��Ofo�]Z�b {�[Jr͓sjK��"��׮�O|#bE����e���]���]�=���B�	�0��$�J����Y�����̙�j�c�X�aN��yX�=�A�p0��z:O&�mr�z�]��kewi����-z�Y�=绹1g\l�v1��*U�J*��d~r��\�����]��|J�Ne%�k3-�T����t?�և��-�˙�1m�u(4.�C���f!IQ�4�N���~;H���no�0�/f�l�t�n*d!W���OR��eYq15�~~]��V{��y�,�Wȷ����6��w���=|h���V��B��Q�D��[�c���$m�*(���i���5tG��ť'퇻���b�\�:ۥ��$�$���>���]l�R� C���P�#;zf�`j�@�K�J����$v(P�Ӥ�ec��M�X�,�}X�)@���V��*�����}���<���I�K�QUxj���=b1 �R܇>RO�������	~$�"�=o�CT���F����� �����}�������n� �U�� ����4P��<�H�C��|J�E��z��;��dq�Q'�P>�a�q����&b���ߺ��m�>� �T��r�YZ7�_��c���ɀesaiKX*�Z�2�W��\<X�K�|�[5��hA�kHp�4Λ[�ٙ\����K�~4>w�Uv�^��0�Գ'�X��c�p��GA��H5���G��ځ&�h�s^�\�G�1m!� Q��j�u�%u�f���yi��H�EV�~h�q�8X����X�؈�fpH��u-�|5��+���nP(T�T[y�cxqG����ωS�^-W4FJpc7�9�1�����xu��Ǌҙ6��G�p�T�a���9X�W{���$����vo�zs�zx����)P a�έAC���+�@b��F�i����y��w 2��K��z�D� =WE@l���#���4pe���
�P$% �F ����;��p�e��ʓ6��;V"{;1W0����$&Fzk��Ĭ���o<���e�`�򱂑�:��&�p}[/��Sbsn�4�u̐���EFH5Q"T�N؅���3�?�Qcl���A'Xt��H��$kV��"U�G����W���ݼ{v`�R8(lŭ3��%c$��eH�P��x�`{��λ|�H3MJ�=�~�.\t����R�e4�4��e
1T=�����i�B�[�E���e:�1��H�ȟ����Lq�upR�-!�<x޻��x�����U�w�<`Y�����!5�vCx+.�I�_�����̈� � ~ǭ��ndg��^EV8�͘V�T�~���)<Pq��p1���c�|qO��A�?�A����[�ŭ��T��Y���I���K5ȴ7�_��C'6��^ޘj	�Ul��[S�T0&h�=�U���0?��,[�6�/��H����1��/N%��s+�~Ni�W������X��7�U���Ej~oZ�P��Ф��,��b#�(�q� �s���ã+32��>��قe�Q�į{����w�ݑ�o��#'Z.��~��Jh�R��̓:yӫ_�4u�ټHÕ�e�MU�'ͼMR�Ԓ�0�rGT֧ߺ���1�K�-�R�ܼP����.�F�ĭEZԱ�[�ל����q�W���}�OY�Y�H�6�I.�>���#}_+!��^�W��E�qq����L>V��_<"��J���?w������+�x��i}�sP�i<�'ȟ����������.9���iC�>"��[�ދZ��X\�+���?���0:�#@I��;�f�X�Ԯ�a�r&Nkɷ��F�D{Ֆ�na�ar�WP�X,�JT�顰�Y�) ;�8�crz�H�J������y������XHQ������20�1&�3��v��H�Ģ���O��@ 䧀Tqة}+�բ�3ϖ�ze� Ӗ*i�/��e���c/I�)Vg�&��L���Rvj"�� 0�Ƚ =Ǚh�����V��jP�QWY�	3��Ϛ]Z�g�����;ws^B�)J�gʕ�v�К�{���u�',h=Gm�״bG�RY2�+�]p�3eGg�J����}|��7m���gGͧ���ڝK�ؙ�o�%�
���fI 3��9�P�p�� 5�9a�T�����%�߭�~����y��Ì
j�e����zo������xN��tU�!���	z�B"���z�䴖��DX��>=�I�����s��02����ٿƁ:�����#da�ջ��S׻	o�,_!���j}z4)i 4�<��>Rei��2	F9���L����)m3&�=��vsP=9�]���d�\�6pO�L�g*aݿ�J�&�J?����D�x��Z��d��Y�b#q��
�L�������54��uv�^jSjb5�)!�*8u����de�M��L�痊NQ��8�T��J0*>t�����;y����Y�RF��&&���������{S3C�7	��N�}Փ Cl����!�w������D��⭣s����w?�vŨ�p����_����=ѯqEANh��p�˘I�`Ԃt����Q�{�};���A/��5�eTBc�Ă�qk;T#'T+��ƶ����m��9١Jz��r�$�#��ܵ�ǎ��׸�?E���q^�j���,q���Y�?��c������@�P��i�vTݯ����]"�����R{���Hɒ0�y|2s���y3�TЩ����9�g�2�s�.1�?U!���o� �)S��9�GD��`Ǧ��Rgu�wl��ρ��-(�mw�����)��DP~J����h�c�3�U�L�{Փ�nhTK�q�K,��2˫Q��������c� p�[BŌ�o�D����%3Gʼ��Y˷�Fo�K� H�ޭ{�#4���D�vz���ըa���|ٜ��(�����JbC`ay��rL��(GB�>H�c�� �SV��U�R�
���ß'�Y<{����΀O���6&׻��Ӆ�Qbnb��w���,Nƅ98G����5��T� _?Y�9�qM��oٰ��R0W��VW7� H���RA�����o�S�~�Ο����g��x�^KY�����N��0�~h/����0¼�ْw���=����|uD�>�Ⴖ2T�&pQ�HJ�dt�T���)<e��b1V��u_8� A%�R�V�?��,~�v�#�pe<���Oʺ���/{�}}1�9���u��ֶbBf���3Y���bK#g�"�s�k4��o^�A� ���&�>:�=�	��U&X�����5c*�Veb�`	�Hڼ�K�n��@��|D��+�똑���������Zyy�t,�*U��p%���p?X�"?�(�?`M�A�~h�#���E�?X��LJ�MI��Jг|���JeA���Fb��|����6*�DNefż ^Y[ՁGc
��`��KV���,91�E0@0�]Æ�R�MU�H�|@��Eo��$��~g��}sp3�XY���kE��t�%o��	x4=�Z\�h����@���S�XK��^5���2j*Ɍ����С��_����B��!��J��D�n���@u!���Nּ9z|>���&M�u����0-}�����z���p�&��Z�P����*Լog��s��e6�\�����H]�CX�~�.��L����ȼ�g�n2�ﻖ�Qnh�Ժt&�.�qh5@ �_���Q4�����3Q�O��1�
����p#f㏹��\4��Tc%�0F�>�%�\�)YI��q�^[L��5�EG��֎���C�w�(��;Kl�����ɖ鷛�qo"����v
J�C���F.y?QB�X�^؎��:ή[`h����<4x�P�Φ�<&&�yI�[S��/aJo��OiE�QTb�L\V��{rG��|�����9�� �	4����vCW�J��,1�}�JUp{q�7�M�%�u��Ҏj��L���=�B��(���z9�y��{C�9�j)D�=��/m�F�G���/�;�x<����&���Į�I���lbQ�0�r�*Wŝ��<�\0��VX��Q��g9Ce�-
ì
m����T˄���FC����EZY@�����;+/�y(��N��&�&3d�8?�2�ȅ*�_��%�'N�	B4�|)� Ii��
;j��,��̨��}:�08��ܙޟ�7�G)��`jMll��'�[;��C�S&3U�;��n\��2�G�8+<����b>���4�j{�	�"�݊��37oٖ'j�C���^o�)���nb�Q���2(�����U6�W��e��i��89qF��I�5�E���.��P/=�P��Ul�x�J��t���hD�X�EN���>�ș���\�WXۇk�~:�{Zc����tC9c������K��5���N�C� �(:P8A���(�R~��	6��Oy!-�3�(����9#dB�F�D�v�s�`��A�Ml��VX�'~��F
N�D��M�����J�v��ES���/��z���EmpnмP��O�Xm/X��jd���MFKgv+Οiڛ�^K�N{\EӉ�*;5N��Ti_�d�
�E���ݜ�Z��>�\��=uP�Կ���f5�,<�K��q(���9�W��8'�*���{N;�>�wb��>�m�ρW�X�4�j��/��i�ݽ�$�V�k�j}�oʞ��n��WM�+��m�.M����V����@��4a�@�fv��6	���0��*��/�|��z��3���YCP�@h���]�cyd?�����;E��rA��3�E��1p���s�����G����� �'�L� ���j ����0�}�x�O��`I�����a�ʿw��B@�U�`�;��ԃL̘�z�����OT�d��%>2Y�m�>ۏ��h*"f\�����x�����5�GH�aS<��{˽��Qd�H[Ţj��OW	vU��������5z�o=&���:`�*�}5z���Z
삥r0W�0�l�D�I�*}�ueT��4��[mI;�	����Uʲ� �FT�(�a�G�iS+��_���! �Z��� )J�)�%?*
ީa��cX�D0��G��r��f��r�*x�&}�>��`ٺ(m��R����}8�`�O�`\��dSLn������pY�]9Q,P9�g�
��~Sy�ls�y����p؋�Ŏn� ���FhC�F$��433��cx|4���YY"��jq�L� 0��a?� _�V�>p���v��݋lv���d2/�����юq���Kb�a��>KܸƆ@-����~RZ����?��&x:I��F��5�^��ES<�|����Үt�:%������
�@�dEY��G���ܜ�]�U�k�p2�k���02��Srk�릢��!|��mYz ���M���Z>Y�jMd���2���L@-O5l|,?�P�G09HB���^�fب���ax�(ٌ�����Ոb��2I�G��ӨƉ��Y�ԁP~���e_Oz2��Ѐ����^�h���ˊ����Q�7jj�h'8C�7�h�������̼l�����٨�7��_�r]O|ǉw�w�*o�s����ߣ���3�4G�Ź��p[��?��g=��%i��Ě0��y����F��
&h=��`����g9��[P�����2N�Rn�	*�ʙ��f��	,F)�a>�XUg4[��PJշ���FY�qvX >#&VS����k��T�<�N�!��ɂ�y.�ubO6�P%:�A)&6���]y��. �}��q<��R�o-E���F���ҟ�>�F���<8|�7 7:9���o�ǰz�,W�ѹ�>k&mQe\J�ѝ��D�ЈcC���6TeL�'g�}[�(\	s�c��"Ȝ�����Uڒ�`��c�y��ʂ{r[t˥̾��&c` �VIL�x���Fh�������2�:m���q�N��R�Ȍ�^B5�1��E�G�~��&}�3��}����Wțe>�V�]��A�/���ˊT}R�J2Z�o��c����[SÏ�b=���=�
�~��}�,�z��f����i�CbnSw���S�������)�e���a��NZ�K�ϤI�E�ĉ�O�)�؊�2��� �xo&��Hހ�:�2���z�غD�lN�m���:,���l�2#R�C�eS�`�����WLJ�d]᫵[U��4i�����QQeY�p9N��"H�-((ݠ`�
J��A��`���%��((��
P�@@�H����
I%�P�(�=�ܺ83��������Y�캧�N�~�ާnյI8��!�A��J����"��~R1I�솜�w�|�b!�����L�D�t���z�L.=YW�3�|����q�O�B͚o{��J����y7ﲛeV��V�1��p�g���]�\[�u��l��jƝ��ؐ�"��>;��R��sb%P{;���6:@�D�>�*|v���Ws����|9�S�fBMz�
g͎������Ǐw����M�FȯKm}���ۙ����b<���[K�e~�l�@��MZ�[�R�B�`]�j�Ǩ�&���aA��5U����"�@o\r���'���|ˋ,_�9�/F@C'�:S��uG�������1�LT���/��б*���NN+�Ӛ��W/"b"L� �aP��Z*��ƀϘ�D��K��1>����m���_�o\��`�ᣩ��"Y��x5� ؄���j7��|��~R���rF�l���`�rwJٛu�)%�W�|fS��e긠M?R���+)\lST��v����xh��.�K��:�s�B'�x�����LVS�cL��|�#	�e�
��WfWz��ښ��di�}�Xaz��˸�AT�X����<\����xY@Y����.����+���f4��Dwd9{�����a����m���<��B�󄴧�gظ��+�/o���MԢs1����R�
�t��v�x��naU(�'#"9�3�=~u"����}#��CQ�C򩣔��"фn��ya_�Q�2�Ⴡ���"�!��:��z����+g롻��vY�J>���9[#$���}rB��}�E�n�F7&�;��+�<u�p�3t��z����%#���j�g�q�R�p�ͳ!�����k�/s��w5���n�io�'z���6���������5fg�К��慬�Z�{҅�4w���/��)�>n�D&�����kG^֏��,����poI�����M�v�?XM�r?��:����4j���jw3�m�m�qeN��zy�4F���U�"0?(���	�s�v<��,l�q 1�)HQ'ݬt}V�t�8�`Ej�_���	�yq�
Œ��= T������4<ߔ�E>+�e��5h:��j���."ty�k���{�qrs���'ݭ<]������0�),����gh�Qn��"
���zw�m��R[���F���*v��8��k������Gr^�D�ls
Wy��y��^Qp�cX�5h�c}�����p���u�����Y��;��9P(�/�)w*�G��1�'���f�H����8�kj��(���i��*�ӏ[z�DLz#4e#��S���@��Ͼ����:]c�Zg�h�0׾D�"�h��z��W��w���R4UN�)�1��i#���Ҁ������CEe��NJ;�0��A�6��E��zW>�\��Z�#mU�&�k��̳�v�fҳ��0^�p�q��lKp��9:���,ȭ8OH#Fπ��U�<㧥��a��S�^yu�F9�2���u�;��F�һۣ� �$6���������͍mor|�{�P�c��3��S��x�b.uc��~-�iq�]�Bd���]�����ՀJT�꼀���pM��pi�'�+/fl��}��l���� ���Qv��-�j�Y�(F�6x�Dz���!�	\��n[�ݓ�%�q=�B��Ḟa��_ ��nμ+^.7[����W�u?��c
�b���c%astPv�7�e��5UgT���'�����,�G���^�ͯϳ?}/�W�B	u�ݸ��M�~2�"�3���]�����	�>�+���sz~�*��2���+����1}:�N�䩛��YgX�̌�`�u�˼@&�{g?�0�����:7��A�Z���bwa2�E�B�ʂj������\��
�a�B�cF������=��=ν��Eh-�ܞ]��M8��t>h��ʼ�њ<��;>�|�X�T�f���h������`��~��צ�L��.�9my��5�'�֠����E�<k\(q�h������w��Jc��_`n��Z�)5['�>���¼�lwƳ�Z��2u����Y�~��1��=�S�ݒQ6�Q�{�0׵=�\'� �[�r<��-�F�5�o��f˟_|%P*���#O�P#����HѴ�ò�����wҰst�W�w�0�E�(�y�W��%�U?����J�Z�]��˅�.wݰ݋������)*�Z,M.|�����m�]��ȓV���*�!%�n
�
���s�P�HF�9>lwxc!�:,�v�}8{{q�FżZ��F��,� ?�L0�ȵ�҇���G�%N��8C���M]�Y�����\qo���8�r�u:���4����X���.�"�6 ���'΢-�����`�T�A M�~�z�U4o)U9���CP�$��3*Sx��YO6Ep����.���7�j�y:��U�+ZT��gTs��|	R�NNЉ�Ivr�є�ީ�4F���eV
�����C�
�%���u��z=^H����C�����Nkj�
����f��aa�g��`�܉�k��:Hq��5�mϰ���	��ڱ�	����!�X� ��:�x��@���ʹn�u4]l	r�xz���o�g��%cx;���.�(�NG�F@��������4�I��tIy�hW��`[>#l��@P#t��&;Y�
j�k�9ۍ��������Zt��`���k����:�D���m:Ʉ�*��̲7�d�6On�P����#T8`�L�j�P�V(�]�#��;�g��aq�SQ���7q;�I�����q\ͭ�Z�~`X>$���6!�m=5�_�2%u����znW����@��e����Z�_K����%�sD��Mn`5NF���I�*v�O���t����)O�z�η�/c�������8����5�������X��-�쇍i���u��M�8%��Ɋ������s<�Π��p�} �,� ��mU�Zâ�  5���6�V�5��("0nElJ���(b꾾�_[��Z���;�ɢR?�C`͡p�SC�92�&:N�D�Z)�,2�AL�b�k��Y0��4a����g�ݐ�5��o-$)�^�GjB�e��Nmw���%�-��IX�.�DL(e�~�����s
>d��&�m9�RpFG�ܼ���|'�iv�Q�B_��C��L�N�_OS�-p�zd������P��`{`�s1�4�9�Qǎ��Ԑ�t�#��c�GF�g'���gG�u��}�<���]^b�=�3��{�����[XwGYz��b/=���I/�t�䡝�"��L}���%i�ߔ}�����Pxw�}��^X����'��E-&C
Ղ5�܅�����dY���.������ݗ��^�oـi!�����Ӗ��\r�;��!.�0����f��|"h�k�����h����\��,s���:��n/vʱ<�k��X\c^6s�m�9��������sH¾��7<,~/�M�� B�ܘ;3�$~�z�M��?l�����;z@ӑ3J�l];Th�>xC#a��g�9�[`k�kZ�<ǹ�N+��}j����k��[���=�,�ry\}p���H���(c���Jx��y<d�wa��I��ɸC��]��Z��o+�ο4�y��d�<�Z{���t<�Nmi'�c	��GU]2�I��Ȥ�����}:�����sA�Ōk��W��Ż�"_|n�����X�6Ӻ�e)�*�
����^2a[�8�P�$E�kh͞}r��Ǚ|qqw��8�ӑ��oP�qz�u�&m�]��-�Ƙ����"��7���R�I�5���y�ft��ΡО���,v?�9Ğ����.�q:��1x�Ξ�/+�1�$@���}����ڧ�B8Xٱ��1�����A���z�`�t��}`�&����84zMa���p�h!�����@9^q��Y2���V���}�@��'4f��>o���@����^��#x2_�AN���RT�e�^4��7a�]i��i�C�{Dx2�|������U��z���	�N��,�N�4��	�:��9Y�umo�ƪ>�w?��	�v�}{j��1Z�!��ׯI�~��P�C��^
z9�|���������)�e.!J�i�)�G�ŉ�X �7* ��a֪ajA������U�<�џZ�߃�a���J�w���/�Ã���5��NKr�Y��>��]���AKz��W'+�Ѻ+;�����c�b��@�~��k�1q�(�|P���1b��'Z�k�:V�;�6������.7� �T.�\4Q"����	�)��J�� ���j��\����]Rh���KĜV���Q=۞�uKiK����D����`��B�=�$Y6�:�)���c>�s$*, ���@����C�[�kc9���3�zP?� ����>IX�Wj?{?3|�n���ʶ���I�D�����e�ƿ�����5
�u�t�;��Y8B�q��Z@;��_n�M�l�B;iHϛ6�g۫� �������S??�����Hf~������\G=���ю�b�)�耲�E_���?��d}i.o0~��C<�̀���s9�/�-����-��K�u��*(>ة�?���k�nv�@�ځ0��u7��p�F[n`������k�_ƃ^k{4.?o-������@����6�1um*�˫�_�M̹Г	S�؎<z��3���r�Z�5�·DLt�DT�꥟c^�i�=m)�"����>0���J,̕�a�+;�ڇ�k%5��M��( S2�����]b��.8����iv�+?�~��NKI���[��}�|-��P~���=������S=y�o�����<F;i!�����n���$dk�u�3w$x�/��Gئ�8��U%����؝f��������h A#2a�O�O�,����=my�����B���M�g�-�?��#-��F�fꎃ�9��3�𖻔=���1+��A8ᑠU7�(���=f��Vg��K2Js�;
>����:��EO����`�fm�vD�t���u��a����x+�iԎ�9)����՛ﻔ�n��0i\7=�$r� ��x8]��v�l�ů���DHw�c�Q*�VW�Xd�1h��s.�(8~�0�ԯM(�tK�Hn&�\Je�_̸�8v3/X��i�_V'ҫ���&	Y����6��ՎNWqe�:-[Kr��lC���#���U�;�:��\g6r���]�,��IX4Z�w�����3�g������Ŀ��{^�.����"�*����!�V�����ڜ��9�%����+�C��xv&�H������yq��\�e��n_�=���]+��6ފn��$k�̭��5L��={�����
�����on�O,�ۗ��O�,֍����w+����sRC��,T1����Gqe�P��ç��x��7�e�W�s�x𾯚$L�D���W������e":P��0_}t���Kk�c�VT�~%����[|+��*-0@O�2z�D�p����>�\���o^�Y�d��_�xsq����^��?[�Yӳ[���)R�������^����+�EG5�UJ�@O��@\]]�^�f�$'g�"��(���D��F���
��7'2c���O�N��{���+���y�����|&	o:��Gχ"6%h���7��]�ǁI���t�ʸ�s0���;�|]�eT]h�h���;0���|i���쎱��r��ݾ6[�������מ���ү��k��7?ؙ�^�zc��Μ���"��:�9V����M������کo�rq��f7븓��եz���~�����dwXk���èSB�)l�h9��a�3Jc�r
7���;�o��w�8������%�z���+{�'���C꩏/���$ǫ�����\+�} �x}:�n��i�?R����������È�=ն�J���ӣ~��Y�+�_��Ƹ�U_;`���.�Jѽ&���n5��U�Gf�,^��L0�5�
��)p]��1A%�+!���k�Y�����7�-�;-���Łm&����LwJC��[#[v����h�R@��߉���R�_��k��u(1�����m�Qe�A`�Wz��1!��U�o�?ޯk�dXx"t��wA�dc9}�A�{�S����@>��*��tDS��b��<e�ɇ�H�]�}[b����8^��op=��4�= �?�9[�b�W��e@�7j�	_,1���K&�9�J�n>�.��<������Q�m
emIl�\7�%�x���f���m�r���͋�*�\��jsk�4������Ot�V5�1,�;��o��x`�-$�/�Ә�F�P��b�7���&�e�%�ŧ>F1�J��,:w�<�O3�� �y�1YQޛ�T������݃�=ѡ���h��f���m�
���M��Z��G�D�ǻ�|W:���{<e`�o��֬��5Y�Mi�/�pe�oc|}}a�N�{��
w9�͢~�+��D|lՄ�hq����G�3�����vsxh=yS�{:�#!��^����vB��E�(����9�R%�����J&��zeG�{�E4+v�Z����;�W�9�>dg�4�˿��9Y��q��l|�N��A�����O*�_��Ϫ�M�Ay���Ŏ��iQ�Į��JW͐2_��D{��{������M�T`f��C��[�S��(���|�Z�r_l,�`�e��53��#W��ROR-���[�Jl<J!���7wl�p�/�n�{5���(�^>����!ioNJD�餢`E���2�՟l�3TD�>Jf��Z�8�#�R��5�4�����0�����'���i�����_���)M�l)������!�j6nes��s=Z��+�3���ٗg�Y�IP�/�y��ce��q���si�������d��RQWN���nU��]�e����¦�����	�����	
[P0���L[�~��	z�����������%wFR�,��Fʍ���O�Άv;1�<A����!=�ۂ�R�I�V�/$�RM��0�Z��^��a��?s�T�K�I�VL�ӑƮ�lf�/B�->�l�/��O�'وN�S�O��Z�N�tS��@��rK�IԣV#fN�L}�$�Q�o��8���yO;]s{�cE�y�X���Rp���rM:���]�n٧f���kb�_�pS�<����j�P~�;e`�3�5�r���V�|/`zG����ϾA=7?�()Y���{��.���[��ݯ���Ӿͫ�I����ܠ�F*���Ƈ&n/�L������Y��Φ�Vz฿�˂����b�b���F9�0��}��5�������Q
c��R�%��E��=��/�t�[�Z��z&L�μ��,�m�ut�>��K�E�9u5=�2C��Ç������Ǆ����
����?d��"�)���o}�_������Zh�������������D>����o"���&��o"���&��o"���&��o"���Md�F����W���[���(s�ƫ��n��s֫l��>�� �rY'�����Đ�z?����IOl�����e���������V����_��&��o�	�&��o�	�&��o�	�*��������o�	�&��c�jW.G|��W'����v�v�&�@�����v
�%�K�(E_&����wyU��k�\m���������(ܾ��8�형�lL�����MtK���/��p���{����ȣ�ˮ��𳔓�/�Ô��WyC���`F*nn�_TT�O��z��EWp�g���
5��̢���G���#��8���Ƿ���7ӡ,��7�-�`�x�~��JB��׷ֽXu���p�C����*'�y˹m��jNӄ�@�Mo%j&7ה�_���[��"A����{�a݆��Ug)�����l��� �ɋ�|imfj�^�ݱ�ɉǺY��}#s��c�˨B����O�XK�Ǻ���U���6�-e��?^�&���h%��o��{QRRr#sS���u3.�k�5q\�Y<��ʲ�X��򔢬ۺ��Q���la~ў0��y�����\�Ù�}��e�w�<�j���gT���	�臢R{�FW�zH�����k~OϾ��w؝�[��X\r����A:䑳�w�)E	K[�>������3�ܧ<��}�@�E"�E��[�X�r���M�w#�Z��N����ػ��3,:� n�8F�f�LK0���$i�F�E9!�c(~�'�W��Kz�hg3�;A�s+k�!!h�ٯۈs�����ϫs���^�(��_7ISeŻi��گ����E՛�	3�.cJ�Xl�?]���DO�@
�9��Η'�eD�1�̾�(�b�������O1�)>-���\|~��(#���8����twKKKg�G�&�~4�\�H��m�Ǧ�{�ĸOHJ.f}Fˤ6��:H�?u��f��f�J��+!�O�����O~�Zز�6��HW,�ʚ2z�6�a��[�����&d���ę\����u R^�7���F���|���+�F����{�5^wY{3(NƁ���w#ΩUUUB�h�)�mX�R�M��_�˾D*4���>����rXU&.d�!(����ۜ%:k��)�*�*G-*C�5mڇ�/N����us̲p�������\]��G��'H]�h\��?e	{��җ\TUUW��AW#��]wumy�/%�t��)؂N-�NY �7w1R<�-�as���D��//�uY�L�Ѽ���T�f��Xu���ER�-w��/OY5M�y��`J��������n�Ͷ�3�e�D�d߂��r�5�S��U[UWW����}�e�y{����u�Dt�����3��Oi;1��%L�������^g�����(`E����`�؛7��m[����i�Y� �#q��Ν;o����A�,��&ƽjR��7�2qm�Z���R'qO�o�������gm� �<�������ϕ+�x0����Z$xq�D#yv95U$ ��[h�O`�WF��Ow�1��p��v��+�:�(�>k�ak�o�3v�8�lp�Ό�rqq�+`��􋰰p�9�.�9�ͷ���=O���n�ދ,z��{���CZ��Ζ����i�q��(+�۳���ʒ������G�1\*�cA'qϽ��=v�#D�T��l`�-{�i�����(����9�G�OJJ2�%�`�Nā�K�L��^���S�|���5�
ПgQU�YN3���}E�Q~ ��(m� 0�9�gb,��n�̒u��]\ḇ��;<&��&ɔm��b$�+J�� �^b�oꞚ��M� �	Fh��W�2'ǣ�#�/�q�)�.fx;��wqD�j�@�m%=� �̯�l�Ǭ]˲^���ƽ�T�VgM��~�yA��=afVzw�����(��e����A��S%y6����O�摈U߹�����D�k������OM��n`���j�U�B'�Kw�l�Nn�I_�x��Һ>H4�*��bۊ�"�2���6�@�:��$�+y7pI��`�k�vQ��.2Y�,�@	Ϸf�c ~9��ɝ�*����#(K"���>�\�돸hPL���C�y6	{P�v��+��ńF��Q�p4R����b�A俬6�/�N�k���A�#�L��VWW��X~0����)tҵ8������L`�L���@��������+�z��'�V/���U�� ﹐BٍT��U	���~A�H"�ވf՘�|i�/S	��0��[i���qUn�ḪaN"D�b�(�Z��"��Y䭱�,��=�� )W��4�.k㘪ś��I� ��x��/��ܹ�d�f\Ov�S��aPf�Å4d0g��Q������k��=�Î�Siii�ǿ�,���?��p�"��	�����}f�fà�,�:�=�o!�}*c��L�g���`���S�#)
�q���x�eӭp�"��}�36i	kU��q�0hmm��I��Z��&�y�0 �����)�����LY�(I6�	h���q�g���VlD�3ov.l� t���R�:�[�)��'Ѧ��"k������d��oġ�$�2b�¶i"�򼔔�s�t���]�Q�%�g]���\aQ|���e��I��&G��)M6���&?!�؋�<2�U����Xg����̩�Y�p�$�_tH�b�d�u��i��O�8*Y&x�T&L���}~077�m~eM��^'6%EGG���Z��kp��v;6�p8�cjΡ��&�R����=�m��:������+B�����!i/�y�J�s��Lp���Y�����d�yv�h'a."�Kn��)�ri� ���C}#�ə��P��xg";^
 W���/���򜄬R۸]v�DZ |g�j�Μ�8��̿tb�d�t�^�dG�Gi��
rHx�S��N���F�(��t��D=h�5n�]�R��S�����eP�g$N����B�2��^ߍq"�7��,yiF4,(����'�TE�n�F8`�ƅi%%�1{�T\�B��e&�z�S�&���ƛ����� m�Xޞ7>��~��.�Z)�62ȔA�2��od���Y29M�!�Ǚ�ϵ�N0|����ݛ%�w#*�ï6|����H��<v?j_!��,΋FN�_�Ci^x9&*���,��=6�*@��d��U�{Oq��ރG=�n����B���ߣ��ֲti�����i\��W���9�'!���n5K�Q@C	9I,�ȅF�}P)?���㛒zt�=t[��c�TY0��fxBL������ǲ,���z⦪��R���T�����ZSSS�g�Tg�X��g%A�蛙�Q'����mc�P�ؽ�Gi҇�1|>��S�$�wR�J(n<{琢��i���x�2V�^�N�,--�`"� ��+��v��+�A�Ӻ��u1�i�.�zK���5З=���� 4��Mi�� %���{OyA�sD<Sx���e�������kݠ�r@I^a�+4h�V����,7ۄ���j*��[����n�6H�g>�u��k�c���7�>��V��:��|/"�J�.2q�4���x��:;n��s��n�����>�|J��y�֌D�La.�"�'��R�	PǸe8�˝��!�
�7���<�H#	H�l�&
Q�vO|��C��6�.J��q�M�F���""͐�[��"���*�n����y�b�Ni�a?��d|3fX[#���&��F�}T\�#Җ�l$��<�j7���ꃲ'�J"����X�Ƣ9���������I�0��͵�Q���~S7V���2B[(W�Rm���m�"Ng�gC��<��]�`Z��v1O8�d�"k�Z��z�)=�PŮ��w� yh0ªk�gS��֎"`n�����y[�W�3W�͇�)M&��
0���~��,*;��Y������VDZ�\4�-�X|i��Y��r#�~++��$��@a.�Ir��|��r#[�!��{/T��N^��ld�h�}tɑ��7���/q(�����d�x\is0��6��)�K2J@7���ㄫs�LN��nwi��A{/������&&姱�I�^g^����%IԴHI��ӳ�ެ�PfB`=�.�27�,I&�������e���J@q�!�Ҟ��^�*6W���V!�@��-�jծ��(T[M���D�!�X�����m����Y��'0�D����g��FCM4��Q����ޗ�>'���ĺ>wo@�b�ߏ8���+b�M�q]��.��X-�٘4r7�f�	S?�b�-��yb)�s���j3�ld�S/<t� uU��)�%L�x�TD3��<�ǒ�Ⳮ��HW��O�L��.��=�ʍ�Q����§i ��LL|W���_#��<0��/��Ҥ�0 ����n��FEDA|�x���JT����u3��4�2&�����r��h�eh�M�z�%�dܹsg2 [�{��ø��J������+E�X�l�
	�(M���G���6hLU@�.\w���T��S�D�n�V��"KS*��q��W^0�8�F���������J:''��)ER�Z�V����fyJj�N�<<:a$�N�-���1K�3�o�`i�z�s�����m�����*}�6�]id\5>M |:�g�'WR�j���X��aZ�uO�Կ%�(����У��4�NBz�3��\; w�^����9���ݩ3O�\�8b���������%����;�t�@�e��2?>>�?Q'-
����U�8��$��˗�	�'1vbܫ$��$<�S����6�Gp_6��O)�+�gK��gH����0���;���c���&���R��OP:n�}�۵��'����kl�,��
O*v{*�F�\�6n`W����_� �w�2BQC^�������	l�T�x�΅��Ԓ��p0��fC�Ջ��3"�$`�̑Dq|���FǕ�����PR�T#����BZ�to�Q~Ď�dބ�4a�?:�2s ����6�B*Lbx~,N�ӕH��By��D�!�>�vۍ��ٗ�-7I#Ch��3JS��j�6�N�ҷng_����ݒ4�'&I;���ke��㠡&�� Ȃ�巐���@��/��07���F&`T��xc��}��d.,�qw� �Dժ��<����e�!�ۅq�Jh�ܐJ�򇩓�x}�+5e��7�6m�m(���&S�O�c9���8'���A���z/ GO���`!���\x��? ����sƨ�����D�?��W���8����d�Y�
����8��Q m�j��`ⵇh�nnn�K�������^�slhӗj��,�XIM�Xn�V�T��p��:����q���ڬ"����\vƟ�;J�҂���q�6:�y�������>���"���d�/�$J���W�V츭Z�B����Z��\�BT�e`�Mc����(-c>��ێ���I��7��o�\�^�+�ku�!�k{`rr�]|BBB
g�'�3��d�)3k�C���o`�8��J�y�����P�ո/c��_��@@E�L�F�U�/(+��5j�8�|AgK-� Y�4	��á����tn�����:y&�W��IQ��C���n�$��LC�6�+�}&���c���6H�cO@�yaÌ��\8���S�ƦqW���^K��'CCC���rK�_�Y����+=s�҄��<�Vttu'�;v`r3q��ϟ?71�����+��<��Kr
�j�%�s��C��Aǐ����y�$s��!������K	D�j�휩�-��(TX�:�U[�e�@���U�Fh��z�VE��{�@ ؏f�Ct�%[����?֑��A�>��+�(:2�����\��=IM�-�y)�Ҵ��s�$&6Vv7X� J~NR��o�"�2B�/�5�2%%��8�@��q��K���B~�\����%�6�?����b�%��i�0\����h�,������(-q`��o/�Ft?�Q�� yj�B��C[[{�0mN�u�V�f���&�V�[qs�?�z'�I>�m��ӟ0�\�Ч��KN��d�n�ֻ���㜜���$���w;�{�YFT����7���C7h����Nt	y0`�����U'�&o�cw�^Pwʓ)���k�͑�p�8�醟y��P����Cm���@C+]�z��Q���h��k0muK3� ��%���e|+�2����=�Η%%�M`��>a�Ά�m�-���3��@V�`��b���y� �%��2cz>jB��G�`��Aט_GG���R�ص�"���](�W���U�_60X)�4�A��/��f����%��Φ�[���\#%��}���4C��C�|�t;�zz�Z6��쮕f�$���.~<?������I\#�uy8d����h����e`���g^� �=�ow���z�о�y��U}}}:k�d�,� �[���鑰��E>�tL´�r�"�>��.�x���3Z$Q�ç��z�$��iw#.���D;QZ�Q���{腧�(��N���M�6�?ͻk(��ێ�O�C��~�� R��~
&`�*���DE˽mm'������(l|�w�V�$�&�bb����_�;<Y	0[m-)Bk�R0�����gձ���	�1ץ��+�� ����ˎ��z�GH�Gz ����.��\ns_��u��cD���k�-ΟQ=����e1��w�_��4���+���jN�&����n��ݿҷ���Ͽ�#�I�q��gǘ[�6J]��:���o����w��=־�䛜t��@�XI���ť�g�tn�5(\fb�%/��B�0O��0Vx�?CB\�#gv�e�0�(�\|h��VIՌ����(���<�}�����b����p�k��/�����qq~�87VXX��:���}���b���;��J� ��=>�������A��$U�ʇG���g9�ui@��wk�t�l�8D�w�����LΕ��ù�
�+�q�@��5��L Ns�@�$<�ʜ�9��{3U!"����%�e�_'п��1;J���i��Ũ��ַ��h�G���R^�J^�`n�(��.�`$���:=D(��S:�=Ϧ��l�*	B��M~�832*j�"ʚN���ƙ���YaU���2W_r�={��H���v�����I	�`Ȇ'�y�7L�͇����q��>���[�'�tpN�4&2��UN|�����D�Fg��f����5RM!R�A��٦g�f#K�Lvq�������K�ž�v�ymT�6c=�Sj��
�P�jhl,��`�FA��8��\��I���ir&�G�f\ll�����Rt�����4]��T1 �64�bk���qa2�9k�٣��4mR&:巉N�|En�����v����DvQQ�4�z��?����N�R�nL\7�.�u7$<\��ral�)}a����C�t�l��G(M�Q���b㔦�ؤ�V�I�b?�*v0i,P�8T�ґ+i�n?_[[G�#�~C	�P���V&P�vD�E�r"s��Wn��>*�r���K�?�Tys�뎹,�l��W}�Q����Ck��b����r��\_��vS�/�!͕�:=2��~�.���b@ ���N��7S}��=�MH(?¯�����P��EP\���n�5>m���Q���R�"(���x�-�f	�a��7<��c��t+|�$EVΪ�Rg�_�N-w�%hABټi��ߟ�(� m'X�Ej422*����C���eY"x�L�U�d"�8Y\�� jN4J��s(��:i�K�VM�I�Z�nr9/w��Zrs񔕼R �]l��R� �-W1P�ow|`ίk*�	�߅Y/��Tt%��?X�}x��xr+�E���H36:&�H$~�AP��e���yү$����Aۼr��=�h������@j���A��YZZb����� �j^�'�/A_R,�r�1,�.��/�!���� ObX\^/�(����@SX�.��	��ﱵA��\�y����6OT��p$�]��f,F@���lr���7#-۾��)��Հ/�0�ڃ(M� Y&G!�g������u�̍��Eg�9�Х������/^5l�;2q�|�t��,:�ejl���Q[2���9	��" x��;�'$%���L�m`Zy��]�u�K�C<...���U�|�#諹����C��?�X����j����62�}X(W�D��}Q��} ����CU�2�
�Eb�Џ�!y8Ya�@���t0VbC��X[��{J��
�Z�X?��y�6�J_�B���]	u's�t,kG��^J	r����2��2J
-c$�zJW((ӄbYId/�qU�j�w��ƺ
gE����I����ׇG���h�U�Do�FRDDĤ�����s��"E��_'+W� ,�� ���zʁ�`_��҅٪X#m��3[�0XWW��Jj�~WkHjjj�J%��e�9���޼�\��7:�6����V��K3�Wָ�J�\~f$␶���w�f(E$õ< ���D�o4�D�7���Ci�����ح�(ÂG}^|ޫ� ��&ps���U���g=]XX�3�7:�<���y3�G�*��U��+D�]���B���
@�%Q�W���ǰ�E�H�.[�/4�ɓ��Q��_���v��^����q?*�se�{�9Hr�nNN�������h��(���2�f5bi)����ӡ�:�-���=�:�'t��b�ER����&+)��4�w�<-�����J������4��6(	~�K�z'�0�xV�|��0��ߩy/�W��)����lx�-7�)��W�CNA����[�J^�M��z�7:A���{�� e$���"�	e"�U*�e�`/��Ao@y���R"��p�}�s���U���Z1�z�~����lC�ߘH���<q͞42�a%
���\���K�*ʃ��/��!Q�Y�6��H�����r�btt4��P#��b��Vu�	��>S����B���6b�|��E�n��V����ٶ5"�M��(ߓ���[+������J���� ѐ�ds�=�En���O�R����=N�M�j	���a��L�"��` ���3�l^���q[��В��~�Z* �߉�8�H��_+m"�R�6�@������ݒ("���H�&�-����@8��{=����{��0O�,�ۂ�KFAI�O.��#�}�y���t0�|�	��cz�}��z��Aj������bo�f	�c�}j�����ݹs�SO�gch �c{�E�to�DG$�*��K54j˯��@3�Y�L_�$ю�^�)��NC������%%�<����A<rj�-��p�P|	b�\�ٶ/K#8@��Y,��de��4*Uj�T�#����^�����sYд����͹�NL���3uĩ��<(ȏ��(�U�𮯡ۇ��%���f�T"��T��?[ZZ�ӟ?�B!���0��Y���@e~�����8Y�Zֳ�,355�s�
2�T�
�-�pY:Z�ϐ~��@�f@wg�v~^� h�<�Gg��K�e��T�8��y���S�L�E|!��v�~�2i-7�A�p��\�KLg�޽w�x-�ȟAЬ���i�B��"�J6��*�S����ZE���ǥVQQQ|�h%�R/��l��+55;X�K< ㋷�~���:&0�<��/�n��d�_�)(�-�J%)�1\H�V�l���MO�R`�����h!Y�������|#� �������^��JK�E�%���n�Y��f�A.Nd��!j��m�u?��g��� mHP�H���f�eA���i�[g���Ql��S��G�do9��\@J����뻻�>:1R`��7����R`��^Na$�F�/��X�����N#ᴸ'�LBw+�C*I�6f*��R>:����G��S�H ����������<k�^�nb�:����S�ՊW���Y��ô�u�ʴ��QJS ��KCf���$T	`h4�[?L�:w��T&������#�����
���fdNy���)W^�\�:x�H�'��Ǣ��B/��{�&Q�`���&�gym�5�~�'�z}����5�����p��O�����lT�^��ߓ���̿s��˷Z:�L��4"V�W�Ł~ о����UG�1؄T��S{����N��J�Ԫ�]��'�@酻*�؊q����?�'hO�,F)W��Zn���9=��4K����)��#YvL�0����V��%�C��y�g���ǝ��� �XE��suz!�]Q8�~=V"lh�mo�a>�$�� ��m[�hQޝ-����;��)�cǎ�I�v����p+!(<���P�>��i��n���s�N�V��pJ���.�$�@v)�"U�����!�1��?rf��5L4y��@Q�p�"n~l*\p�[iEx,z ?��<X"�\�;v�rp�f/�y�T��O{�����u��)+=|`�;u��H�9�E����ǈ��̋�6���1Gz������z���as��B1d.SWGgBj+��$+�?����T�������|;�R��[���˃��X����#}���u���W}��6O���5���3�C#r�����(E�Y�5��vpY�&i���OS�+R��w,������6��g�\��4�R��)��Ν;_����X�C�u���ʒǎ�N���S��a����@u0����P#�6�oB,�Qi�o�4 xu-�f�T�Q�hOQ��L��~#�ߞ�i����3,\����]-��&S}\Q�Ͻ܅Z���haG4�~HS����Y����f�eܜu�Im%i1�©���9�RiF #��ã�Ux��&���2�@�^�
�y{@T	�7C����>�#ӆ	���<l�z ����ܢ�9��N�[�'���=��R�8̿�Bf������(��
|�?9[�7J���j�T�3?;F&tnv�	h,�/�[��%��� q��;�;�<\#���QH�'N���36.3���Q����v�NUL+�t�:h�f�\���.S~�"��A�]�[��g6�FG`�#�'m@���}󺛑F^˺�����ss�Zr���U�c��@;]?YV���p�(/�X��� ��'�ɐɃ�*��9��@y�9���iu�Z'm���5< �٠0��a��@&jb���D��X��$��yo������1�s\E�2!
��~v>H1_��Mَ������rN'c�Ϲ���v��b� ����D6<hx�9�ďM�k�T������TL^�����|����ن�C��/{o���B3��
)|:�'������R(M�T�7,!�@�Dy�ܤ6�%�m:��\���,]��Q�;��z�|$�4Z�Sy��?��v刃�ٖa��i)NI�f�Q@��7���
Ӓ��x��)����~Z�j�:0�*��6Ee*�AAQqG�
deY�DA��j�4aɰ��(� K�,���w�r�������3�w��C_ov��1j����F�7���?4�J!E�
�^ǣCW����!�Ą�ҹR�/�k,8��o=G�[J��	��3����)�3}���}fUku��M_�p|\��=�%u,�c]Gkkk9�����AR�/ى��Q�MaRRXVRVfq_��n��Dg���anV:p#��w���e�M��Ōҋ\U�#z�\zh��Ǒ��=����g=���5P�l������	�g({�:�s�T_PA�Z��Bk����dp�����|wq!��Ǧ�#��5�?N�IS�8��0�Xy��{���\��s�[�g5�^⠅��6nV�jv�mX�(�x���\���#�������ǙuO@�WY���t�����e�n�f�� Eދ;>��K�y�C��� ��*'��s���P��E}�VnZ�5ZI��fY�s޻wo�@������}�?`:9ސ��t�޽�cy��I���?�s)��ܺt��/e����x��/\͝hD��9uy�����l��Ӟ�n{[���&SZ�s�����ㅀ��S�}6Z�!L��t`��t�vIFg4� , ��;��!@�:���r=2��xK��)3e#��i��ɂ�.�u|m1;;��4d䩅��+F����^3<6�������傕�5io��G���b�r(`�j	��Q��L�5Y���w���x��}�&¸t�̕���줾��] aT`p.=gc���vP�i�z�ܹ�{��>Ҳ0���Mj�ճ8��;ǜ={<�ѿ�����^h5'�ɚT�GsȀ�I��]�6U�Wj�����R�{wd/��<�@�G��g+�b6��*���o޼�B���V����" �X�y?źf�Kt+�f���>���т���w�)���K��#�u��8ٵ�<3Ea�.c4��[1d�|����U�cGM<�L��������n[mq���K�c�x�N��/h�=�I�P_�F*A����^�;d��f�MH��Iofһ��Z5?��3��_vLA�<�>{}u���%�θ�k�Wo����a�f%$h3�,�-Gx�P^���+D��#�^�w�Y��^*&"����TR�Ϳ$�n�u�3���P����F��K=�0��l���2:ԛ�M1�Ը��P���y ���0���֞�~<ߟǷ \�x�9C#������v�in%�?��ry<[�Zv�H�:2��?"���>Wa���qH������_��.![��٘0mu9}��]9��l^� � T�;a`�t+�t�l�B�s$��ߨq%�粓�<VR�vU���q6ױj�������[{��1שJ	�"H���1f�2�-�dXE�{C���	��򢷇��S�qZ0�ʺn��		
���:*� J�i]:`&�l���e�{W�1����?�]-\����Nj�Ff�C �*�`y0N�D�����nb]}L���hŀs�@*��:���߄�5}n%�v^��f�#j���B��}ł��ʲ]��1u����u/�&" �Kr"��Oѱ����<�=�fy��F��\�)����e��z���]Kv,�#��d_��`��
��,`�&J��8�߭�g�?��ӈ����B��^S}޿�j�,��$M�ka�S{���m�u�=�@�M�Z��4����)N[�\���F�%��}� �:��l���@�t�: ʤ��a�H��0��_��,܋aC6,X�[-�+��p�O�l�6�.<@�#me�IHxϭ�O���h��9@���ѐ��2Cn�Y����b�!gT;�P}��dY꽒�����.�~%�%i� u��TQ�~l[6�Y� ���GaŒ�{�����
�Gv�Q��mY�<���T�{)e�A����n���MK���nX\	��w���f�MZ��޽�4j���utܵ��/;��MG��Ka���>W�o��B?�ҭV_�.9����?M-޼��}�Ϝ��W[_�:k��)k���s+����By�[��۶�¬�?���l��fz� o���7|�����|Y��*nȻwʮ�׫�v��<~�5W�ox�CB�Z\i[[��D����|�f(��j�P�6��*Ca�&�*ԫ����ȍLG�l��4���[�y��־�	���/Ճ�c��|>�~d�s���J��X^dN�b��s���0!��P�HYc޼y��!j�� ����Q_f��QZ��]qs���ن�����f���Xu�ج�*⪪����^���d^s�ݳ�ɥ����2��6yp�nvke����'�����U�r�8�gb+�a���D]m����13739��:�8K��ϒ^7��.��9 ���5���#;�!���t���?����,omjXɴ����I���@-2�X�qʝ�� ś��k}����
�Z�^�\r��ms�^^jjW
�U'����Q�Za���ɸYI���U��s�����hů�~H�;H�������ޡ�pt4&�}C����+AS72�}.��B�ǭ�R
����c �^;PYӌ7U������DJ��F��G�k2�����ϐr�[f��t�1$�y&��>��S@�be�����ݟ�*S��:�fGj{5��Ǐc�mթ���&O�AH~(//_���#{�)璲�'��IN�[˘a����S��0���!��G�����|������] zl(+�ml���@sP�?�ĭV�?��ƄS���=��Fx���g���D_T����)L��r7��X��<i�-X��X���X� ��j���:��Xpa]�C��t#�����i�'���~yx�#\:�|}G��6��5�k�ɓ'W(#N'�n#B\�M����2m�z�ii�1E�el��~@"�0��������ξc��vWG(��Y���ř��7�%sY�Q��UX�?g�(��6�Uc���{ۈ��&�v,�u�%�����b"��&_/{482������3b��f&
F��\����w�%����P�����6>��%+�z~�,�$١Ƙ3g�z�	SXk�v��z�wO���8�"�Zq�~3�ʹ 2J��'��r�X�%w;-��P�6e+5����>���Tzk~�޽�0Ʋ�@iA���K�g҇����bw��\p��?�j��Q�d���+L�s|lǳ�m��}��R-s�[񈾩Dx���c}(���Gg='M���'�̭?e��(}��<�=ɷ�τ�z�|���=�Q�^gѓ��ȢR<�|r����~�X�Xga���6�N���U�X����V̍�b'cQ��]�w��1l���A>
W��+���1Vw)#�"&(��j���Ȍ<V1ŝ}��s7��S�l��u�SQQi��!�!W�^rH'��r�lʄ����l#TfLv�G[�Z����B�	ǽ��s~�����4�Y��d������&�j�n6	!�?�q�ܹ!1��8X�^�>q��! �2�kb��D<��0n`��V�6'�����O"4�w�q5�p��o�7V-���d��q^>��_��W����ɹ�/8���e)[g�k��q��]�x�bU%e����nL<چh����Y�s��m��|��3���s��5���`e_�� R]�(ɰ���5�����x�s��u�L|9j�m��k�ǭ��5"��^�Z��ו�V��E�h�/��>E5w��}/�5��. �B�j6�Eg��\���/WwՈ�))��Ʌ���?�Q>�E)+[��
cR��?>�zZ��n˱ts��0��F�r�X,�RS�YN�Jl-��G�=k���1���K�c?'W�:��yO��%�c���V|ށZ �1f�/N��x��8���L�q��3_(>y�孅&��3�u��SBe7�h�{�%y�������"tkx2N{d~(��sR��=G��ID�v�4�r�����lǗ昃\���Bz~L�:˖_���T���*'�[���$�C�����eDEJc郗�b�}��$���#�W<���k�XB� ����`�K����^�.����Q:���M�[�&�T�,�����~���U[o������Yqqq:'y����ku�	�2���=#�)z��l"!�"*�O`\oqnΪ�:�۸��Y�����@O�����+11��1�	4���B+ԧ�S��֬×Ń�f,��`#wvivY@(�F�c��z�/�xs:h&Ke�ps���$���e����>F���B)0Dq��atC����F�"K]YK\)I�j�Id�MW�l���7�*������_X�nxx�!"/��=��K���f��[��6l
�6�q���Jɷ8ڤ����o�Va�G�r+�r}��=�M���,�i����
��Ul����A ��l��Pl�g+4���9_ӁX�B�$v}�ZG9��Y5�hk���2��N�L�n~�=`�F����\J����e4�S3��9����D����8��4
R��֥\�������q�T@ů(&[�̖Bo��^�P�ۀA�O69�V�v6�]c�*1�"p��ڐQk�����%��hA<�}���E����L�h��@��0,꾥����+&��� ���u&L��$K�b�B'�%'"X
�oː��`<�!�T���W��u�A+�	B��<b]�d��VF�Az�e���-Jr���jʼ爪s�	��o�?oE���9�)?A��_�4v� �w�jߤH���c�X�q�\"�?�
:=$X�u�]���1���1�%�r��.{�H�-��w:�P�b�-�ލ7���/.���ת�M9�U��=gR�
1�cm�sZ��"?%T����D����rO,�(��,�z�h7����"	�MA%�����M�=����oH���t'MpZ�z��w=NH&��N�ژq���O�ѳ��ϯ��ɩ�O?��ƛ2x���^&#7QI�B_�4Xss��A/�@c�'M���c��5(��E4�*_����/����jb�:�7o���*6��5uZ�9߂�cʚ�X�y2�ܥd�GYǄ��i"�5c,�9zכ�_!_���[�Զ���?A��d����F��x�gr=��?�Q4)��.�V	����ty�)Z=e6��*=����V`�1��� ��)P�@�z�-��.ct=.��2�ɓ"Ui�7�ڤch�[
NOҘ���%���d�t����u��h�� -���b�#�wd��U��M�x��XA�ܓ�]��75�ɜ5셾�*��>��Fx��|B�ƂӪU�@n�k����h�Ն嘠:$AY,h����W�M(��C3���-	�ύ��'%'[̒������$>��*���x��@��퇥�qm�:�p�2�hy%R�[@�:��F�[c�J*P�ʔ�e��3������(!.dܘMO��f��h\�`9��4���	ǧ�������|�;D4D�.�st�����M���I�r�ZO��H��m�33�m��H1�ܸ��^�x0�[����J ��X5T����_�K�gүnuQku_�5����>W/�4b[���F�3�̝|��vE@]�qՍ7�7�=0)���e����c�*�t��<���^:jz����y�k��bo��W>����/w(79�S�C`ͤ�������56����������=!K�x���Z�w�o�L�~����P��hR<�i��Q��F|+,�믿b6�N rU��f�4E�c@D���P�R�]��L�	u�q��j�ف���ٳ�]8�d%�b��4;�wS���Q)ӡͯohwW��c�^��f�=��感sQ!�I���������������R6�������_Ϡ}�_�M_�1�Xԏ�o�ba{ �	z��(� �$)A��7[vlCK�7�����G�TVV~ĺn|�h?c��Z�sv�ЗN$�)*Z@+�.���*ӏ)8���;�<�y� 	o���@�6�O��>�%%3����&���ك�c����$�������U��
�FXJ#��r$����|�
_u�Q�Q1;9'+�ݝF��o�P���(�����2�|�U�'05��遁�J��P��照\\>��0�˳���U3���d(Gs�y�P�g� %Hq���$��Zn�\��!�!���v��Vj�`x�͟�4�n���d73V������i��j7`�h���.iZR� ��
���H�mA)B��u�g�r�= ���C5�i���,E˗->��k����Ѱ��'�bhG1�*٪��dܙ=�9�7m��E�?Kz�����N����cyFaaa���$���z%���  R�J�\���`1.A,E����飉�5d^��@�wQA�[����8=��ö�9�u9}Kq����p���f4� ϗ�� �|����y�UW�#Vg�&����;ȗH��5M���Eˇ�7�&?ߥ���%�8��PJO]�~���W�\H�-�2u���78��N4���fՊ����ki|��8GU׻�Q�0&R̎��X�0G1��C���.� ��JVp������9���pw|��9$y�7�-����|�X��`E=�8�"��>9��j0�,�Ӛ%��@>���A�Y��-%++�&��I��fn�,�A�A��rٓ�%�J2	��a5uS���Ji��h�Ϳ�d�� "��`]�xJ��2-7�ŉjkk�}�ҋޅu��N�ڙ��P����qf �#�����=������
]�N>ٶ䪡 ��W�&l�ީ��f�ٔ\�t���
;Ŗ��$��ݑ��}�gZ �i�D跋�s�U��s�Фxu��O��������\Z����{nC?]�ZO���Qs�i9�Gc7�'���$�L�#�����e�޲�S�g�}ǣr�@�rr�
zY�%�Z3��8dk�C��[��E>,WU��wb�~�N&�#^��o�u횗>kx+Z����޾�> b�kB)uL}�<��Ј���I�N�/�		�6��^x�;�#u��CG�{���3�-!�:�P�Q��|���P�������[(�*"�c$^G�1��q� ����Pw������?RRtv������Pr6F�\ �D�� �w�c��%=l�u��U�q|�YӰ*�^=J�>�%�h��}�@��)Q<x��C�����_s�2 ���s�|=MxLn4�s=}p���ӈ:�=rlI3�ʌn���Ŏ��M����I:Zo�|X����0+�ˉuOr�S�M�����z���t�!��.��.�����b?"�-�I��i��q��	�qTS�]���F,cw:�T�2��Q/tV�vq@#���V�
�5B���j-�7�ɚ���}C~3�����?O� |)���7Ѐ��{����y� �����/3`�{)~�A�儘2�y,O���r�${E��[W0h�U߁����x}v����g�(�n��&��\�`���jw��i@x݄�"�Z��cT��J��j.'�k�
�������Ƚ� '�}���<R��{�U?�u�@T��K�����(L�\�]�+�٬ex%��؈�Ox�4���s���,/���KӫG$��7�m<��Xڰ���8�P�����D�KG �۪S��D�ϡDI��%�y)ѹ����⌀���zW!��٭���z�XT	��!s�y�M��0�����\`���^U�A��5�-#~���0� ����y���K�q�oA��?��j� `���Q�J�@�A��1<7d
*Zt�2F�����c�d���ʠ�n
lNms��6'�UԚ:uj��;��d�{���G����_�q�e\�a0���-?d!��cµ�z���C�|=ߨ�k�o
bL�^��T��kwo8���rQ���_��0)��-���b[�BM.E=T�g��W2��!N�]�y�&�PF�'���	�yO�YQ����\�L��|����nj��f١�K�x��u�Q����ܔ P�����΄�� b��l��x8ڦ(L�tj��^j�����pQ�����=��#@���Y˅�n�d�vv�?0�G�J�y/=)1�b�2c~�m��k>�;bbߝi&E��?���Bk�(X������#���]�Q��u���߬G����sKp�{�ă�8D\��S�)����>V��f}�k+��-s��#PC?���c�#1�X�T^� Рq�r�<Iϗw�5���`��=�s���_�D�pM@�}�;�;����B�U��{�%��% \ރMixنl��"����֯c��B�7_���
-(�������C�$������X%b�!Sa���E��>�a?�I�"��th�jh�Z)>g����紧,Ƕ��(0��|I�ҙ�z��uV�7~s����nfZ]����3Sܸ�����=Z����1������;�K�҇����k#}răg�������]�0v�%�zI����X��&��X�&>��h��p=�t�0I|r��6yT�j� 9�R`�Đ�g�A�=��[O���gCX�9�ܖ��<0����r�z�:h�����X�x��%!���I�KC�Н��O����,�q{|�~�&;�i��g�+��\o���2|��j[�Pd*��$�$��80���?�
�ί�H�'���W2�Q��Z���>(��s&�p8�6C�&d�A[�45��CeZF�4�^���\���e��a!H!�4l�z"=-�A��$#��?�j�,S�`�|ve³��B�i-�����A,��3�M��o�mV� ���J��V�Q"�q��zL��������/I�������
]E:��[F/���!2a�ؑ�G_	����CPR��1��'�2 �7��H)D	�&����G_$��`�;�wX��? �6fP��L8���*����������G�����Hv�Ü$� �ig�62��{@��,��@�}����<�������[u-�R��Lg�����6�|��w٭-]�$���Jzc�,Z�7�'Bܛ0�Roo�� �\�`���8F/�6��MUn#GR=1�K |�8jc�����P8:�� 5��;�+�g��yCW�~.��18��XҚ�p����苮@�8�F(q�Y��BSz
��qC_����766����]V�����a&�Ka����"W@�qiii���}�OU�%W���聀���"# *hqޣ���kt'����a=�<�Q��u���~{|>w�Y�L�!��E=&œ�Nx��x����:^b�(�͕
�\���AZF��b�y1�i���cJR�qKvR��j���Zu�eh7R%h?����9/F�7V�+�8L��H+X,���J�u;��x�DQ�h�y̬��˝�ܴ@��;6L,� )_�״U	��4E�y}����gF�@����6	"��h˶R6W
��Φ=����eR���(kV}Ύ���zտ��hjz.c�^�M:��5�G��Ϡ��@͂"��_����6(NЧ�|[�~>=����,���J�~?�z�N~�	���)�͊���>º��ݤß�r�4J+��U�LE���Ķn��i�x@a��E�U��ڿ�rl����a̐e�F��iP*s���Z��ߨ-_�Y�č?]n�ә�I9��s- 7��ʊ+�_���K��9S�[(�?�I����5p��S�Xd�Y󯉵�_Y�ڀo�5�&qBޥ[Z�]�vt�a�ŭ��~Ox����b��åf0/�ا���p6��[�a|�� �Ԏ�XS�	�f-+!���dO���R$�m�[��:��XުG���*�J,�W=�!���A{g���]�-�K:6�F���Q�?���������c8�����Ol|�3�����!��3Q[��bd��
�Kp���Ƭ��Y��PK   ���X��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   ���X����  �  /   images/25cd0dd7-bebf-4a92-94a8-2c258b16bf7a.png�W�[����%�0�HǨ�H�tcа!)�]JM��5i�)%����o��y�=�s����8=5b:,,,bue����@��� ��?y������m�l������S���+���������[w���������#(��������
�02�}X��t�: �W��^�Mc����*��?�\/����;�~�*[��aQ��������H�J?���S��.N��oC�ģ�~�}����Y���b�����ǭ�o��k�I�)�a����WE��q(���_2��_Zg$'�T��y1��W�V��D�xVn����K>�;�;�!��#/��GyȎ������	�KŇ��Q77�-�F���Đ�L�&RN7��Eg�-d�$��8��''���T�@ �7���B4�wwA��nt����AAr����1=W��^l�������P��� �sa��Hz��N�[�^e�wc�a4��F����k�w�a&��ڷW�\1=�H"�)��=X�W~�s�@L�r�S��������N��a�W6w�Vrw=6�s&*_Z�G����"�����1����}yyy����)�:݇��L���E푐S���Z�7-j��qڛ��5G�|�y�H��^�ٝyiS"sܖ!�H���Yc���Q��ؿ�H�H�N��J����ৎUOPJ�%��<r��֯�宭���32?ڼ!�^u�x}���T��v�˥�������j��ꋧ?|> ߐ#����onl a,��aw�������z�����z,kjj{��g)Z�'�������2G�l����]fJ"��:ɮ�C1��TT����{������'�Dd���3�t�N���ϰ�6�ե�0p�Ky����Z�KK�u�%;��2¢s|*����d���v�������+�����8^O�^W^ν��
��]l$�U�bJ�Á���@U>>�m�.<��򪪄����Xo ���Y�o�j=�s�kЃ�%a��P���c'ēfP��
��=3=��;Z��:�{���_5p�3.**
Ԧ�j��=�5���̹�9{2�2jxl�_�HO���}2���x��Z���Ne�mieUU�n�\�]>�u(.&�I�G�Ml�Z��4�4BZ-�	4z��]F̆�r����=�sm49�ri�Y��-K�̤�$��'_Qw{7�|����su����I���ߠ�'�����aq���p�1��'RKdو����ɢ��$:1����d��N���uȿ�2:BY�.���5A��v��@�g�8�H�#�ʶ��[H@�M""��,)��XW�v/�꥛d\JPO��s�_��W�s!e�f�"e��n@�[h���;|�ZXǇ���߯i2��M�����ӿ��P��1H;Ar�I~��aZ���|��ȰϼP��+<}�	���aziV}1���.����g�ͧl;H��C��VGloKy�1��h��7Mfk�M�JxO����z͎��=^���y��R�g��Cf5� >8$�ٟ��2��<3.�O��%���zdE��G�M7₇��ԔW&ڔC���2�:e�<��ؕo����X8"m{��(�u%�����Ur�A�Rd�f1*���e����A[=����b<+�/��Kt["�ŏKo.�3��}.O��,��GΠ��V/����ٙ�;+~���5�y���T��?�	>���Q�����%��,Td36i�φ��^�eIrT�'E5�-d�8,Q�c�Y��2�3�����P�9Trh}�i-��~�Y�T ����T=7��:֓��z���i -o�(7D�?���P}*>�o�t�U�<�E�mU��m����)�:?�=�����f#���g����d谣n~.�u�~��wش�3��6jGȉC9��̸������f>�����D��w�������GvKF��W2\V����DM��$�"8�A{��qm��g(D~Va��|��� s�*&0�q�c���E�Еz�2��٦١J9fᣌ> ��*~f��'0��ʘ��n}��9ߟ��傘A4��e�Y$�U�S�����z�h���dW�Pi�8�Wr�ɍ�]")\��"]�R�t��Y���ʎv��\�L�Xx]����4Џ2h��¾�^s�z6�������À�ܧ��,�
�~��z�m��/��Ѐ���ݧT�/*�XkSd�|���4	��GfwRφ>��a!TX��R�}$}𙃁z�O[ L��z���HP�;�C�����;������,�)_'O�, >����~���ߣ�~DL>�{m3��וo8�`�W"1��,\���ؘu��Ԃ��������F?eg�$g���=�&,��7P�M��?��̖��S+�-ҷ�u�qq�t/��gv���ɬ�[�a�j�1�I���C9*������P}�3X�7�����'��[k�h���B^�������T������*m����s(�[R�x:=�W�p�@����w���B,Y�`�
��+c�@3��fO����;�����aZ��΍����=�ڎ��3�* +쳁yJ�71D���&�!�̳�孔Ϝ$ߓ���{�k��(��Q�����;�-d��+j6�Bʇ�Kzd�8�%{q(�N�M�q��k8�nh)䟰		�Yز�n�{�j�����J]{���ohĢK�0w%t�_�E=�W�ѯ(��/�8��檭���Y����ڊ��.��t(��d*�<>��5Ө�a�A�� Z�[&�4�����c� �����J�%2�8��C<����ҝEHS#�j����Y ��֢�U#a56
� ^��l�~"�l�g3~��Da!�g���e��6��T�"A��[y��s�(���d�I�P��d:�a�!N�,�̀g�J���q{�!��H�9r��g��,G�0g�t�ȏ|��Ίh�p�$���6�qɅ⾖��ga��.
 -�f���p���ɍ@,��rv��:�����H����fY�h�8.��Yҏ�ͦ̑�u����L�?�~�U�C��R��R��ox�[	0�4o����8;s��B����<eZ���C����"���p��w,��ts��}�\>�ΐK�s��i㘘���f�o�4(���6�:��>Ж�J�����HX��y`�� 6�)ّ��]:�M\�'fJ[�9\�D��\����t'雷�:#���k���Rh`���V�I�d����e
��k��Y�B#�+������$��+�d��G�47�-|GA+SP��H1=�bݤ��ן�l�L�&�/�yl_ߕ�b�u^8k��� ��R�N��Tm}�l)ƶ��==���}<y�xt^���@lq����q8�B�M2����Y���tX��]{�/j��;n�c
z�7lX{�bcM��@yKڰ%��@R{�9!1kgJ2S7һ���I7:V�p�>8�S�����\�vZ!�2�WF%�g��֦�(MҹdT�t3Z�����<!%'���.��_�l���B�G϶��
���[�w��$1=7��;�׸d��2�$��"5��6xu �1���D g���S_��Lުy|c�{''��~�)8��_?h�6F�ڢI�O@������GSx%΄F:|u{+$�0e�m�a8w<�92���%2����������[,��hWg�����E�[7���}�N��z,��ѢZ[��T�ö0���M%���'[�w��v�H��s���R�b��`8��kɏ�*$�1*}ֵW�϶L&i������|-^❖��#�f��.�UuF@�� ���$����v���()��g�U#|�ߜ\��V��7'���U�Խc+6�Fʡ�(��Y�ׯ�G��	/�Q5��G٤maD:�P�R���\��d��=���,̵)�7�M\�+ʹ����1�@���#/��<�X൶��ׁہ�p��;�5�Rآ���#����Z�_X��b�w���J�Fߪ�VRۃ}yG}���[n<]5[h7ĉ�EӺR�d�1�jw%޲�b�q���S�T�+�0�yW���XZ?�KI�R/��s>e��'V���Su�/�I�_.��D}�oi��6zj��9l�<ܯ�?��lA+��椬Ba��g!�OL0�xnM$ �O����d�l��9�xVJ�[r���4��݈�.��jQǭ��y���fy�*~?��k%�tFI����EN;9�|ahaA��:��`46~*^�9m�V�gǞ%��JRR�h����M���|"�¥6p�j�I��<�O�w#�-�(�מp����%3��V��hq�xWj��|���.��@���T���ؒhE8��n��4��z%B�-��ʼ�O�0��u\�O���	 &햵�]�^N��=��h��΀P�$�MB뿠���'$�����C�-L4f�k"�*��.��]�GK|�SP���MV���g�~�X��]��W��U���8*�|��A�e���ٰn7�D�%�(ɇ#A�g��������1mP ~��_��HlT$�a��p�Q�p�ԩ����-�$��{E�î����B�y�aG����8��V��Ew��
��R:����U����R�H��Aj�d��q^���~���M�_2
��]d����si<�"nV�;ك����t�;L&�H�GU�}��4�@���te9�Z#f5�P�9/2��T�Yu[\ �̖KDr�����,��K�����֭)��0?��P�7a�xLsվ��.¼.�����v����Wv�@����W�'��A����0
��y�R�>*�u `y��vR<��A�ܥ�"{i
e��T���^Q{��,a�	1�6�
�%^���ؘC��7�a`�Ҫ�. G�B���#-q`D4&�x���N�0�g�Ȯ�B��؝���**���aب��8��9����d]�3�ڮ��j�;J♮���,h�*�U�mO�s�p)O����?�:�ud��P�<�����(�Q��(M�rmx�������KYj���n�����a���������l$���u�Ӓ.�dQ���t^]4,��'�{���P	�<΢/T��m����*��!�Y#���|E�
DWG%#yh����e�_t�wyG�J�xT�K~3�`��i 3|��5� �^�LE�7RSp�L��e�r���~S�H��\mސBe&\ʿ�qY�$��h�^��Χ�k�`��F.G������&!砚�x�]�ӻ񄹎V�j�t��W�|��sm������p~A�ջ�����
4Pt�n:��fu�j|#w8�A�x���'w+8�i��+:D�U�u84��q�_If8٥Jβ�rÄ!Y�%��?ށ/���Ewc�BC�o�:wS"c�*Ce��	h���av�#%�o�UK:�N�������������Z)?�>�Z�����B���o�j���~�1��n��3�����i��:jpC�G��f��<�[+�]k���[�O�mE�W�HϞ���q�v4����-���>{pB����l�w���X��?�#�N�{�<���U�Tl�?�\���8e��~�-y��D8��׵�O��W��
�;�Rn�`��vs*�G����R�Һ��#�c��҈���]����`Tm�d�M�(��Nn��~�HW_]C�s�j�ɦ(����O�ۄ�O��0܎��]�F�q�n������Ec;��0aN��-��F ��Y�곮�v���$M�*�w?-oի0���U�|:q��g�Ib�㷓m�>�z^��j���A's����1ۭhݶ��]���X;b�@��%�->n{!zvh��R��@��T��3$`�tgfNG
��W�wO���C:�Z�tL0��n=��Y!4ғ�m﹨jS��!��b.Y��P��kQ�%/>�V���F����8_%�5�7� ��d��*�j~ִ�j�e��*x|����(T�Ŭ�0s5T���psz��u�6��Xڙ�H?%v͌4Ū���-ߜ@v���g�nI�]*�P�%�m8v�DFJ1�Jm��?��AMY� �����H���cX:���G�Q�<�������2f�PK   ���XhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   ���X��НR5 �� /   images/52cc771c-8bcb-4758-820d-da79c3626c72.png�uT���>:��GApD�tH�CiP�D��;���i$����;��A�;�c��3|������οg���zY����{?���u_�u=C�e�����@��r�з AĨ���/�eo��[ί���|y�c \�u��v��~�~n4[�S�H�"��fo�7r2��pN+;��������E�(�$}��=ic�#$�؇��o?�W,i��O���I2�j��(2���qS�a2-�"ؘ�*���AS�I�ԋ�TV����/�����J�ߦ����� .�����������N����ÿ�/�׋�9��>�mP�t� b�������׏�4���+�$n��x��p�?w�ƃ��T����T����?S�oSY����&KV�M���"E�����b�����	������KJ�y0�p�_��3E�~�@Ҿ���@�g8,��?����������ۖ/SZ���+]be-�sQ��d"��AǑ�����f���\X�Mq����U� f ����h��h<�G���U�,l違��۫2\f(.'FK�npo�ד��!����z�@mU{,)����&�/IK��#`�z���Z��A�?.���c�KN�*��}������������_O���.n�sOX^Zm*s�uzc�N.��:)�5J���<Z�`�\���wR08�,�9��J=ux
�}�T��	�j��s�:$�!��u �Jl��)����u/����_ f�m�3�!�K����@����އf��S�ͪ��/�T��R�]�_yb��[��u�(Ij�CJ˭���]?]}�4��G�zE(���]Ә���4Q�,� �ި���'5T�iy����L2���jbeg�VC.�2z*C�����8�\��$q����o��T���a9����O&���
�jVk��4�����z��q�P�㽵�8�u�Uo?�*-�M5Lz=n�s��҄ bW:k~�D��Z\}L��nxm���Y>����g�h�:i��5��w/t��s�*����3V��ʖ(0&�����U�_�W�5T��TSv���w��ް:�xyS�ˡ��Gc[��6�&8:�`����ӧ�ri�����u/�Mz�+o~zj�vTM��9<����x�PG�!�A^!T�R�>&7��p�i0.A����i�����ш-J� !�9v\����� A���J�j���c�T���ݭ_-* qNXhI�r���R4�z �.&09��AA��m$o���ȅ(��d@Э9#O+�y�`	�%r��.���l���ӖǪ�|����R��lߑrա�T��ʁ��,�k(���$�٭���UOˑ���W.�ɻ��@���|���w�U)Rpt��}E9�d?aqi#�G�唻��^[��(�L�^J�/!A�G\!�:��v�FaR�ա���A�������7��1�؄�q���z���x�3P6�?A���]�|5WD����k4�0))�$%�- ��t�cI{��R|��h��/(��t{V���?1V���0�܌!�RȓyeK��yV�n�O��*��5M"<u?��2����i���b���X���#y܌+���b�5�1�&9��N�>���F6~=��,��"���sn9��$b�&�f�&��H����45�4Z#��2������/�w�{�/P�8<�Lz��4z��)�\.��={�˷ O�ӊY�M.aČ�x��n7᠍����)�^'��՗I�5o�x�5Gm�GYr���:�_�n���Mi-�q���V3i/`3��Vlڗj9=K���S�;h{p���L��k��&���D����;s�?F��~�+L�t�X���<�6b-�l��Q'���s�$���c�k�0L�x����x;�����yı����2d���2J�/�=/�=��0��773x���O���I�e �{�ol�L��9-��	�K�+���1��Q*)}��F�蚍M�5Ml�|����=k��������%�^>6^IU+�F7X��?�cޤ>4�Eb��(xT�@�tf����&VC��Ӝm|��sn���/��j�p���B.<�����ȥ��	��C��0d���]�{Ι2��ȳ#H�%�:B�E|��|����{>�ф�(�_na#������^��oܹ%�*.��oH�U�O̙B
l#H"�wb4)�4��b���a�����0�\��:��Ւ���W]�����3�L��P!Lr-�|�}gL��+�����h��V��PM�@3���=�tcCV�V�{�F��A_�Q@F�p���a-���Q��n�z�O���7ۂ:>R��K�8�O2S�lD���׺�ǻ��Kf1���k��Ή��݋��2�#��^����`�S�E16�����	���T	�h�#|� I^��:Q�zGG�IWV[�'а>�0d�fK<������3��,�݉3)raĹ~�>Nv޼��ո/7.3�ں�N��0�{�C�D>��E���or�DV3��1�'(ԾV�!�N5D���}rjƵN*r$��w|�3�>��P'�=p\Xb ���TR�<���~I�|�<�S5�&���oK |��̬��"�jk\�d7O"�Q�4����G�w+��7M� �$&�?��x-�FǺ���F=h	��lRN�����r�3�y_��Pƿ�������ܱzG�:��)Y�Ǔ[g��^#m:0t��Q��Eiح%E��T�������M�D� ��E��#A�U6��U�h�vP"%|�ߵUԎ�P�r��4P�O�������^*G��⎩9-�-�P䳛�~Uu����1t�A��y{���|�C+�[��(����7衳�Nr������"�wۏD��\��p���G�ʂT�,#\�[Q�$��h�
�����%P��f�_�P�J�������T>Ր86ϟ*� $�aR�Gr��mR�n��� �\���i��p��Lj�9US���i�4:�,?��6�����a������MWq�x`1�fJ�|�6����}Hd���s\_Gq�-6�	����L��3���4��ب1���(K�)�&_X��^��;Y��wI��6��ji��%Ƭa�∿�G0���"��R����g�ｅJ�E�	�y]��(-�I���h�`u�{���~x���F�������2�D`�D��^WߢJ}�Q�H���M����*�nN��[Q�0�c/���}��ߩ�p�-t-��jj�TԎ��2����n:# �?�%�6�_�|�h�~>�F���m�'&V�-3��N�Vư;a�n%\!"�H��7��Q);������S��S�����|��;>���Kt�	`3쎎N�Gx!@�Ky�&�m�d����������*�*���B��vh�h����o4%(�,/zRPжY'��=k����9*�3g���"��׻"��'�Q��0�? Kb�b�
8ZX�ƌ��(���G�2Ι<#�W��b*>g(p��z�c���A��O".�!F�)�@���5JJz^!Z� P��]\�;�!�f��NW ^�`=�X�Jg���K�U�ll���#l���\�x�URh�}�+ٸ�����֦���?���0�o�4[�qT����cM�!��7����|�,:��$���*�����(bt��R�w���+у�G����tn�.朏�mxۏ7k9���`t�Ph
@�go���Z���*��� \��N�,G���������g���]�0��+�������	okϳ�0<�op��Re[��d��~r�B�j��Y]ip)�r��-R�!�X��K�	:����m��Bj�,Y��r��=��������Oe�S���-�����Xs��U�w�^V��oRe����V)��)�O�vfa����¶��~�ʖ���2F4kEa2�ULD�)H�Gs�.#m��	�'|oQ�@O{�A����*�V�t=�+9��Q[�LM��n� ��K�n�۲6����. �<����y�w��l-j���Q0�^g{3Z|��A��E�*�3�< U�� ��R\�?����[�� �"�g>k����&�M z[��vp�䂤H:�nw�lOq[���\�g�������G����H�.
Y�C|��	�ު}�,�¶j��?jk��z��
����O)>�>�� <n;$H�,|��j5��z����k����0 ���l����CA��U�I�n�pw�Е���6�E\���s��[W����<?��=�7?���8V��u��zW���5�r���c&�q@���}����^�@z��ځ��)�m��V�S4|��ʲ¿�]�ud�E3��k;�R�;���j@�p��Wa�G@�\�1��aT4��hK'�zX_��-�a�#p�#�T���(�qWa�²i��uo^W\�Y�>�[��0����#��kp���~۷8��� p�H� ��}�SN��6_d(�����]���͐�Ҝ�}��y��
�]���5V�oܒ��Gn�_ɍa�!@��/F࿐Q�TQ5�H&�]�n�D�H Nj1bv�t�(�#�}���ΘIp���v<N8L2�\���Wd�-<?����yk&;����W�_S�;0}d�&�0���+|�N���޲���Gղ�
�ݣu�v�㵜���:��!@`�Ϡ�,x܌O���Eϖ��aKD)C PZt`+�w�2��y!m�g�g��C�ne��)?�A��H�>z-?������+����K�n�e���&��ȍ�-u�.a��kd�P8h��JC��;��J�n��l%ƶ%S���r�Z·�7���>����
����J�����gQpƘ��nK���i�^�;ޖ��̭&5B�Ϻ�7Aa0d��J�%a7����}�@��03Qw��ׇ���m��]��,`�8�7��/�Vns�	*.[�W�K������-ӏ���[�&5́*)�6Iq��k1G?�����Q?*5��'M��-�_�>�c�h	C��M��Q=�5?�*���1��I��}S^>�6�/�*�3��C��3����i�qFO8*��>_�p8��o0�����ƻ��R�/x�N+ɕ��ǚk�va���#�s$���6�?���x�p{��}��� 2���}2W��]z��q,`���x�����L͖���x`�L@�ğt
�"ị;H������kP:��C��b�x�8�h�lf��L��{��ǚ��=�?���O)1���bk��%��� ��> ��VZ��nO�h��ZT�2���s�]�\l��y��a��^R���7K�����F�;:��,���\�,��gyl ������ �&��#�E�{b�/q5�@I�e�"-���!iriJQao�T����[�Q���G���V�.R�G�r�����X+���
�(F����[�w!V�Ph$����e�+U��	�{�`+��r&	Y�P�/N�s
ν�����\��D5g��AM�"�$�����f�g5_��e��Cr��Y��&�Q�L��+y_���V�+a��'��BN����թ�<���_=#���2BWe!��.��r�k	d��߈2��frQ1��DB�O��+���3=��
��;�U�ȟ�k��f�s��IdF�U(��ڒ,��`�	��s��T;�
&d9B�"+���Y�O��9դ�-�:���y%���c�)��D�/!��z�^0��2��1Ƒ��<L�|��f��&�z��NF��Rzc�c��%����
��xջ����H`�6�x��CJ��Y>�aN�V �d��ҋ���2L��-2ڣ��Yk�o[r^G&��.������Ọ�����;�$�͋]�(J9*%�'��qҼl����hi����F ���Ҟ��D�k���V-󀓖��)`璈�Jqm돡��e��t����`w]�Ƚ����$K&ݒ�C�2: ď�[K��CDZ?��U�6�w4���m����֚�-���|D*�������G�0H`�|II'0�l~���2�+�2!�8A�14+�aY��<�;k@�R��L����_ :o_IB�������+|����~!)�,ٌ����a��y�����W�>�� �(���;��`g.�?'�3�GZ�k�O��9�P,Jw���v�fSO�cs9�O;e�V����?� �q��j<�a����U���Ռ�c�_vޖɳ9V��h�!P�dsE�"=r�z���l�a�ҳ؉BJj����R��f/��RtU�����zV��6�
K`&���>Z���sC8�H��ƒ� ���%F0�3��I?��{2�IC3��$>�t�������ߎB%�
�s��V���¨�U���n)	�Y�z����6/h�
����YC[�����������u6���Nb��Ĺ}��fPN����Ģ����K�֮��u�����Y2}ip�A��S�.cv5���a��������d�"~yo��^������N����Vr��D�F'���������t�5�c�%��rz��[��)�㚓Q�:�臼��I)��盄XO_H���۪���$�o�v��=�>����D3V�e���@�*{ai;��� @��H��f�zA����)����)��-�nQ��hH��tDKbDF.�>2Q�C��rU$�q��G����u�!M�_?Tt\Q�zFԞV���|���w9�n���;�A�J�nN{�0�"(@ b���K�9���o���������g���

"�ZI=Q�ɔ+y�#+@�D���gCJf�+��O^6�Zg��}w%�o*������(
��͎_X�_͙4���֢%��è����V�?93E��ӳj��Y�+o������w�Κ�K�"�Z�k!		%a�rk�z<ص��0�,���l��)�!Ҋ���+�8 ���� oO��m�!�#�9r��E���%�Er<�����Kw]�]����!['���b̏p�"�$W,��$����Y��=A������gg֟�'|��B+��%�({��׫%���`���犀���HdyN�]�xTJ\�J�8�Sav��v�@�K EM'���Z ������*���BƁ�ȷ����K�)�.�zVjj�o��KX�
dM���r=j�	����oڹŵ� 1p1d�t����v�����K�!�C���6�e����,3ӭ�;�o���6�����0!R����x�pX����KZ~-:��+���N��*��j�w��E�>q�,%�jw�T�(����9��J���6�1;u��٫:��:��@a ��֎0�&#Z�#�ֹ-�%�k{��ә���t����p��v4��g���_�e�+ ]�xXc�-t��rs_�i@�;��h�:_k*�۠[Z�uԱ��gl��d����R������k7��2�ohTf-�xD���ki�����l]���PY�`Uз�3����Z��~�ZG����V����ٗ���V5�ƶP#[O�q��o S�KP�f��L��A �~�k.:���y"]���2

X zuD�8��g��R��$�JZ�BfF�T�;����l-��`m�΂�9��&��F��	O}����|���Жm���^�F���C��B,��BY��u��s|wGL.��(E�m�
��XE���㩓�ψnR�m����)�:;޾jn�r�2@�lcG��߳�G�:�F�J-�:6x�/�p����m|��pXf��x�hb�đ�q##�uY�h�H�ӋګAbe3��h����1xw��bӞ����n ��Ӟ�؝\6�K|w���8�EEqq+���
l/C��lx �nߖ����ɨ9o��R����+��6�Q�-�H�o�
VMQ�&�:���k�p/JK���@m؊r=y�~�a��Ү�)1��QKC���h��?�F ���ϔ��	�LXA�8
 �K�)� J(��֠�/���H�\-�c�}.f�,�
�8���#]ӰV¾�[�E*2���?��4�j�)��&H�S$�6@=�X��0��-Z���}��rgE������d�����"��h����y��xQ%t��`�Q�v�(���m���+�Q __�N,}��ta=P6��$"���pC���}���-����F_&�(`0�g��.fE�����J|��Ք]�.�N;YW��O{��1��mL�_�Zwڔ ��׽.k�������/�����+q�mPC(+���^rHK���} �%)���Y�у~Z��l2tm|/!�B4�zA^9Y�LlP��<[���8�,7N�)+�a&�b��t���\�8�L���﬇����b7[g��N.�<��m��ϧ������υ�N-u��6��{���X3Z徤�����n���Bj����qt��E�l�]Q�.{.OjW����bC��Fp����VC���&��XX�ǩ�q�����%��~b��:��p@W�d�6�I�cR��Cb��W���Z	J��BHi�~l�v��Ka�}�JA��@Q�?p&`���͓��eR�>�D��1�0�V����PoH���F�r�@�B�l�x��`�^����"��٦2X������7c��$'�jA��g�i�#L٬ˉ΀3�MQ��!�՜@
�׏�$I}}G�H6e0����B	��s0x7���c��v?ĸw��D���{5K��hO��u,�nL���l����| ǧZ�Y���j�����ȸoݖ�hc�y-�e%��i��ޫ�˽픐��}�e&m��Y1!����4Tx��i�2�12Jut<���z�l5�6���,䆠���h�����;�T�*��xU\lw^)^_U_�P˲����/tc���އ}]�E�mm	�_(~��3�{�g�\��B��Ӓ;��j���Լ<&{	�"�0 �!�A?�7�x/>s�&Ch
��Rq���ZFA�H�7{'��X�E��h�Z�
��H�zZ0v�װ!7A����S�/����`��U^$��la�$Q�1y���g�Щ�M�1�>�������)�)-��$i��hBբ}%�n�~X.]���o����U!g�w5�$1\:ɳ����d��y�Ss
	�{���秬���w�L"a��˩����N��ƭq�����iO��w?C��Ro��9w����G�Bd�}`���O��ｍ&�� �f~��Q���O�=���K|����W�ܢ���+�+���n�/bCw*�:��_�FP�ǲ�����H:#�1����j�st����Nd�_�$�$�a�,@�ݽ�њ){�>OҽR5��mw��Q����Z2��2�B.����S�X�#y�r?>f��wj����|>��a���&P��@c$�Ux��`�|��{pM�`�i�eeA�Ƌ���*�	�15h9�0�&���w,��$�Qo4'�yYV/%`���N�d�2�u�f`�Ŷ��ö����I�s4yl'�CD�T�Q���1T�l�;�h ��?���E5IQ�6f�c"�n�w�i)�<�QKEm�xrE���2a�ecP�2��jX�ƽ1��=�9k�THJ��l�*�-�bX�Ҳ6 ��gA�����Y�m%�n�����0|��e��� �	2)�$jh��+��ɠ�l������Ѐ6���zV��
:��{&�;D7�AM)�E�:~A��>�z4�-�-ǸY�VTn<��ZrA�.��#r#ƴ!n� ~V�Л#_�_ޘ�r�!w�q���5|�\[�^�^؈�L�u�=��k�'�`��pe��
�[�X&����+��O{�я�}t��!1�=�}c�"�v�bln���3��j�a����`�˖/�?lt�'��'�a�N���a����~��:�)!�b�o{ϸ��`[5��<XQ}J��׈7��<�H�R,b�|x�R���p7ϴ���\z3�b�kʄh�3}�C��8�>J>4�#��������c�mO�UK�S��g��}�	�@���mȱ�QU��"w'�f9!�:AS�2:�qΡ�l+����Ǝ�f S��N'ZoЋ��·f��v�5^�Σ���L��R[�њTi��[R�v�b~�EW�K�g�����Y���ղȾE�׀��'�r�Vy���������"K���`I^w���'񄋦�5����S���B��n�T��B�m��.��虚��m=��:�E3�}���{���{m)u?�7A�.�p��o�n>i��OJ��M�L)�l��#;�2+(=-#{R�>҈t)�,��Co�A�֡SV{�"J��FP���*�jK)��hz���sH���2)��T�CX���W���k�ݻ����VR�;��N��m�����Z/s�A����*�#��w�İl�^pq�w>�!b���3�������6b3,q�2[}T�Z����nP4�?\A�����7{�h�Z��B�x�%���w*�K{�ߺL�t�Y h��d��u�7�q���fV��@�yG�\^o���=��3<��'�MQ�d&�C��໒˼sEy��d�j]('��_����Hc8b��ԥrzхפ^�ѣ��A��֊��c_��&eDR���A�N�.���ͥ �ZZS>	�)w��~��o�͐��c��ӵA�G��>���{���m|�c�`h����@�A�����!־��e�y!αH[��)q�����I7���D��;>	Mp������o#��LZ�j"&]v+��ѳ%��
S�&�
�`+h�(����/[����7��g�/d������uPt��V��Wb����W��;��jA?�>���a���&S�7�vaͣo33!}�B�˾���L>���2ϰC�'|@ �+N�(�Fy�V'�{�ٚ�I8�>Dk�.���JM�E'�����9�#~�ƶĦA�J�Ge-Й�.��ޯ���=����}�����]�E�N��`�X���U1��¤��Ԛ����F/nSe���i<����x���u�yDx͞��ή�wOJ���+
�c��ӓR����#h��\��uT�l�4�q�|l���~-���eh%%~�[փ��8Q��TUx���:�<�-��:c]v�����b&U�z������4�L�s�t�ߧ{�;9��x\�`H�̖�n��� 9�mYo�h-�=�~MfV���K�
���I�5��9ƦC�ώwhƿ��[-����h��b��o}���cؾ�+ezb:u����ϟi`��$�.�Eh�����PX㚌��q���x�����ՠ�9��PT��D5Dwլ���heJ1��$�%UR�ZK~�`����IG���U�[	��I��f	>V�?����Ͷ;l6�E��KpI�Y�o���5�p����ﲹ�30�1ש9s���*��n�׏��$U��gY����c��xc���5��e[�**i���[��k����-L��Bu�\T�:��Z�Q�xi9��Xd^@�s���N�,��5�I ��7O�̻_k1�н'4A	5q���q�8�vc]~�LT�@�p{��������I������/���L�kA��i9����l�V��t� $:�-��C���Υ��p}7A3��_=-=T<N�!���K�����]��y6�
׶u]�������F�)��z2���YZ�@�~f�L������P��B10�H��`w�K���v����	�)W͙�,R��>����Q�Eܩß�Od�o����E�����!=��X6�7P���&+W懗��%���n9z��V@~���:j�C��\j��Aְ��Xx�{���)�� ]��ȱX҄]$���Ɲ�(�(��5������M.�d�_C��� ���[e#�TDW�~�C�{��y&�(ө��Mr��#/��8u�g&9�8�?Xv����FIun����~�|�ψ~E���S��7��-��6K������ޅnwv4�I���ª{i%ֳL=��)%j���^z����Y�t�͞A U3���k�p�?p/�����٠7��j�)|[	>]�DD�tx�;��/L� u��W��oݞ����(*(xKBx�-PF�}d�uC����@^s��1]��EH�5��_���mQ��,���z��X�Y��M����?��_��Jߒm�C}{�=O�e򾥽@qL�-6�6.QO0-[�,[i�7���Il�TM9=��3:`�.I��6,���nҞf�F_p>�̆��Ӈ��[Uf�=�cEڞ]��m�/q�=�R�Q�]��`[���׆�*���.~xK�2�ga�x�U0F�a��r��h����a�<:[l�Q��c&?��)�>��0�cj�h|Q�FM8���y��OPFu�O�4l.�Y
mU�ۏm�N�)�I��I��>�|ϫ �wR�D���P��<]G�	O9�OΚVEi̞-���9?��&��X�R��b�D���g�ު\�/aX�7�X)�.��'�?�Zk-�\+(I�|����\f&��w`$�~%/���R���%����c����(�ĳ�r�1s�	�΍~�!Vӌ�q��S��9Ǆ���:0yq��M���
�`"j;m�O���_.�<�pX�ѳW	�:�h�����-rd��N9%�'hD��b����:��n}A��(e"�N>>z&k���ϊ�"&o9�9�\����%k� �S��^T&��P�����X=U[��Ng�@�OFs�=�Kt3�i�B�e2NH��[*�׏w�sD?��Z:z_�5�-�n��%�{jZaC���Vybt"]|�����*ذ�"���9���q~�^!A��NcX�żW���!�e��4v�Y�/�K�H�א���¸w�����m�l7����į�/z�*!��J�8N�35��ŧ;�\�S#n�V@/��$���!N"|^T&G�|R�u����q�$����A�V��Dǈ��V�c`7n�[��P�΀�xe2�;}��(�ֿ�����h��W� �=_��ӄ��xF��"_ګ^�%Bx��M�0=a���Q�lNE&����H�᭦ᕑ��_��Dn��~�����[s9��K�l�����Z^��q�D%f���%�e�[��>�I�_��\yǿ/���=1��cb�Xm�,�_5����3uP���7�83�uTK*}d�W��/p|�6��/y�˳'�Ю����gO�m�q�����~VA�Z�ݦ�񑑍��2b��@_����a�r+CZm�s�U�Ã�є���6����������zk}!���2>���ӀUN�^�͙ݼ6uk������B��Qr�SK��Z�l5���l8kV;�p3۠�ؚY���.��@��;_��x������ET�+_�F��&^�.E�6SEK����3�#�i<���o�&�	L|��2W3�1�_D{˰/�{C�s�B��[����p���<�=I̛��e|̭a�[ڽ�!��ȷ�b���;�a���[��?��,@���;�kI�,%)��W�9~��i�_�
Y�L�885K��ي#|a�0�
���%Co[ �j;�L�:J�$��mX���Q8���ʟ����[��P���u��1�Y �rc��d�}mP2G�7���3)���CM�~J6uc#]���	d��@�5��8
@A-e��z9�s���?�)O�X��zut�)3<�i�Ŝ��Ηa�3���٘V'=�o~�SL���y��[U����{fc|�jMxmD���~�I"1�$_�S{Nd�R��ۮ7��8؟��2:Ͻ���@g���Չ�G-6!&F�J��y�@nA�:�)�<V>o��*u�Ҝ��B�]c�nA��˞.~���	�jDH1F*h�����jv�]�YZ<ғⴷ�\��u�;v��ļ�&���Rm�V̯gdĠP/��[L�sW{�Z/�*3g�W��`����V"ƞ^�K旲������F��l�IMPJ�w��̈́���W|g~����N�(�cB�me�| ��vpDqn+��=���C���$S���r�}��ֆ�c�J� !Ը"����ک������$$!>��@�SJ�c��ң�d<��ĥpL��m�Sk`�Z�:��J�k���n�]P��������*����lั5Vn\�q�^�Z~d����8A;�Ŷ��ix��{biGk�Ab���,x>&f��4�Y*RՅ����x������J�Ŷ��9��Q��=� Џ���tM�����wA~7�1�����o/�1Y����I=��:��v�O�$F�\xˋ���͘zn����Ъ�d���{�|���5�⧹^�R�x$��p��m��K>�\y�x&IW�	JV�������6�u}�VpÅ��"W�����!s�_�1�C�0�!R��k�r
cU�ϒU,q��Sѱ����~����|�����dR��^�۵�K�oUaK=Ht����}�$��w6�@q��Ux'>ƽ��q¬�ӽ�"oBdG��F[��c��������0)(�K,D��{�ǰ�^�u������b��s��(�M�G�d�\����M֝�<&�F9����wd����^�ϸ`$S�8�ҦU�I�N���^�H�`�O�R���;2g}1���}��|�w�m���*e�(���A�/ \2��_cD��$+|�o�d	�Э���@ ���t\{ ��-`	 ��;8bMQ�[ۀ�z���)�w��V���|��}|u����8^�eJ�y��ܟw��u����v��yY���*
�8%n�s�|_{���U��`TD�pZUQU��VD����wZ�k�9*����ހ8i���K+s^��"�A�� 0�
,9�5�����`c���a��/�<i3^!{(�v��6�G�}��c��n,��R��B��;�Ѭl8DQo}�YAjC@��m�6t,e�f����5��V��eM�D��^�^���E?z�g	�@z��6*_���\)s�^K�*�z��?�6�+a��
8�>��;]�������(�4�i�@b��]�䷖x�-?ޡ���<}<���2jab�Q������� �J&@x�lGz�`S�Z?��I�3^2��:���U��F�?jE�lz�^j����ѭ��Ќ� ��2��,k~5>^�,7��� �Z��aG��"AV�Ӊ��|�pE���,�u�]�
? �k��?: �36^1ɽ?�)w�g3$-����]hHR����#;�_> �xx Jg�+.�zn�s�ӎa7��0D�|�� �`��.�a (�  9=Z<Ā�l!�H�S�WwF����a�t|�Ы�z;5��+��-oqCo3EϹ�Bo�6��T�vD�(Tzųɖvx*�<E-�^�S�tor�\�[h%�!m�"���u��y�� �l�-ڭ��ҵ�M�W�g�#@��ֺG|NY |N�N����9t�.\֝�Rt8!�A����7x��#���Y�R�~!_�C�1U]�	P����Z%�!D�[Cɶ~�|t���&�b����X�j��&��	���V��eVS��6}ha��۱@�D0�ݑi 4ʟE1[���Jԙ\�|���$zۯ��筣u`^�ya4���Ʈ��c��h}���p���m���̘�L�nh�_��"|$5z���������������󵹕�1�@�u�L���@`D +7iՖ=����T7|f��`��ęj/��t-7��<�/��m<�3�y���@b���DO~{���g�M��ͮ�L���Qk�J^=�U&�}:2�k�dp���`��8��-�KJ?djc�����m3G7����@.�_�X9d�č�q�l��j��23�"���zc8���y�(��o�� j~�!�ɧ&�j	����5�7�/j{G)�׹�\/wZ���g񯬶
�V,�z�F
�*u�͒�m��/�ت\ y��0�M���j�b~9�2@b���F���� n�04K�u�#�Uo" �F*����UMe��� q.B�C�m�:Cx3��@��[/��,Z��ٟ� ��F�I�� � YyJ$�"`�
Ck2^�(#]]_R��O�p5̛V%D:S�����X�-�c93>W�-,3�;FZ�1��{5YLI:�!� �r����
:MѱÕ�.?D6v��13<�ù HgPFk�}
4�o�	1PW����ǹ��8�'�vd�]&5�4�=~�c�W�"$���&h�����+��+[�Cv���l�t��нXW�ֽϖ�}�j��`3��+�/E��=������P�B��~:�>�Ѽ�{��-���N]���x�0��	�� ?>A&��m��Vk7�(���S��
����j����>v��0��X�$����qU�w�^��?#l��Wn�� Pm@�ۺ��H�%$}���z�tȂ 1ڱY�}l���s��22T�����5�� hô�V�K?n��k9���\����b{9�=��L�X1`����>pe�&��@_O�),e�qw�k�ҸO�Ⓖ�v�57�����]#�Z���9<>9yz��#�O!����j�+�K7�����o��hz����6Igz���Ԕ%�mp�g��Sj t���� �o���5�m;�:}�V)��j�����n0W��t�!�Ȫ���l�z-��y��U��$��`� ��{Pm���[=����*�RF��Z��$��b�Tb����q
�4��Ry�^��&J>�q�7z���/@48B��8����O �(�@0�����Ҳs^KG/ 2�q9��2k\����Ŕ�[~�ó�%	*�s�r�{�u��ά�hMb�a�҉h١�k�-���J��ȟV�ٟ� ,k��&�G�����&�6}C�}fo�0��5�#s�i/�G�����2�f��դ�w�^�O�#xmx�ƛ-|]S�ұ��@�C+��uq��p��PJ3f3�ڎq=V$�Pimf����g7�
�Hm�$)ۗ�T�j#yߒ�����$�/�{U]������M��6�����x@,��ߟ䑨��c�	ڿ����"�[����ﮕ�l~�����:p�G���R�
��E������.�#�b��ꯨkС��@U���b���L҅`p.l���;�<�Q��"�nx3#�kKq���#�C'��7�[�z�s���?�W��Srh��a�GAf�����j����QD% ���Hu	)�%��ӤA�CE������a萘�c`��ټ���g�zV��׳eb�'�#��C�V���%ti�c"8l�w�Us�\)T�W�Lj�e@��8l5�z�>:�O�IP�e5@6֙�ww���$�U������L�C�|x�Đ����q;�E� �B{�O�~-,�g�s����|/e"�S��1B����*eLvD�a���9�4i6�Cʤ�/�j�@vpz>RIa�ޖ���0���.��/���O2|Y�c���B^�w�7{����A_L�"���L��&m������ZMa���	�J�Pb�!���um?R��o�.�����o��9�&��;���Zk�3��g��C֜j��"��@w���b��p�"�*�ST�O��],#��җ��ZI<Ix5��١���7��8w���O�ki�x�!�1K����`G��!	���S�#7>����妢�w��d� pl�����q�HzS�����qdk��=<E/��עBg��S�k��:�dk	����'Q|�Ou:�{���ݑ��˳1:�#Mx�0�����󹤭��s]$ޯ��-����bI�ϗ*Bax��IKBP�P��w��7!�2�s���ե��ѷ��_&��T�v��ՍC����7��"$�g�QW N�ON#|)۠x^���9L@����ό�9��>=�~���"�&2j�E��͗c��=;G� }䫩��:H�u�M��������w�:����9�G�DŴ�zS��M��8 �
d�
�W�� ���L�u��p2��8k�V�Ua���� E��o��������]-/(_ �;*f�:�x���$1����>E��J���D*�C�4��� *�_(�a.ں	�_��<2=/�4Ȕнt7'���q+���R��T�L��+��>�f���K@WS}+&�,���r'�Ջ.�ڭ-j���対]�x \�M��om��/�?tD��Ҵ�a�T2������G��F�����aC��������9�������<�����|��C������~�WW�*���63���W��jFR���T�[!�}��0�`� ����p���=�W:�M�j��V�J))>�x�s�������ѕ����8)/H�� Kc�����ξH������bR���#.Gui����x��"�/��)�����q����U��6���]XFo���CP���f"��~��=���щ��e�so�"J= )�Yq��n�'&��C��������/U�8�������ѷM����]��b;y��K{���D�4�l1��z�5U@â?>�t�$�!�Z"��毖��u�s�o�Ju!� `\.��X3@��e'y�姀�6�C�@���\��kL���ր̃V��].&���d��{��kꘗ��1<11Jk@3��|�ƌXK�%̊ڪ�.ꈺV��>'�eFn��=���$A���T��c�:㰜���=�֭Qp��i'C����l�]BRcQ6
��v�J&��k�YΛ�������!	|�@�9��X��4Kį���@�����s�����- �d��d(�0\ȕ}bc3�+��z{/��#���.�o_�:_a6H�WY1���"V�����$��gD�g�pݥ��O��`��6?��$hթ���w��Ϫ'$ߡë��q.=���Y�k��l�g.RG^�EN��n;䀍W�K$�(�IUg)}"�'@5Aq"ȍi�ٴ4�bU�X��������E,�F��j��,���J�}q��gM:�Q���U�_��;�h��pՂ�r��~��;�t�I��J��z����x@,�Xsn�I�0G�7�1!�H�]�%z#��
2e�!Y�W�Y,$Iy����7.��Pb�R��Fmjq�UۺmVmH��t��k4����6�� [�0~��][�758x+^���U�9_H,�;5'E]w��㙘�p��ԇ���ۍs�� ��n����5��N�J���ԟ���7M�u����z���~\@�+��')�^��^�/��P�6��J$a/��ҺGآ�c`�a�6���#�m�E���k�_g���u��=;��~7�#�
�b ��JR{;nNf6
L"&u��@H�E��`���
/qHLQ�
3iZ�C��P9�\J��d�vK�GE�oes�k�Ĝ��NGωB�D�נl.d�=�����?�e�����= �^���O�V�d�7�:�I���oU�|eo�̮4�\��|�U�w��'���_4u��ؓO��E�;=��~M	q RA���?�'=�!���`�S��wR��bM���\F�G%���X�yxYp��Ӓ�I�xU�Z
�\^����Z��Q�5���'8��hh�����J��0�^oڲ��$�y����hrK����^���e��ྮ���M	t��.�PA�RjY�[/�־�̜.���;H4-g)�`v�b��YP���L0�����ĳ�[���&,��1s_��]��Uo�s�@ۦ�f
�ߩ�g� jQ,����j����Jsԕr�7��< �1�����4�(�.�Z������lj	=���\X�[]�)��T^�H�L'c�?�|6Il+c�`(��x`ò�����	�����F|J跐��p�j��x��A%<_�e���CE����;)`Pv���#4PZ��������c5��y�V4R"����Iq��饎���#������;V� �0��!u�^`E�r|*M�moc}�ը5�?@���g����'V��� �ʽ�mm�E6fe�r�S ��2-�d�oަD�.�6�~�R0�,�F�
��eq�0IK�b���V�������y��:�p���3��|�Q
`���c��6]�t�k�W�\�W%��A����B�3�+{r�E傧�������P���o\ QD^��3ɭ��ݘe��9 �(VOH�vބ�l�J'�6��������Q�Qs}�R �c|��6ю���N#�U�>�V���P���k�G�r�◻���K�M��`����ڳ#� ����mx=��sQ�j���?΄�7��hu�.�A&Z�=�K�j;73&N�T*�:�4{�̖�~;�_Bq������ò��a*��審X�DA��N��Ԃp�G��8���@���fX	�f)���!�3��p:��9��[,��!�JW��xpq����ǉ2�ne��an����1�>Y�ܓ~k_�ɹ�C�D�@o����*��.�5ww�q��
CZS�i݋������l��'�PP�1�i]l�C/T��.0�4a��"��>E�Җvs�ƺ�|���_}S�3���X�݁7���Z���x����֩�dU;n(����%�<�p�T!>y��f*<�gO�О��3ßkMz�;:A���{�ۓ��{^NuF3��gluN�%_�e��F���߆�W<������v��1�M�1�>��k�ts1�3U�M����ZP)X���,�:`y��i�����U�q�U�M��a�����4��G��J���ӌW��]��y� �.o���m6�D�G��"�n�^mX|�_�Z�5�x�ރ)���w �[��5��~�rs<K� �����}ÏzZ�΋�Ğ���kkd4���*~��?�[��9%��j��������5�٪RK F3g�B;�p������.WRj١�JNƨwŗ<6Y�IS�{�D��J	{�A�����/ډoW�hbc�O���Ԫ���ݦ�;jRJ�� �Ei����5�]��!�{�s�ݚ��
a��W�,~��6��ԇ_�l�?��_2-��pou� ͼ�.����W�R?�v�gw�~&�&�}<���:��#�p(��\*�!`ۊ��c;�c�\�6"�-^��`���}e/��`��s+�-���O���ձ��`�~����;ѕ�/�5�@�s�Z��q�8y����<`�G���b!��'n�MB�w�ٺ�q��^!�ZS*ɋ�����f�J���Y:��w�&Y�Ք���>�p:�|���Iמ�5����m{����H�t���a59�.(,���|p��7	�F��$�%L*�xw?�x�0��V�B,qݺ��BIJ��#�:I<�xi���M�pR�v�������Z��3�Pn��m�rlt���6�'�|����TAv�܇J3�W]f&?<���틧������y�Mhz�O�P�궡��gW�����5��3���@±��A���o6�6��)�H^�t��m�v�Mk�4�W	��U�qDJ��TE��k^�m����d@��*�RMS�t�|�C��!
,5���� �"����uPt�/?�"�;�G*'^&�X?���Uv���n��J�9 �W�dui��Ο����o�7$M��Y�ʤ���j����{9 ��*�܍�uYA��}��f�e>��g{�A���,�L�AR��z4)6p��W��_@g���u&�]p8$�|K�c1~�#���&"�؀p���J�,��nQa�Z,��~�:gZR���|�~5Y�c֥�[�"L ����fpRyW�l1�a�0�,ITB�]`��1�|���e�y>��d���qw\{�F�?��]u�s2t+�����AQ������j�C����O�����M�7f_�Cfa��d��M��E�%l�-����(���{���Д�~($R� �|/޹ы7d�	<�:�~p�~��e�>{4�ָ]=	���0�`�p/�k``i��w�Vd{w�쎨5!�7�q�4�W����$�]��p��Iv�&��0,#f��0���\�!W�q�O�_ϳ�%��>� �xP�����,e3x�Y���~�JQ��5?]u�B�c9�5�������W��))�J�qڹ�?X4�gX��F�Mk;K�U���?[�+D�o�R�jZ��Y���+�����������BJ#�'\SS.+��ύ�4i,��b�\�B�$'	f���5^�p�H�[6��#q��i@�h�݉`���;�N�U�h��%����'��S��k�'I�ѹ#�����9E��zT�E�u��1U�L���v哅k�
�$޲���қ�)<�b������ScR��q�W<�
��|���$�������vGJ��/�lU`�<o��
 �l��ζ���']���hh+.�'��Fm��&Ɣ
���ʟ��L!hZub������v�K���f�'QAb����5��7Ԝ@�?b��+��?�_~����F�AZa���b|������:I�9e������曏��0q�ߤLy�P����YT��a�Y>qeZ*�=�I��Ƞ9������Q�@�.�2�Q4}Dt*�����zc��j��X�@j?m.ȏ�)���E��"c ݦ����'�P
 �J)nD��a�'��L&;����j��m��p����T��<JtI�}_QU���l�0�}D� ��!��>�� zܴ���hX&��i����v)�rן�V@��t�|n5��vk6�M���]���אں\"����˚�"Lݍ�L0m���������=/E�\�ܖ?�3�?w�:���%}�5�R�L�oR!�3��<X�����a8�5�=���q�����Xm���(<h9ͤm���d��''u�
?Zw�
D����n��j����-�� ��}i� �u*ӵ�����<���;�a+ҋ���昴�	 �D@仓ؙ?�F�#��7Mq<N��Н*����y�+��R��X�Qv��c��R���k9�`/�G
�G6�D�2"�NZ��D�D�5T%�6��қ��A��x��x��vv��p���"7�
��{I���g��vo�q+�6/���T���Fs{�;VG� ���v��ݿ(��,`U[�a¿j!��X�y��$aݼqCej������������������eq�᧸����R�>�$.�&$Sw!�W���v���]�g:W9��]�;6{�Y5��������c����Cfk���Q���ɜ4�VKX h���F���3LT�d+̼���u��O:�~<�[�\d*ڹlRؘ'N�$��j�xv��r<��.�x��W�W�+o�2~6�U�"�Q���@��V�-:��-P
�ծ�����w!�{�=��ߢ +���	a�y���.�u� Nn���`�CQ2�@�����PR�=��h�u��oq���=�·��}�ڌ*����.�8�3'�Us ?1}]%ַ�UD���&	�������Z�7����0�Y��p���.�� ��$�v�zZ�3K�	�4�q�vF͘�R)���6����t���A����D �����m�^Q9x��Zr��<$���.�m�{�hbw�f|Fi'8k��l�7�����T��HZD2�v�y���K���a�D'�O�}+�d-e��N55πO^�T�9�.�u��C��Ȓ(6{��ߖr��y����X*(���o�ʣ&��`���hK�A�a8�����9ňC%�Y�#�%~��,^����H�K���󂖕���=U�2�����f�&;o\O)�
\��V�����l�Rm�D��i*����_�dn�O/M�NHDy�ރ�g�ʪ_1��~�{ŗ���D�,<���ހp7�~������b�ѥ&ƿ:�^K�;��;I���GL�)���;��l2 �>h	��^<�_�Ǌ?��<�nv?8�h�	 ��)�ܳ;I���t�Ip8��n2��l��K5��c�M��l��r:��$�����/<:lͩ��:��3?���	�+�1I#�q�+OZyh,���|�2*f��B4&S����U+A3�������#&��K��!I;-2��Xk/Y�?��,,c<~��P��N�����g�Jߋ�W�� _�۪����0�^���������s{2ԉ�6��Yx�B���u�3������U�>��")^����߻P6v�w�(�gq�����;٢閖�+U�g��0�6�`%n�b��� �BS�pIд/T��	0��q�Eq,O�6�P�����2��Ŷ�4�ڸ���F��o
?�xgąT���jT�l7���M�8|hZ��cw�
nw�$ou6�w����>΋ �g!���?uU�&k�f�6Z��n-�s_�MOƃ��_Q}���Ԇ_q�2���M���c0KT/t���9�J����ܨ� n�� Wqt�$C�Ѻ��@�ä�T��ەRf	�����R�����Ei=����䡥�Kx[Q면Y`�쨬"��*L|k۔��N��۹p�}̬^�$5�1��}`��>��5u���K�`�j�+���;���S��} ��N�V5�]���7F%jNX&��Ǟx�����.�v���lX�c���:=���J�ܧ����4A7��S�*"��YHd� /�j@9��Ϧ~g�M��2�j���Ϯ�Z�\��ܚ�\�Aq��bP*A��n�e���$�mQ���߱^N����JR}\Ld	"�-�yr���,�+5c����ch�~�@ �n�'����o!s���v�����ȯd_���������na��� #��;M��;����o>����e^��sd�A�Ұ�!�|�o�_���Tßr�7��Mʝ��
KgJo#A����}}3v�u�OF�J7�����M���� ��`�ΩR@⹧��e�b��^��F?��jL�7��D��S?B�m��Vq|�K_L=������`Y�x����2r�q�l�:��-<d3�Ld��J���o?0�5I��	~�o)����YfL���.A8��(�w��s�x`��nmx�����x�����{��m�k�K�L�1���խ�f��M���ժ���H�*�ݩ���uV��8:��F�!�Ӭ<)*���K���4n��o@{��dԎ���I�3��|-[?��� �����Oٚ���^�>b;�c`j�yW�!߭#�aL��i˔�k��jW'v���S�X�B��SP��"�ͳ]��y*�p��Yڐeè���
�AfN���
�����[�>tZP���~W���i�
~��~�4�CG�����N�ܸ��mg`����>y8v��K%{S��ik��$p��%��W�5����������A�d�LĚX�y�g�?܋�������c���c:'�a;�6]�(ŗd�?�L+�&����^�����8?���=�W��zyJ����T�w���k���P0a-{-�Vm����hU�Um�ohjqF� �Y{�Y���y(����0Nۦ��Oϼq|���+ǥ�O���o�UӔ�8�J�����"�'��8����� �����;θ˃Ѳ���]E�}���#g����&*I��7�a�	%���c?��/����S.گ^L�hę"YhY�oܔ�2����g�F��0L�LX���ag���������t�Q��t�f�m;�j�˷W�x`�W��P4"oc����~��CT'-M�`Y�Ф���7�O�ߝzA��i�����!|�����'?v�lؙ��dr�D�"���t
�;G��QċW��Q�s���_M1�x�P�ӿ�S?��b�x��z�qzm�ӣ�PfR�J��$�a����~S��E��L�Z��M���n�E�s���l�G5���)����DuHm�J@B����:N^�Pޘ"���>8f	�F�������oM��\c��	�.�Ac�f��G��m�l�吤H���X����ܼkpU'��1����ze&��{
�����w�@�/��wa��t�`��>+����Z'���`U��m����f/���D�u�"�Z��s�*p~�ϱ��/"Y���ސi���u�
A�-��u��;�'����ad��˯>��P�!���J�}ۀ��$Y_�m��k6)�-�Aua,5=26�*��A�����ĥ���>�a��Ǎ��E�+�u��l6�M���i� c#�F
:iI������Ք���hzN ��1	���9��!"���2�_�����H�c`�iM0{�7��Ja����?s��+M�m��@�S���vߘb��)��	Aggt. 5�WX�@?Y7�~��KH,�zd*KZ|�x��|O��p������cM%7sN�)��9�sϗaA�K���)��y���7�H��%9e�e�	�lL�ǳ��S�F��sළ��h}���k �ܹ���_�^�+�e@)�(K�8�1�������^\�]��U�m���F�w�d�|B��M�0��D�����(}c$11%^Y����WWc��a\֡��RҽM�J�!�m'����{��Q2�XWW���`���ف[���ON�Z'�8�*W5�L0�d���tq>���o@�@��fff�I��p���!o�3�
*ۍ��)A}X���b����,_���~Cݛ����ܤ�r��/�o�@j5���lJ,���zG�n����.T���r����0�G���F�Lmޜ���f'�u�u?<�h[L�O��8
����\{�p�t50��K/�w��D��� L�'�OA�� \��o�6�'�#��ͽ�P^��]����ng����U�r�z�c@������`�O��j
�`�?_RW�ʼ#���5z��y ��H�O�$����b��_D+'_��	����)	'@0�IAh%����B!���� �7�$R��rԕ
*Pob�ݡR�� �|�fl�=�.(��x��r�C�d]�0:a�::��/���i��H�is��s#'�AM�E�Ӛ?����4e���[���HF��#C���
�s���A񤈏^ϲ;�u��̊���t��6�~T�
W}��	�O�N����M�s�6e�R�1Px��
�x	��a��$�x"��e� @#Y�*(N�昷iZP���l��v�u�[���ȖN�Z�'�ꕼ�xd_���n�;	���uQ	L�Qd���^����nu��W.�*7�w���S��Z��Nw�qA�e��q����R�d�w�OJ�;�Q� � �{��ii�
2!�Z�%�az!X��KH���a�~l��+T�׻�_��G`�#�4�"H'1��S�;Q_):Si�u��V��c�NY:g��\̫��ܰt�k���ݔ#0��@7�o]�ى�s��b���U�Wy^�|��mN�����;��o���Wk<���@w��/(ߛO"�W[���,��$��񱉣��	@}�-H���O��u}Z�"0�+[��v��m���1}�Z_ҁ���w(:ƈ�4�G��eGx�.1X�p�a��c96՞��[���Q�U��׬\Xu��H��>����J�P������gҠǘ� 6x�Q�j���=Kpz�����@�bY��'@���++�N�`��b}T�� �_S])�<��7���$@�d��޸g��}���q�I��JQ@���_�hm�f8 ����)������p��8����*G}l*^o��g[���0���\�6����j�A~�S�DmFQ#W��P���r{s0��%�������h�ԶiXD�-ۘ��ٟ� �� ���'&E]2I?���Z�fF�T%Gٹ�{�[��r�r�%��Bn�#�u�[�A���Eg�۴�Y�{�4l��X�]��~Զ�W<��bj���V��˯��!����<�\�['}S2�q��d�� 	�����DW7n��p1ֳ��80lCC�>����	��Y��X�/"V ĿuV��_Ⱦ6C��Y�4�}މK��՛���I����̡�ܠ�xL^g*�x��叔!�WRNۿ�h��By�T[�s�B:�t �������?���5^Y�)�c>��fi{X'��ҋ�=m�DӖ��;GưT���3�0UW���q���h���:�}�tr���L:@&�S��� 4@g(]�E��'��r���.�)ծ}�sJ+}: GPVnQ�v�$���I������!�ޝ���qȝ����r��ގ����µ�Zm|�a��9��f#k��5���rW�lu�<^w��h�j�U6&��2�%�<�����椖�>��8�Z�7�N6��6zX��_����$�'W�9����!h�9=�0_���|ܰdh�ȫ��Zk��죬��d^�\�|�m�`�O�Z\����<��v9?Lr;��_��E]�M��U���}�;U�>�Lpn2$��~Vnh�`b������/�2��� =W��!粦f/��$�����u石|nwVƛ�=C&L��^��₅�x�-4���뿄gz�u��m���v^�Z�4��)+�����Uv�}v�l���֣��T�9��&R-]$'m{�0��mW�Y&0��QB5Y���C�^Ub�.���d&�Vg�tE&!Ӊ�L1�
ۣn��H����N�[�D��>){��+Ob|Kv�Vu_{<����S�a��M�������Ґ��qe��OV�u@�<���2�r6e�x;p��˳s>�h����8|�f��Y3�r1*Mr?k]�dZ0b��@,�^*[����[�(!�^��>N����:fH�H�����$��iK�>�"꣥ �g�p���٣3���5K<\la���!2�x��l�4~@Ur�]T6����F�����&(�|/�r;QA9{ 
�:G³��lT�u��%��Z^�S�i���ai��&�2A�~@_��A1gKd��6�[���/�m��>�L]�/�ds�փW�vS�QC[��L)��p��	$�$�P|nH��4�H+AGX᳒Z������L�S�����褣�>���N�ቼ���n��L�W�O(��Lu@��6���䗙bZ�њ������ϥ:~Ya��E����˃.ee2����}����K��2��yJ�m�:	>�_���7�<=z����zz�Đ�K�V�j����ۻ:t�Y���zT������fg�-���:@!]����)A�����k�1E�"˕^e��ύN�Z����g�x����t�h�]t��&r*YcK��`b���m��saIA����8��%X�GDk4���I T����>���J=#��}9�_�/3�Yhx-�Z�WL8t�,?�[\�:�Ջ�m��-W�e5n��z����j���3���堞��[T��r)j�d����Az={]5C7u�»O%KS2!�S�����48�p�c�M�ǳ��
m�hM���eR&ݸ�I3$��!���w&�#�?T05-h�ط�Hg0G�,����E<�^�"�l�}Wx`��J�I�Sɡ$*T`��/��}K0���j�`߮�J�q��?l�I��,y����v���[y�����S����rj!jA:Q�S���Lf&�o	<�c�7�!�y�+����6-�	���oۍ+,=Y��Ҳ����ziU� �Ʌ}A�H'5��~1�^�"� 
{���^=�0�n6ڷ+vs������s�+�g���1��K@�'���l.������8: N����ESQ�[�
�:N&$���e�s9�o��`� ˄��a����P������e�MN��UK�ȩN""`i��(�,��@�Ȫsn�x�Rʄ�{ҿ�5�6��R��:����䀠W���l>��x�B�ۛ�Eݦ�=p�5~�&j(��o?���B�962��Hq��ۊ�G�K�7\�o�����W����L2Br$牟nnf�Tڣ0��g�y��I�f�!���S>��4��I�-RC|�S�u6nMz"~+�;�B�mh�oS����5�b~�i�Wr�Q��l�D>ǈ"Q`A'�.e�%y˻C�G��#��hݳ�_ah}���O�5e�C�ZG?�����/��.��+�IYv�Cv�L�~�4�n��hO��*x��������,TƘv���8�9���@�8���\�<��,;��HYsF'�-��8��aVT}rIu[+6Dy�~Z�]�[���a��h43�Q�v�-@!Ҽ6&>l_���b�@�˱�QT����]���5��2���1]�̡�fZ��d�3G1c�IE7PIt�ы���*0���N����"�,u���5��K��c��^t�U�@�Fֱ��y1?�R3W*�����ƤFg\��Sbki�+����K3����I�a�V�����kcr')7^^^�y�9�Ob��E��Lg�}N�8�t"1�ձϬ8�7�=��+�~��u_����n��"i�-�[��롩'�2��VCU��)�H��x��<M�ը�D�.��p>=����/�&��v��>�E�d&���Ug�38U�*��!�Yw����nrlV:�e�&��M�N�����M�]9.�Q�Z�& Zeq�����I��n�Ȳ��Ɗr��pb|����5����2~_Èف����	py��+���ݞ.��~�X볃X��6Ƀߞ��,m�o/�(M6w˸'���Q��N��µ�T��(�&Ɠ�"�)�,s4���\ҷ)u�0ik�L��Z�}�?'f~&h�=��u?ҴS
��~
��a������[���py�U���Cqz�$�<htK�p�}��@<UX� �,\;cj���*x��GL�����'�r�DM�=~���{�:z��,08�����[�� �{!�o|�H����ZK$G�%��x7T��}�C[��äo���R��iP��Jd��Mю6{�9�ZO�~@�X��|�[W�i��=^\U|��&����o	�p(b��۱%f����.H��M��Uk�5�}�ZG����+��IdVN�CeL���h�<�`�*>0~����T�rSbO�"�ҩ�k�M��Ob��jk���&��ɑф�usO����1PJ'	2�:�D4��[�S'�6���ŝF�=V�=��:N������o����y�n�b��qߗӽ�������Z��:��F��/{N�M�ɗ35k�$QyZ7��Y�<��n��p��44:���:��{+�W��<�#�z(�e��`�|U_�o�e�����X&1�<�p��.��/���{c#��E�~u��;\:e���D���b�(;6����eA��\��[c��UoR�F�<]İ[A�3�|^~�4�z����(8�Z½�q�\�l!�����}����۔��ZU{(����왻�J*���|�)�o���m��#1;,��X��~���j�C��	��^j������}�w)�T�Ͼ+�����ڛ$�϶ě�a�G�_��&��u��.��� 4-U�8zU����#�'�9��b�Nz>]x����{���;�)��Vy�tߝǾ���8RW��6&�գt����Q/�԰�U�<�ZV��%j�����>�s�������D}��zie���[�T�n�
����y���2��)�����\`�.�w��J��+5���=�Z��tǽ�u�NQ]�����S��e?�p����)c��ř�[����.�� Ӎ����E��_�18Fs�y�R�,�� KצU-3ӣ0�UD3��L��Yʺ�즬�3�9m����u_�Dl�ˌ-�,��W�P��/�&l<j�7�*�C���Ḩ��Խ{�Lw��S:(��ט*{+ ��O�?7+F�t�t��ƺ�F�7[�n�B�m���<�����3�%����訨A���嶍��1�v#U�Z8���	C�2d��Pj�ͳJ���I��3?��M�7�dD�p��/)���������O���w�j��Օ�����7�*ta��A����Fle��k2E�p��R%�PpOR!�V���*m��n;u�Uʸر�xs�͛�_�U9C~v"���O�T�$J�҇ݏ�?��6�4J��+[�#,mK��U���ޚR�~Fqe�k�������|��q�c���:�0&�qk�uA�Ã���#��2Zw��&牻�E�z�H�1aldj Kʲs�~⏣�~�}O�M�W>�s�j����g�wa�Qf"�7��ԆY����^���D?T�Rm�;�qX�W0�6	��%���ݹz����y�:���a��������$.��%���*��ȟ�j{�:OV-M���e
���7q�'N��Wͅ�ll�n�Te��9IE�*�a}k,�\�N[7f�E�fy�xO�類��=@�-N��L)���fJ#�S@�Ӯ�ZW���p��uٹg��m�k 6����;���>)�������ʔ�[��lXWTp�,#�xm�L��)�:\�.Kl����f8 7Oْ,��4D,o��?��u{��{y�Ξ��]џ�����2j�5�o�N�����*rm�XRo�ŝ}�]�Q�}��5�`2���~*�߾V���ѝh
��� ��T��
��6�!c�,��g�;�f�s#���n�j��{ޘIkv9�8�3�ōo��˱�T-�:
��2����A_�K=͋����!���;M�V�;qW ��ߪ����DH�U*���#V�ٰ�E�=BA�pc��Y������p��u����MiM�++3��m�m�����'	%.�4Uf�>�Ņ6����R��%zP�|�^# ��DW���S
w?p����h�E:��P�b��稾t��1>ŧ���݌`޽���3��LE�/v-[�����J�$_��Y��X����}�1М^�9C�M4g�]hJgTՙ�x�xb���gUs�Z�nS�K�e��/������1fJ��X�Z;U�r�?�hP[t��½�>]�����#`n;�s����N��c��~����!-�ISwף)oܢ븖��J�O�CS��/f�JF��jd��N*��?�VN���"ꃫl����3��O,#3�Z���/8����>���g�(�=�����ӌ�ޢ!9Y%Uj4���-q���n��=q����[=��rPA��C�6ϫ��X���f��1n2��1��K	z���Gڧ��"I��8|����*5?�r���j�-�9�oN�m�Nzk ���>ə3�N/["��m�n{��Y����kB���з���M�4��u-���v���w������X�-��^��gU9r2m��J��I��u�F˹o�_��fkG:֘hw�?��}_'xkk�=�Z敆�㝻��v�^�6��������/���٥�L����m�Ԉ-��w�e%wߢPߕY,S��s9Yg0O�F��z��Ú��]���d�:j�AK'3�)i<��I�>��is�[�>���JU����:���	-bJJÏ���2V�4�$W�1��J�gCݓ�;��S�#!��@춸s��Uݖ���]��J>�&�s�P	��u)�
��޴z䅂���/9E_��HH��������_eV�:x�U���c��,`�}{�2�zpq�Fs���94P\���ל�6�+�m7�p�b~����HG7R�3�^��B���4�b�B$�by�?rAc[چH����\ק��'��^oV9��7j"���¯(���[�#�{�=�c.S���2y�_������ݕq
�oH�a�z�
�����I��x������:�~��~<�R0��:�
�e���ܶ�8�m�و��Z�xL�3�_��W�i��N�Jޅ��xP`��Ʈ�ɥ?�FGm��Q�߸�l�
��Z~z�ހ|�R�)˓��k')���#��Ȕ�,a4A��.�-�y=7�3�=B�%�5�(C;S��P���/�c�'J����gݷ��+���BO��G<49i �O�Tb�����6ƙy�_�'S�����ɧm��a͖�нE@�Jc�I�v@>
�ngZ>3�+�e=����Ѵ���+�DR�>E�xDN.�K��`y^�x���
�n�D\�t,����2��^D++}��NO�����+锋B";�Q���~v���&�櫫��=Z����g,Weo��CshC�o�y���M�R��om#�eO�B���w�V�ٗڱ�+�x�������H_�|��%´< � lW����#��O+d8⬘:����a��ct�O�	�e:��fñ����3����A?E���b��)����P��m[G��J��v83�$�^i��C\b簚,�T�Ы����v��ViP�mF�����vw�t~N�K�h'�m] 6l��!��
���g������#�� ?S���/��� �N��t2��L]���LŴ�m%��&�P�|��ڷ[��6�9��:)�Hp:IH����R����?�������k�7�!�a��Ώ�@��cH�.�^�H:��G�W@U�}_�	�@Z�)��$$	A�C:E	)�CB��n�HJ# �%!q���o�{��c|w�7��}�^{���k��}G�R
E�G����k���Ն{�i��	�r��޼H����3V�Z�n��y�V�q�>���6�����ZH�bhA��y�{��m��ٍ��N�hl�7�A�)�h$���
X���Z�%�6���� ��m�s����怦�n�2�ÕZ��-2�$�����?S\��V��J |C�L�7��%�:|�*�oU�	�B��&ҽ]��HS<������2���@������3��Xj[�#t���f���z៬�GL�{Z�WsG���n���� ��ʯo�F�p��
8���]8�oY�������v�R[�S+q�pR��>f7f3��[��ʷ@-Y��o{�{�����0�Z��
���cqgQ��(y#H��b)�g8��x�t�@�t�d�=�cf	�?��.i���Pc��4��2��u��?߮�D۞�j�S<|�O8�`{q��9#�����
ZU�-ֹ%�8�D0��HN7�|"A���(g�K���@�%�vZ��h���'
��>	'�p�V�*N�jv��w�A���ݱ��}?�F�i�U����ѷ�D��1�&O����϶�5��ΆtDo�IB�/�4%�k����w�[��䌊�nlÃ-N>��I��F&V�I�o٥�S�n�1H��\YϺ�4>�����̝��q�:�uLN5��'�1q����/���U2���
�g$�Bn���L�6L�-L����`��ڽ�	��p�M��G��=��ñ�!��	>�w��G���*����RE�
������W]�a-�x��wXr��b���-ajp/
L��(��m(h��W�&b0[�ľ�6x�3��:SS6�����?�ꆖE��;����#7$�\TJ�+���ig��,��]ߐ�{�9|���qkR}�ȍVN�J!Bg��N!�Y;��x_G��p�9 d,%�-� ��EUt�-�1�1u7���xj�W��!��~�e�)].�\�#>k��B��6��87���П�c������o�:��wy~�:�%=��:��w�L[�?������`�é�����v~�j(�A�J��k=��:������i�9� >toU�����/=g������Ѣ�j8Wg���c����֫i�W���� �^@B�fD&Ji����
�[E��~��~s7��C�!�488��%^� �s���v���Kw��.������@.o���1�Hq��	�9��m��|�����٫�r��;)�@>h�"��I�43Ӳ� nɏ���v����]��\�(v�*��߿���'�7=HFnؼ���}��<��	x 5�������`������Z���9�LΜ �)qn�U�?��}'nL�@�����h3� � �7|Vk}�Zm!"��e��n��m\k"7/R
T:rjc]@�,M�m�K���o��{�Ƿi�U�t�S�~�s��즼t_p�3n��c�?��%��ܴ-� ��/��;]#�$�\$�qT�o"L���W#�1A���'�6Fh"�C��ʹw&�f	C���[��K�KqJ9��3?��q�zB{����G�F���~ޑN���ڛ(����J���7���-��D��}���1�`F ���t��0Z
_��1���>�6;��8������pc�ڸ��
nzq�]��ǩ�6�+?�E���힆�"�/W� h�Ҷs0_��v����.�@�*��?�2H�y���������[�ʌ��#.R~ߪ;�}wL�m���а:�ЏO{-�X�q��R�
�7F���٧s3���ſ�&D�M��v%� N���M��DG����Ȱ_�V��8�#\�:�W i�o�t����QM��to�,!ƭ�0@Dk�|��ƿ�aSl2s�A�����<"�w}j��@��ڒ��k�t�&s��J��DB}l�al�괲��<G�oCr!_�0�_Ť��-Xn�� \Ap�t��j��A�#R.��Q%��1�hŪ8��E�$�����j�M��a�}%��:���e�Ϙ�C��Zn&s�mⓔ�Xwǲy��j@|�ݨ''�����R���k>R'͸^PgN���א�Ƚ�'	�&X�LO#�Ú��[��i���s^j��0P��f���U���G�#������o���%���u��42���_}\�J6V��7�M_o�#=�?���~=MM�مk#4(�F�Gq��JI�p<�w����2�[K�;�R��h6(�fNx�`gd�2���,�k٫Z����¼���Jo�v� к�TA#]8��m�#ϛ�չ6�/B��;t���1���;�
H�AGDY&��d���FS2d�;����p�
��T��1#�;��̫�~n�+�\�<y*����j�=v>u+��/��U(�!�,1}�ýl�W�v�"0�\>����g>�����C
_�!7KM3A>�0[����0{)���`���p�Xz�!
��,�V/��KMg�#=[��)�J�t�'��Em�Iq0���Ý�:'�����qQ@Y��YaQM����m��^a`�5>�C�Uq9�2e�x�':a¬�̄�S�h��v6�U���]�
����\���4Hs,��B��V|��U17��G_f
_1�~��e�.�-������1�i���g�iQ�G|�?VD<��'1K?�y�!}>4�����9'pL���H��&���R�:�Ua�y�_�(�dM&AnxBt��T�ϡ����$�p�� K�)��?D��ϫx��?�y}�9W��'����/S/.S}����p�ET��;�(t���t�)��q� qA�s���f#��_���V�RN�V8�H�4�{�� N=s�X�֖�i��'����w�di���#٦g����ʳ&�l����ˡj^?Gi�$�A�a�N�g|�ux/��Ÿ�E�!_z���% ����̄�%(c�ǳ7���l'(9Ll�3P_Ɏ�L����͆?%���4tC%�Ø�b�M���I�fkd�����7_�w���W1�e �7�:-|���d���R��'��iD�KB��f�A���ql�_7�T������1�H�ɑt�1��K6���H̛^��W�K����\�?��
H7�[����J@u�-��/�hoQ�|E���:j��#2;�����X�����7�TA/G6Q�R$S�\a���� �u���94�v5��ذ?Ip;_�D��1�+,��")�N^!+�Dw%`��:���sg�@0@��҈߯�D �X1��E��?��C`�X��i�xJPR8����Y\�؛TLS�k$>�/,}L�Ql�F=Й�">�-蹊'�p�K2��^�{ b�V{~y�|��^��+��J-��]��~h�

SE^R�х3y���O�Jƶ��ߥ�2)�}�Yr��9�H��AQĞu۽<�3Q�69��	|��E1f����*I!R�G&�pÛ�eK9L��͢�5ΥY���&(c��-�/��{�;�~y��uἹ{�����O���������r(Z��kgϩ�<��\M���U������G_�x�W�g]�/��~��Q���d7���Sg/KWvb��v��?+�F,�G�n�Ir.���{c	��<Ț�
q�޽o-����`�!�#XE�|�TH~���ջ0�7U���;�"��s*�����=��zRVot�T2�&:;h�B�X�����֋�`]�4i�5�4��v�Og�BX��tX�r�d"o�
%/�p�P�Y�Q�WLʋߍ�<'�.��4�r\F�T�YfJ#�o�ƞ�����V��)N��^).�}P}kCW�S�ۭ� ���ø��~Rd�<�|��<-�ӫ������e?#ۻ�z%\�t�5��Q�^�������4����#�&��qK�3_s��{{��B���%j�����ѭ/��yV�I>����2J�bI�?����f���	m,�%���Ν4���?�,�}k���v����+O���A{�_�y|���R��m�=Z�mn���5ۢKa��-j��+�S�@�����6�xj��ZT�y�^2��̈́�e����#���u��i�0����]�q��svm���kJQ|&{Go�U���.xo�eڽ^K�jb�|k �aX-���_*O�>���w�i$�!�������F�v]c(�7r�j����@l�a*�讟?m������-  W૵J�t.>�yw���]�~�"�ȕ�W3���)mKZ���UAz�ߟ�j*�E	�ˢ#׆����lP��ķؗ�뾖,�?��*�3\�bi�Ԥ�!�__��F����"�"�2��M�rB:>,�p���XS��>ڱ
:ވ�U$����:%r�ʲ��kf(����,]~
P������T�B,�N5>�4w�y�2�3U���j��K���n�i���!ыX�*�ݏ����"�8�R�����+i��v
X��>�-�M���AF�sm�����n���>�(WYr�:���H�KqJ�Y��WL�B�\�u4mL�j��W�^�W���t4�I��9W*B�M��h[P�J����@@f�*vNyJ��h��;�#_N���fi�i��q:W��bE�����)�Y���A͏���=P�2�����DMN��1e��ɥ��O�K����/���=Cs���A�#�Dk+�������v����~y��{� ���}w����������}���B�4�i0��e��M]����E��^�y{�7��kz#��˜�/���w{x����dE��VX����q\���J��=�]�E���G�\�$.��� ������������|3+%W�U.`0Ҥ{w��*\��=,R7>b��+�
�����3��k=^�Bu�#�݈:Jut4O#�����mi,.۾��z%f���W�^�Bp{�
±��X�������^o/)��ɖ��Q����Z���T�����.ե�?`ZP�B~����Oݩ�99���Ͷ?��ֻ)T�Dؽx�P�U2$a漨�Ǽ��b�͋û����.xû7���0���������VC��7�Z/�婅��[з9�/K�ݽ}��<u�� �}��.1��	�9�Ѓ��][�&�ٰN������������ו���<���׽2�4��6!����8��6�3�h'���+A�����2!��>ՠt:>5~Ԣ���;��_�u�(�~\~}#8���o�lA�{��K���gh�m�x�/faں���������mN>쓍4�ĘW8_��p�'�O����s����a I���d����z(7m���S�U@��ޣ[��
�$��:B����Y�����e��%���_!��.�LR�@�G��^�PF&�m�!L��jb�����5P_X�'Q� �K�n���΁ �Fs�?EL���v+���F[l��߈ �5��]�Bg���;�\�O�^O0D�R~á>��+�\qjO�9b���D��ۈj4�N������.�a�'�'�!mx��5��o�!�#1̕u����d���~� )p��:#��<af�,t���4�7�p����*J��@#Dd`���L���h�<�;y������
mx�
-t����ᓻP�.��×J��ڝ�5�8��	�7�_[�/�����nrѧ��'�4�% �6�6���[55�s��㗄����C�Z��|�*7y�����|j'� 4���@���۠q���un���bd��o^^��~��	�9�Z��`���S66N�-���4Hb�3�^����i�ysV||��vF�D����S�Fk {�\������^��i0���w���y�5���:�l���т��j�vP?�|>�
1��RRV>+nr���,��4 �&/��%ke`p������i~1&%ZE�Z�#����ȸ��A������7Y�=:_�?��>k��A��
5N���&N��w)֟���Rڎ��k���y?�z��Eu�%��5���/�ɭ}[8M���m\�V��)�g�ٕ(N��6��PZ����kgo��ZM4��mSA�|:��������U�D������χ˜붯u[�p=T\�����2>&BP�O5��v�����hl8�Їϗ�����f9��de�HI"���[�����*�B�w�n��Rn�;���˷�~�AP�,ec��;wNP,A0V�.�s;�|��\�:UM=z ؐsެ��r0]Lv��W��9��=fp �o�1�ˍ\ɭ�~%4�b�E�CBE�p���:⏒�n{Vz��w�!|
��^��	�~�U^|D9�<��k�c�*\t��q��f�W��٬�UX���1�)=t�RK��e�go̓,���q���ӈfC6�(���Ysݑd����yӚG�>Ix�|'!��^�|�?Y!ގ�ll����	O�u�W>_��dv�D)�W��
;�$Hs�����1O�%�(��Q�n�f��7<�75k�U��Y}=��s�>�H�F�'Ҭ���b��������9�6�e���<��}�f5�����z��Ÿ��[H��Y���85x]��?`5Ŏ +v�S8�e��\B)��3'�(X�]ܢ�hϼ@mU\��K��Y��d����*V^�#-����~fu��<$��������6���oL�^��̡D�u[��݀Q���H�Zk��ڑqů��!�A�"�p٬���B$X������N�#=
"/�	�j��f8��z"V�)1�<�?�9P�
pЅ�G�̄>�1�����7��@WQ�hB7�_(<�&ݟ�۸���ͦ'�>�����]N�� �����v<t���3�I��/��bp���ڸ�zd����q�C{(-�^@��r��r��!v��#��}��o��v�b���/aF�]L BR�$��)��X@�p��������AG�@ੱ��ߨ�=
�qմ��-���}����_����4�l���%0=��-�	���>y7��ʿ@���=�8ΰ�j�dJF27iq#L�8氻ؘݳ[)q2��O�L	<���G�,�M?=��-�ky|��lM�H�H�3�	���%:cX�r�2N[A4�����>���S�y���'-Î�����t9gK�ǨI�
��~A�_�*��`�0�P.���E�T���2fg���X?�a�Px;U�Z�����>��^B	�E���|���l19ě������C�,�[�לAz(B���`+�9uZ;����f��S`����B*h޾Y�02iI
��\= \d(�9mV�)g� ��S�=���\>D"C7�H�U3#��q���$6D>fp��sTV ���4eV�?��"�ر$���ŉ�	I1@�H������e�}A��w������^`�,Oo�n����4)j��}��S��Mcc�q9i�y��a3�&&���V�N!]>d�m!C'����p}�f[�~F�O����?�e�}����`vd��H]"06�2/-Y~�
玾����hv"520�2(o�Q52�Z0sB���1�S�_��A�(#�/�w~��o���?��j�D�8He&�h˛.8������a��m����#�BHX��D�# A���>ǀ�{�������ȠUP�ua�]#0����S�D|���RlJ��s�az��)I�ߌջs۬�U��G�mt��/�w��2>�P�������'��T��I'H�����=��_����Z�o�Ǌ��k����A:)�	m(j�����ł߼2�uB`�}�瑅͆�L�Ѫ���R����3`!-d{�9�'��n�\V�4����EO<�T�Q��$H���� /(\%DĬ�Oa�`D�RY��T�(ʝ�j���&��WX ���Y�K�J.ê�i9���]�{@��B�Ӿ�� �(	�  ��4�p��x���+ß/nsU��"D��67��.1�j!0@u�Y�#�{rm �"S�!����� �a%���@���."�E��D�� Q{����'|��em��@�����	������e٠7�	�J�j��Y�ŷR\K�zQ]��X�}����"��A�S�nu�%�缐֭������R֦@�kيc㽩x�� Ah�lS���h�6��c���;��,Ȼ�	|�ע|ܤT!�/Q��1��y$e�!	fB[pM��}
,@��5� ���&��{�8��5��W$X�㗉�b|ܜ����+/�q�Y����3L�Fa�������Նed.�j1ό��p�|�Q�_��kZ`��O����zH��6/�+9���~��,5ۂ�<GCW(a\�����#�xz����6P"*5���b��λ��ȟ�_W���yqR$�T�Npi��[VV��w��N!cjxG�dXP�'�����<~&̚{����_�.PA�<���J����G_��7�eVo1�?L̰�g��,���oW%�<{�|����b�*޿w^1�l�������l�2�h�Z2��US����!:q��L�G3�pW�sz��u����A��Q����L���e��8��5%EQ^a\�}n�5��O_G#e�B�l��S�UH�9��>��y�@�:��Ϙ@?B�tHho�3��e0�ѮK� �Q��#��n��(�)T�4׼1�Q��5֘M,��o� ����I{��s�L`�{^z�#���%�Fc�� Ra�wo���(s���E��y<�!���	�늟�P��ҧR�c�ģ�W�O����~�AZ=.*~��w�ga��X�(F)/A���b�fY̛Y�Ӧ��pؘ������0�f�y�h��i5Jiz.j�R#���E)��a��7L��D�����Y鄲s)q�{#+��"
�c��a|��#@��+���e2��
�N��Y�ck��f�J%���
�L&vX?Pl������gr,=�f������ȣu`�l�z��V욹��О�#�oj控��Ox�2$Q7� �+ �] K7G ���.$������yKht�z��<>�U����\'�8������<�I�HP�`�1�<�X�
������xl��ag(�!�wH���ڦ�\X�����b�x��Y ��UD���F[Gj���c�k/ �ڒ@7�Lf�,1HX�kw��>F���i�7�W�k��@u
�g����o9ߑ%/wzR��M?%q�_J5o�j��_�ѐ_⥏�'�EZ��I� ��if-�t�s�E�B�l�������.�?����7�}qW�yy߿@`�;��U���{}8Rjp�X��z'eA�f����~�N�S!)$}}�O�+B:w~��wB���{����,�=[�V��:�T"�7�pYKC# @~��<����1�Œ�'�	C1�wA��ˠ��.*x�d��/��$w�@b��Ak�`�ȉV�$UET�ܳ�
b2 ��ac����>"�4��ro��D�Ħ=�{Cr��#��4�il�	�pl���F�1V1���*�=��?m=������=dز��e�	���^����:�\��N���������<�UI��)�HQ��^�����!�=��N;)��k��鵏���0PKzx$a]'��-!-ȵy�˺�-V������c��}�vL"�8���	�'���������6��v�O�6ҡ���o��K�I%�kf�n�w����L��f3��tL?�H�&#�~ ľ�S�2�6�J7m �i�Q��)�㝰Tϙ�eB�2�b���ů�)ύ�^wtX!+�jm3&<����fw���6-h,l.�͋�N7^(�����p���?��u=v�[�rV�U���D��n7�CO������d�7����t�qs��>�{� ,P�hc������%��q4�������"���X���T��O!l*��[;?��V|���.~��:�o�s��c.ĔY�I��~L����I��	`�R\�!ɍ<�t��!#��0Ւ����!MCC1&��v4��#
W�8ʓ1���0���c�}	<�X6���#6������բ ɂ�o�䢥�NO�S�ɫÑ2qf:�����ސ|�H$�'�c��g�S��ne�5������I�͸t��D��xh���Z��d��O���o(�A����Ź�ދ�����hv��N�%�jxR�7��(sHRM�����:����������O2DZ2�&���A[�JXHϹ�o���^ǚ�d��E��Y�c���炾�I,�� �?)���[�f�8�3�:B�+(`�U$`��RR�vYtf�E
c��.�J�n���Q�,�C���:D"��e�ViF�/Q��V���yFi�5��]8r1�|�9IM���A'���@��45|h�P(<�fϹw�OE��5��Otn���Ue��b���2�ho_��\���k&E'���W�Ĕ�~��efj!k*���馯�D�:<�p###�[|���|���k�E� U�&�(ʷG��pa�j&S�0�=<��k6DP�lZ
AEEG���O.@)�����)�<lrbAPrlă��o@� �2��}�"�M�{��Zd�-IG)�G*���w5A�'P����[�{��,�t�rR�E�?%W �"�����������}8v�B͙ 3=1�˗�Ђ��	G�%�`UbV�o�ҵ�BW��@��ۚ\�џ×iT�tf�B[fM+՘Zx�0E�glZ@<<T����.č4HO�K ��9X�@T\ �[Gh�%��FT�r��Y���E��g�s2᥽�%9�4ݣ��2�Bb���O��`/��'t���Ƚ�x�)�w�S=o��Ӿվ%�y0�U�0���pp�C�>�3C���_��T<y���#���h e�F
��3!z�� YY���hx0%��*z��{|Wd�T�!��kg���#��d)�Y�w�|�l���DY���;uOf��N4�uA!��I�d���g�ZK��ڰu�0Lc�S#D.�!��~>0��M2}I4|b�ɒf���9^A��d��ǈ�"{�`��T�[��E�^�L]&֋����S�?��I�")�P-ӵ�и�|�����222�3c�Yv�V�
2������R����1���X�a����bϰ�zB�~�FL`�'���K�Xm�Y��B���8��-�͛?�8m_#����3%=4�E��T�]�N��_���V�m��߼B��xv����{����{Ńa{��xNެrWT;6� �r�S�����U����>eCAtU~�ST(+Pߗ|�W��k&[��ů�3��\��#Ԇ�8zWQ\� R�����z�>@@Lҧ �+�{e�=q'��yB�#6�.�;��FG��fS�+��)#���wn�K�}�x2C :{��lZInY!2\�e��[�R*��� %��,$F�+9nV��c�p���<���9����Peљ��v{!�9��W�nd���6���O|����� Cܮ) 6�[vI�#L#��0`el�L@i��y�UڸЧ.��7�H��]�u�[�����-�l��L~ ��mT�$MQޝ���=�֙��Գv`�Q&s��a�M$^��}¤��e�q�k�=��%�p��/2��$Kp�
�$]��cU�8��G�[吽` ���BAI�'$�rLe�wnpL⧊,�>�Q����+�pGB9j M��K?ӄ�ή0B�s/~�1������s��[��!�BC�@�{�����R�*�w��)��B�t�"G{/���B�M�>/���Y�u��7���L�����K9�:���({(�|���Si�GeF+��K �bb<����X��ө� �#pSX�G�&?�5MJy2`���l+�< ܢ)��������Y�P�0c�U^j����	q��XC��J�ps�������=���s��@�숍����	Z�6�w��ت�����O$�#����ʔ�7����(�5 wܸ�b�!�b�q���D�
��L����N]:W�hA�phpx:E���6��J�uС��0�6�KpT��0�'Ć�1�����i�!�ϔ���>���RNp6uĕ�jj"�X	ǏW����#Ӎ��	�~���۠!�3�$��._&�8g��jK�o���2��'�"���ζ?+\�QJ���8jx�h��S��+4�d<��<lg-��WB^~�d�;*� VbǄ�)V:H}ZQ�b�~^��Gʌ3z��7�ܧ�r�bel{ftl7E�dDثpՂ|������ARj�S������ue��0��n6�[�H�K-3f�ƫ�O��.Hs��W�7��$�4Lk�tetkb�y`�"�/GF�L"�棂�u���A��+�nO�������a�HN�zݑDdQ��"��V)�?��h�Z�K�s�H�B��#)��W�g^�`��U����'+Zf�ᔓ�k��o�f+��Y)��0�p46q���Ϡ��z{/�6�֮r�Y������[�]
8���x�k�[Y��IrPt�-{�b���ǖ�#��κ4X'@
����ɮ�Ƞ�Pq��*t�2)�"�'�eļ�@t8]d���r�u [����쬉���^v���	��1�N���^P7f;*���j��Da;�=�=��0�G�A��+�g�i�$�'���#�[hj�-g�@�`:g�z����˜��U�Jy����\�nN�ѷ���U�����iJ�?e�*C�~��N��Q�P}�_�����@��V�SK<��]��S�Nh�����Z�I��z����P�HB�'��nw��|w������}��o1��ē����D8��b��W���dU�����~�LW��-;���T8�`�6(��LK�+����*����'L�:q�%�x���\����uS�M�!�m����v�P��a��Rh�X�8�殽!�C��ݎ���)ey1��	�����r��D���n�MFn�wsl�V.�<wՒ��Bw7�Dl�b9��i���`K7H���X���;��!���ȍ�P��6��"..O�H�v�MI���q�>�,? �Q������@���z:ޣ���O�����"ƾ+pJ����⧷(�a+�3+#��=���?��Z�M<���f2���x�|�UN-��߹�/���'r���%w�ً��:�^;u ��Q1�,l{0O��R�1�6��\Ծ[���{;�cބJ����)t"l!-�l�Io�pް�z�XrUL�*��4i�_�����=��5�q��Z2�)�1R���m^�j��D�p� �f�zr5�p���*�>����k'.��:�Mp�q���NA��h0��bļ��-Vݸ!^7k��_K^,� gU?�u��.(�b	�W&�:��ǻ������{"�U���}��3#�-�*�5Ի�����J]h���[�`������YWs�wW]],�Z��7���\����x{�qb���΢�!v7��r�lb����QnO(��˥(��dR�����!�?eZ�>y�6ddmr�rQ�*�t�J�ŭA�#��.YgF~�.;h�?���%�R���d.�L&��( �9��I?йQDO�}~P�z�#׮$�
�ȩw�:��+2ɚ��!m{�.��Ԋ���p�SBݍ�e�����sn�|�p:B�O�Ͻ \�
D:�|f��|�ee�C(�<&�2��{)��q��/����x��(���%Ѿ1�kX�ٳ��a]���p~vO�I�zT�݇��{U��u2��L^ �޼����kl��t$��N�M�%�?�+�"M5q�s6�8�������vB�$]��9�@SW�(��3N�^q�{��/_N��oX3���~��Ǭa.�786(�)㗗�ݎP���jH;b�;�����D'{`@@={��^(V�U?�q���sit��p���[����i���h���$��f僗��^m�T�a�G-+$\##vÎm���S�%�2��]�m��9&�����hp\DC8�Ћ�B ����>�=���<�����݃PJc��_�В��:����YKn����3�;_ҼI��?�_�N���v��HV/%M]m�6���OO��/�:�	0�*�k�z�Mű�{s�;,��$i�5Z�6+;�wi����:7�_h�E'����,���K`�9
]�
���.`=��v_�(���ls�_���ȴ}+�=PR�ʈUzjm��4��� �#ױ�Y���O��F��DJ�\�Me�#u�\��t����2�4u�	Y���(#�(�v���_���	_�$wb|����}��Ğ�����7c7m"�\l4r'��2��\�q��wysr2XC�Ws��DAJM^n_~�����x��<gy�%�7��pki���& ��K�'F;���Pv�ʰ�����h��Ù���	
�������;�oI�GtDW���@3�����)uwt��[@�ϩ�5^��L����}<���(7�T
�K%Y�d��r?�[�y&Hߢ���9t[(�
�%�ޙ7yF~�m"��=�yRi#����2򧥟���}L��t���Z,ȝ��~a�,�q@�=N}�����I˄�_6=V��b��t�=�{���0�;�a��佯]ع(>+/e��M_$b��N���*rm8��乪#^���q�愻�#�hO�9tX�l��m��I��p���F�a��f�ůL�o /Q'��������v�bV�Wa_�o�}�Ӷ�w�/N��$���g޵���a�����Z��M�XȘ!*1��ܐ�?~\�C�g'<\W/��aؙ ��vmIj��es�#�G��J45�Ii\��IQ��|9��d��I����:JyZ~�y���������7į��Y:�2O���o�[�9��6X����r�����X������"zlI6d����^q(��u� e�<���فrk�.Z�����p�y3qU�Fܦ;	w�O����>7��*�L�qM��p4�0�}I+?(@{��x�����z�(���$蟺o*%G��p/�㗼�al��/��=�����R������\����kA�0Y�B�zj/��o���G�ՌU��_P���7|�͵OU��B�s˞�q�vZ��M���R1He��tw؞�WI�S<�K��~eXÓc�H۳�?�C̤J3��a-�B }�N�#�uHx�$�9s��8�;�����[��K9�Stf�]���_T��t��,��eee��o�m[a8�-��I"!�w�>/���'s�i˗�I��E���e1̠?٘�i�r��XS����6\*�	�Q|��9Diu�W������~��fH��[a&�³��Ze�s{	�����G9�����iG{�q���J�p�v<���P�rW,���}:)cU�R���x�b_r��'�I}����6�bJ[OG��Ϋ�ޞ�J^����U���<�"� ��H_�]�<)�v۫��"�e �A��1KО����\�Ia��;�ܡ`�ڏ���P�����'
+�7鮗y-e��#zz\��Sm��Ġ�DUkQ��g��
�g��ٮ8��궆"�.eNO�D�T�;Y���,���C�TǪw�oGn;!ٕ�#'�Flg��8�Vji�%B5�#�9�4���t+��{�,V�u�{]��M#ps���ɳ;t{�r�!�g��V��IȌ@�)ʋ��Bd��qz��o��'ѐ��0b�{�� ���4ґ ;�ٻ u��9i�����K��m��O���H�z2R'^�Ywr��=�j������Z� ��#`�t�Z��ҝj���d�3 I�. B�ַ:�/̕�g����Cwx�xJg§����t2�Ԝ�"\`޽<�4�#>�v\�4�d���E|Bk`����ߴ�s�<טIo3���ಐ�(��kF�0��������ny�N~���B�t��,ݩkA������VW��!1��M[�muP�U@r�Z�����>m|��i�5�Y0�k�C��}
��|론��|9��Ӧ%�;3<,���h��`����Փ�S'w��������Y�yA����0�PUᚐ��2�i��U���Ѐ���_�
 8mN^��K�5
�,�����ۡ(���6�n���X+��0OR�pl�M�IZ���U'k#|	_:����U���-O	g��)���q���x=F�{HDu�b�O�����d#�.����,��Q��,4�
�Q'J�4���kɞ~�X�b�\��_���n-��
E'l1��[�w�OM�¹M��,��ܟJ�s�Gť�*�~�?��Ϣڪ1˼p��|�����`l/��9ރ^�� v͔:@w����n+�)�,\��q%���hW�e�m.���݌��1�wOW�.�eg�(��
�]}��b������NLH������E^N�x��7C1�"��Z�\\n�RL zw�8�;[y�!�p����"���S��x�V�7�ca�� +�I��W3��\M�>���^!�E�ȣ�gy�`��>�tE3�Q��@1���l�C
�gq���͒��Nf`���^j3��/�C8J��Ռ�g��.e ���`?�y
Y��_I{���d��Ί���<a_��؝0h�-�Q>`��)��Ӈ�3�d/C��*�^ԍ.�U5W�5z�K��</�W��!�ڮ���L1h��_0��9!��GdM�U�k�n��d@���ǿ>��pQ�C�)/�f(��M<[3��h�2�][��?�V�˷'ޯe��U@���I�Ī���������)� �zo�&M�G���_}LMD8��߷� ��v;O�������_z,�&�� �₊*���:�c��e �q�He�El��3*כ��3na��k��%��GRvH�l�����5����ci� �� ͚�\ �0w�uƧ}���D�繁�rd�x���o�uf�1���ܽ�J���Ȧx��B�1zx^R��t�"fne�H�Ӧ�`Kމ޽�m7���0_����j<�R����|Ȧ�����|���7��]���T{ݏ��qB{cB'�����$�>�n�c7�@�[�8�b�}t�� f�;�K�{��)��ս�Le�n�p,���k/�������x<�+�`h�@h�W��Q-</���@�׃�.��ܖ�ڪ���'�8�d�(ｖM��칛��_i� �9��0Cӽhip�k|��4����`��ޠ얫J����ѐ���b�Ɍ��G�W��Cr���=�t@��5~�w��d�c�ZWW77�����t��-���N#���W�l����h4ٳ7㺥#����E���r�#]L74̴��e15��jqIT���zW�̗,�<}��@�@��{�F�v]]��p�p�Þi���	U{�>5:jF��Bd����L7�]yש8�x~��f��P&v_E=�e��wp$�i�}��ȳ����#�/g�E�r�YJݍ�����ț�&n������}_����H0�h�z�ۂQ��x��c��4��m�BcѢL�����D�U>zMs
�z���
 � �p�RĮ����y��~{��k׫��tqR��x'����y1��wC��'���[~��$���g�����&��B�?�[�TOO ҾV�Z.:���n�����L�SV�淹DA��6]!�x���3�����5%�P�,���z��]�2U�����T�?�i����;���F2���+]Senq�~�����2S�a��̃�n�Y���.��2�.̤�g�������n{]���f��P��*�ǎ�eo�F���Y��A���c�@At����j})�z�m�D-ۡt_�	�x_'�ϳ�$����n���S� ��
yyj.p��ZXVQs6_�o��h�d������z$�G���9PL�@��]Ƴ"r~��d��w'QCv�|����G' (������j.X��?ҾY 	���{�.�h�~��أ/�f��=F�+��Yxy7o���{�A���Xo�� �;�y����MmM�h�#x^<ǣ�
X(ґ*�r,��t�(MB�%x��@��B�RC ��.��"��� j��~���Aa�5�f��yf�w�����/��ɭ���um�2��y��W�Oݫ�˴����Ta�6��I;���Vg�L~AY߇�c���U�3����fՌ���� K�Y@�kgR����Ǭ&H��/��xd�4]�_�_�����>��jnƯ�3:K�6<�F��i^�cYJF�D��Y�����)֡�����K,GC�Q�=L���%9`�f��|�Vi�}�㪱�ε
��kLW�JW7��bj�fK|�u����m>����O�<8Yw��@����^Kq��zgk�lׇV�Ƥ�����ϟ��Oʈ1=ѽ�~�s�k�qB8��6���
(b�f,d2��s�<)�N�eLMYc?��Ĉ��	����s�\�KvO�'�ħB��[^��SY����ʰ��'����xő� ��՚���e ���<�@Pk1E)SBcf�6W{b�>tn}���ʦ��ut�Ts������:P�y*3��E$��td��t=}��:R)qv���8͠�/Ap���#T���
����8?�>���[`z��W�\�Ҹ٤��I/�U<B����x��$-~�
��ީF� .t�J�9	I���W���$$FP)���nkq5�����/D��t=�e���ZXo�H�^xn nČ�+y9���3z��lE�ԥ�͛
[�Sl��2�ޅk��j�W:���SiR�]�e�~^����}� Y����>kT���zcӹ=S[�0�
z*SY��:��U���BC~D2�ڒ���߻I�ۣ+�>2P�|�-f����$V�����U�f]�+�~-('���Y8�hO�l��ڢ�O[����C6��G�a�D����x|��؛��M@;ۑY�
��!o�Pp'�P���i���"$B��[��]�����bV��ab����iUي	�9�*�<Z��O�Gj�qJ��h%5gS��O�<�������U�͒��ǘK]>B��/���f�jQ�3�A��Rl��b��I��E�=[�в�o�R��/ަg��v"�r��U�$W�ߠ��>T)VQ'{W�q< ��L���9�=]k�M�VDn�O
M�-D.�C�(����AT���5|]�Jj��fH�4<�_]�if��w���*�8�_D��ux}E.e�B��ɭ���z�㜠ᠢ�;����b���q
�X��@$��Lz}ε��J�㚯�����n�F����M%^�;�N@L�Z�Z�Rں#ս���\��*C��P��7�Sg/#ϣ)$N����\;K���T2�X,�!�$�#�%�|�|��,Ĕ���&˕:� h?�Ӹ��Y�������Z�?�����O�{u/��6�#%����>��#�>�����B�)�'!��zq
u�C�w2�4���s�7�#?ǟ6�5�������9v�!�
?�&�Z���꧕O�=��I���a�yE��HC�'��k�dq����th���\d�v��j� Z�rw��k�(Q�������2��}�V��n��旮���f�?*����O�����'oj������;�@i��䞝�n%x��"&�g8n�w�k�7=��+}�/�l�|&3��O�����8��i�L؀b�[Lj������bY)��,]��l4�c�qU�F�C�Lv���D"�����������A3�g�+綗����ۙ�L$a���-����QOKJ�R�ɏ����_|L\pc����S%���"Ԃ��\.;б��:{���޲�g�\�����H��`��IΖc�:�RX��fPc��5V��I1��^�g��n͇44�b��������lfIy+@��B��f�p>	O2�g3��'��
!�@�~����-���?�lT@	�)猈�����l��r��"^B#��nMo�84U,
*_y��sH��Q���ŠzQ��}}�E��e��)�1��ǎ�PEܶ�!���S�WNP$B���\�������-���H�����F|	����V9Ϥb����GgLܟ4�y�w�����>8
1���mDR��kBf밣:�Y*�N"N�����j!�䏑�����+C �a�sfh���s�6L0K/m26�~"����"k�}���n��M&���ҙwex�h��Q�BC�ӿ4���:]'Q��]e^�TN�q�h�`���,�4�5�tS��
Ώ�{uxHDD$��/;e�R�]B���9�nfij���sZQX5�x�>a����޾��47"[�T(+�|j �cIo}c<����^P�$��riޝ��B�1�M�|mrb@��V��T B�n��W����M�g_(%�V�1�־\����Rqfw�כo^Γ�������a�����k�D�@�&�:�l�"Kcp^z馒1i�U$�$���@sp\����U9Rz� i^�R��WG�O,?s��Nuos�K�����3�<��49�~6�A�F�rS0�:e�c޷7c�Ѡ��i�|bǯ�%��?rF
\������0_A��:
.깲�N��<n��!Rn������2�E�*G*����
޽���ך}��V*�Nٌ��^l�����G^��L��H�*q�q�d��'���C�b��L���&�f@�E@������SC3�Kol��2{��fi��H_ő�K4!W��z`u���q]i7H�����z�vcS��|!�c��0ϣ]��g���)�Y�(������U�f��g+h��ڴg#4��]r��^9@/�^t�ِ������2�
h��#������"�$��\�����7�!�V����M��ju�a�ɷ|xV��E��ɩ� ll�f�Z��!��@9 !�\���v���$r�Hs���'�X��Q�?���_���������%��3��J�e�0<������KʫO�i:�%[��<�&A-Y��@z�f���+g>�?c���r�\�d���BA����L�����x�I�Ec.�(��fQw�;��b����Wř���6k  =��D��Ń����8���s�n��b͡?l�}W~%�ר3�_��h�H0�S��U���c�,η&�����/\�-���5��!��`r�ɋ8	�BA4����W�X���4�~�7�Ѳ�?')-��'cӋ�Q�����t1E�,j��V �.��~
Qt������� �afj��_�rc���z�q��6��9�	�@y�'��B�ie9���|n�� ���}(��sm�YN�ҥǽ�+���L��o����9d%~&	x���Ͷ ��R�vV���͍�;�M��8r��|�1(;���"�?Rw���PP:f�eP�@�^~&y�aS�����쇇��J��,)N�W>%��\���%^��g�Yd�����%�J�vz�d�S���`�,�i�I8M�'%�������Ner���T�̤]Mẅ���yy_b Y�k������E�j�l@H-(q5�S���UE>ԉ$�S��x_Axy��i^�h�*{���4pw�7)Z����{v0��D+�g7��_ ��4�o���M4�f�|������[Iq�B3�\��J�R��D-�,9����=mJ������{Rn����N�{��E���p�&4O��>mꁒ=�Pd���; ��tR	�Uט8^$��,s�8C.7)���r��I���6��\1��q�oD�F�o��Sz��(r��,r��Iv����f�h��B�*�]~*��+���=_�%H�R>OɜVl~�F��	En�G�"m��y+��'_�Go	�Xz=��jES��hS��%�\@�Oи�{��H�L��R����,1akѾZ�{"�w_�|�샮{�|���__�ʝrU��������|�����4���c���J2c�w2'zz�^x帇�1�$e�'�S���K����-�=��d���d��8���&˅��F�#����)9��\J_�������'��G��4�{�L�!K/v���7�_�7h�/�ɚԥ+���x�0�Pb�u�[&��e��ɫ�S"';S'��g�of�a��A�Oz�Ir)��z�|��{�������o���k�(!��u��m/b���T�d$���n >�=�c2YC��W��ww_���#�r-�2A><c���h_�,VZ�U��Ik/��K0�,+�!\�wҝ`[�0�G�
w�"�����[�8����U��k���,���&)%7@g��vx��==��ظ�S�ԐH�Sﶎ��E�A:�l$zLVO3��w��'�s	{\�e#�zN��\��S��� =B����>��f�v��_}�d}�xSxEZN����[/S�Q�x
���M����l\�����G'l_�����"bZ#�(p��U\Y����g�T�"@�=����W{#�,-�ў$/M?;p���d��t�5aGI�l����'�S+��[�=�v��
���Q�Y�8��	���2_��}��i�y�
���Ʌ>�B�xY����cB���f�);�oOF�}/�2��6r�^.���Bb�i��w�1CÇ\އ��$��sg��RvPZZ��2��h��1:ȭ�LLj�N����c���B0�:��s���]&��0���/9aT%�4bs~�o�����P�!��u{�tW��,b�}02D�{%��ow��ښu�^N���uͿ] ����.@�����4%��e�<���[L���5�XP�.����R�f��E��}Oa�~�) ��W��Oϫu)�=Pb�dN���}__йCh
S�����*�S�A��N9���N�Pv��H�3�(qX(�8p�0p0Imμ[�I�hQ�xؿae,+�����;R����s3��y�x���D�w�s�+?����n�Q��w+�_�䱢��$n��1rC�T��\~��pb��*��T���0�T#@"���F�sP@4vm�09�q̝�<)�qs�'��%0���~��&�/�����*����L��@�;����6X���}��#@�sP�z7=��RC��O�	I����"��3p��d���Z�	V�iFw�e�z�)S"��Rg�y"�鹖U�|
"Z��GCtm�Y{�!���|�t5i$��WE�%��:=�*&QH	���I��x����`��{�-ؾ�B��v1���k�R#pg�]��Պ�0��I�
�������yʂZ���*.k�=)���΅'���4y2����~�]���T^Y?��'����w�2�7�;C��i�>']ט��&�ՁX���P��&E�M�S\b�L��מ�Y=�y!#����eZ٥m'!�?:�����#�Π"����������}e:aJ�h`��).�����|풰%���Zo0�������@�U�8��pI5��Ͼ�T�gWj�m#מ5����]	�U�q�l��@�)��;��g��KKx�F�Vl��|r�ڭXa�? Ma����t��������g<�j����H)��k�u�l|B�����Po��k��f$s�+N*~X��q�;����!�q�S��-�U
��Q��'��O��
Y�C���%69*pM�X�$̫ޔ�/�,:�rzI>���QS
:�\�����:$+&&����Z&�⊔���ϫ��o���
/�������]�Y|�� K�́��������Q�� ��k��:�a��:�>)��wǨ�?�P���;�=[���}�n�S�d�+'��|�"
���h�7�n�w'�4�;_���I�R�k	�\70ܸ�\��3`W����=
�o``��+Qp3�����ّ?���|q��[<�Ŷ���88�>�t
	���IR�l-���5\Y���ɥ���.�݃ B><����c�ʫdը��+R�4F��-���]Ս�F�+��g��]�wW��/�9���7s^���]��t�t��������2�\�>��e"�Ŏa��B���2S���ȹ��M ���C�ڙ�8��07('��a��/26;�S�����?����D�.�F��wI�.Tt;�?���Ӂ��ZQ��A��n�`����=�p�ѥ�4ԗCB�D�iS���o	��+��S�����d��-��Y6�Y�Y�o��U`)s�d�����ۢ��I��!�K��;I?���#��N��Aw���V��h��"�At{XԕM+��4W(7������剋6�}�ވa�=Z=l'�v}�D���o��R������Uy�.(������ҤW�ȥ!NEL��
@��>�6ɭ0y<��0�w����T8` ��N��H�eOh����ǅ���N@k}5[uo�j׊���X�S�O��0��5U~@�"ԩee���x���4?��i���s1��I?���**ĴN8O�=L��� TQ�[ g�� ��2fR٩/Q/.��;�ؓ`��@�=�i��&U�T��ѯ
f]���)4W�'��ϧ�!��^BW��m�#r���)������V����)��%�s��U���[6�Q0��|�~
`�W�'Ń,� �r����Jw7�|�l8�yA.4b��J&��ط��(��	����ppH�X�2�W�~�du ;(�k
Q�B�~����)��sLU|��d !�P�W�#�SJ�S�@�p;�~c9�	jv��G`f�ڵ�kW���
jSԷu
n"����:��T���q�e�'�v�{��X�?�=��r�	�o�Wl ���YIW�Ĳ�&��,V=�+\e�9 ���*͟{��	'��!����LW��l!�M��*m���P?���,#;D�F�2T����L'�yӒ��ˊ��c9�U)�n��g�K�ZΉ�{�k9b^����d�s�2��s�ܷ�8����P���1���F���)9h���y�r�)RU�$���h�tj�R��^�Y��v�MG�O�J3��w8ry��*,�Z���&��7�z�_�؉�| ��@�%il%����u�M(��8<�('�,��,�-�v��~�h9g~Y3�+0���JX;]V�o��s�c7���`�CZ�r���h�UY@#Υ�)ʆ���=o�nrO�ts��s;�Y�lN�dS����ɸ:g$�8���י�nk�؍�H�.�8R4��G�W��٘G��ߋ�H�%�VK�,F�UA]�1��R�����.�����l�ƕק����)�����W.G�s.�Y�w�L�8;�s2�t�=G��d���﷧/G7��z�rD����
��k�|��6��Vu�>l��#:�r�X�hȉzH���~�k+����V��������ߟ4Y�ٔbqy�L���;��f�*���S��i�� z���BW���w��MM���\���9U�۔�kb��,#�18<D��n習/����ç=p�:�2iQ�k����#�Β�=�����4�t�u���
�P�Q�@0C��?M���m���uw���$uŨb�V�ۊ_(r��P� 5Z��*���_g�:^y��[�Mw�Lэ���TUe?�PB�v;��jCs�9�z�]����h3�CW�@��M5���������JT��\���
Vo��X���R�~[h�`�Q�����l1x�@��[�m�4���	��������2z��Elm�(�$.��s��"T�/� :`��g�}�8���"ˈYxRSӡIx��r/	K�)x9�ڣ���-3�}YWegËP-�ve�fa�n�J�T�rC�����)��U/�6ҕ��aS}$�NMN�GS�؜[�2��\b=':�z���/��gchUE�U53�|�x�RO^Rd����Ыu����Hܝzq#B���;U�(��h�|�oD������逩�de:�N7'ڛ��Z\��Xq�(�����~�0]�Ê��_��2�{/�'�|2iH�i]7���D�Ay�����ϗc��r	�XЯ���{%�s��{*�֏�v��=��uV:��;���;��:Ċ��ˑ�c�EW��N[��y����MJ�Ϳ��e&�^~}	%�v~���e��S
��@��@"�3e*a���>��f�D��	�\M׽�'u�"����,|ۋ�1^��OW�Si�f�^5G Eǀ���/t���G�$Zz�������2,��[B�����3��^bsm6|�l�����v� ��a�|�Q��%�o936�N%�<��me���4LP��v�L�=ss��r��(����T'���|�}-��ԝT3>M7�X�*��B�ŪJg}����f?�>rV���K~�O��^N�S�5q�U�>[xOw�O@������m��>x�����8%9��o���y�d�b*�$^�k�����q�u���Y=n����r�h=W��@^r��l,7<Meκ�漑�,-vGk�4��o�n�������	\j�&&�S�'��[9�d=�$,�q [ʟ'&�[�k��B�_�kڮ�J�c�-a>o,�:�w�u��~O�wJK����~*v������Ԋ�_b
�1iI�|�$�vb�Z@�VS���>��
��u-�HⱩϕ�G)�����g{X(xoLn56�����S�c_����Ba��k�f7�N���I��=!�Z�T���#����R�g�M9�ι�5`<���hdqik�5r���y�E���h"%-u�`����i�_��*��4���j6��z+F����EW�u��2?�̅U�(�uq�*�6��`j�z�=���򞈿��K�ʋn+h�A� ��c S숖���tE���m��ZcA���ٜ��Q��!��Ό��͟%w�;��h��Gi'v��̏��$���d2*�FZ���	��d��e_��U�c�L�������Z!3n�e�k1)��E��]/�����)%�֞�3RQ3�S�$��x�{C\���F���4됁�¯���:s<�e�����ˊ�A K�Lڳ��J�ۋ�Qa������ЇV\n��[e���D���J���
�!w^�^�Y�Ў~։�-�PJ%d�wL�n?_��+�S�r��1��%F\p��?
wEˠ���@�YA\�x?�V��2��sF�.�#��0��E����W'\,�>�����_w����8����[-Ut�e��]X�&>N�-��Z��#%�*��QJe��)h-=fQ�Gdە�D:e8�������p�H'�X�{Mo�3�2�\�-�|�#��Sdw�5��cG����M�X�,s�Ƹ�^���B��rRU'IDK�VL����S�Ů�ʑ�4���_��zA�5����,p.���K��+ʅ��⥟���+��I�$��:z�($�z_S�]�\�oPl������أ�%��-m��|/I-���ˎy��uJ>��Q���i��]>����IC4�l�ԝ����L��)�7�]HY!Ng�6�H=v�>�1�S��J�F�T�OV�!.�p�hc٬r�1�c���E��D�@�Bb1��	���;�U�-//|ɐ=�y�0�����=�[����Dm2�/J顔�TNw֫6��y�.M��}��J��ܺ��7}���9��X\Q͵��������8�#�ڰ8��:i�F߯��^�NFU�f�X1�%J�}�w3:�u���\����!���V�����h��O!�T�ĵ�x�dsk%��f��f�t��4����dDt�Vj���BpיrLkk-��c�"cϽ����ٓ�B^���,C�8[ׄgk��Z�FsT�j�l���!z�E:0[.�4W��+-XxB�B��I���&�@��%���6jZ�	;��e
34A�M��{[�X�;wշKG�/8���Ҋ�_f��0�a��X���/޼�e>2s)<���J]�]��?>��&(,r`��)���\���23���פ�eհ��6N�}�*d�����	�����=J�;٢�͆2�"���m��"�""n�̽㒶�&��T��$S#�I��8H��1w�!���!c������1�[��q� ��Y�	�s.$I��{{��VmKv���;j❓[��I�0���L���r��e���?�<k'2c�sW�����x�����J�xa��^�l������%ΛbJ��f��v�綿1�d?�A�R}�0�F�k�~�pW�)��"{X�بCs���y�>��๾�t��k�3�ƽ.[D��y�Q~�LGr�TR�K����4�}�%s��~�}j*��+�1Bg�rf�
-���c�'�������=�������E�Z�Ԗ�m[�SӼ�"�VrR1^�Q�n����!C��}b`����Fs�Ub�f�n{��-���XՓǎ�N��v0����Z����f2ʻ�sX��*B�|���ư����H�;�dkTs�K�'�j�5��uj�`��?��˺��C�%�1�]3���A:�ݚ�~��#���N���eY��]X�j�@�����3�����)��:�Y����	��7�T�<O���"�k��C[��\_�f53�.�eco��z���n��9Z��>�925�X��5.;���Ǡ�ޫ"��3�T��K��e�n�b�~���wWR&B�&2��Ѣ�S����7[���_�փ?�����y{(�G�)p��`K���bk�Rq���X�V��>��э�ޟ�P�߬�Y*��h&�	�̿i��9@����^
�Ԍ��KYN%���q�p��4�mw�X�\��޻.��9P���+إ\$�(�%
���m���҈7eb�qxԦ�����^.(b7�@���Hܞ��1�9H�i�IRz�0꒰�y�t�����Rz:���v(1�����m5N����L�_m�0J�b�]��Vf��Ւ@|ޒ��%*+[�i��}�a��B�3yl�5�j�����'��W�.�x>�]�l,��M�t�er���"�5'�htKQ'�r�d��N3(n�����f��+�a�ξ}l�붟�g����������8\����魙^.E[Z�
ڡ�|��5}�cl,U�u����E^E�s��R@�'��F13����e�b$�iM=[ٯe���添�ˌ���(S$�$�)o��f".��>@H�?��uf1�T [���b�?]����ѨJ��]����{���2!���5�i2�>aR!&C��b���߳9��Hqi7N^4��.y���h����c
�|�!�?z��1IkiIYm�|�[��������HlM2ٳ��4�� ���+�-�c��r\��X�f[3L��p�;(bv�kavQjT���ǻa��!���a+����[x��;��b֔�_����՗̱�x��v<��v���\D�j���xg8�d�ѫǚ䪃�q�����>���=Yb>��B��dX,��[*������A��v�莨w]��p��ǖ"5���a/���[�}�Y/�3��8�FpfN_�x�;����&�_K��d���᜚��	[��E?�=����/��6WN����UX~{��rw=v�1Ps����h0��i���d2*�u;֮����B�vߏ@���K~�U�i�U�Io���%	�'�D.����A>8�p�	Er�%>�~4%a�YX����G�~��mwд���i0K��Ihzx[xRќ{4���OV���WBn�X�z���,���U2�&��2�ɸ,����ڋ�慅��ig���f�(?��*v�y_4��b�n���?VF>}�rާ<��UH��Ug��w��R�"T�'qT1C�jI�Ӣ7�ʽ��ߖXqkQq��D0:X*��봳�ވw�����v���Wq�WAnr��aC�J�g&p9�JPF����Ut�+�������F]�SI��Y���&��>��7�m�w��M�;�%�R�'��;L+쭧�$Ó�/�mkmM}����'��^J��\��d�_Y�V)ݕ�S噾�Ǭ��O��A��;*��C��c�~|�	j/�EA�֓
=n�c<<R��rH�����e�ЮP��g0C��n�V�o�������-*������`�l���h������B���8 �Ǔ
7�P�5�Ɲ�������=����Vf)��4�������~��G�~ :	��S�ʅ��XGi��Y��h�<oꇸ�=q5��1���F�GF�����������C,���.]��'�Gc'(m:*󗹾�=s����ܸ��j��wN��S������Ű��X��/I��	�0�����r;�_Ɍ�&d�8;�~y'�)��ocE��;���?=�rvo���H�t;z�)s���c�D4��J�/��@��}VQ��B�ʱ���7��E=z3��ٚ��8�H���a.�޶fc�5�E�9���%��8(rkV�s�X���cJ��Z��~zO���3=+ l�ԝ��c< [����j��辕LO��8�,X����r�B�u�u�R\�fO�z�����sf���B��{X�	��!��G�U���E���U��f��mDf��5�Lܽ��/��-5T��o`�t9�/j~�h���-
��΅��z�pv,��4V\�����ffl�4��a�Y#��1��s쮀�C"���s�
Ųm�M�Y��Б��9]i��"x7|�r����w�]���������Ǽ�������������_O��U��-�=G���E������N?$�ȯ�3ʧ���bk��}�i�0"s��o�gu�obe�CoGE�4PI�A�t^��vo���wv�hW�a�!�?�5�CZ�Mȍ�[9y�ćp���lTK�v�$1�n7���4�*�Hqơ��b���J��S��z���)wo����&&o>�V��mf�f�#G50�+�	�q��G񲃚[�0�7�g�M$�iD�<1~���I1�w����bb�d�E{*��*E����Kdajxӱ$N�p�,T��őJ�J��g|��:��rx�Z�ƪ���*?�հ��l��Y��;��ZFH�D������n��[���͟.k_�j��J_��#\����G�/~��9��ymӚ�7`�6TV7��2�4����N1{�5��JL��#on��kj����ᡢ�&�P��*A��³Ғ�_F�|����\�4R� �;��@"U��N?�I��*�r�?Z]ɸs�@�����>�F��vt���Ei*9�TS'�0Ƌ'I�m~L98$7�TC�;��{�k���r	M�Wlo���pH�j}L����l��	���c����|BT��b\)��װ��{V� ѕ���^k�=��_�AQVP½>�RF
��qݖ-��ƨN��M�]�vJ�"xX���P����s����ȁ�#�/fd�p��P;�S�5��	���L�[�@&я�,�t��D���0��mDt��!�6�W+������S���^��۾��\�K���B�e9rP�7���$�*uh�1��GC��]XW����U�Y����@��O�rnU����r���+��:X�e�SJLWcc\�I�S�8zǩ�f��W�B���U|[|P�q��90rV�x-*��U��n�J���/ݣ�}��:�*�ۉ)_"j�2��Q%��+��p_#Y�����R���+��	��hu7�	s��l��a��(a���[�K�q͙z'��>�c\�E�<^�1I�m@5,�18U���W�-"hϳ�r7m��9��`TI&�p_¼�����<e.���:e��
"ˠ�jF�<�4M������F����B��/Csl0T)Y�_�]ϙ���h���|�d�a.������;0��_蠴��8���L�\����:{n�L����]Y��.W�Q�k8��&�A��㼴�[F��-���lܮ�����g#���CO�:m�����e}��0�|�jDf2'h,�w݋\)wV�:��mo�b��~�.�[<�m��5��$�0�-�@�>��WH�i��.�WP�8�b���l������f����1^fb_�7��5=�A3D� �C�����#��K_��ǟ����ۻ�\<%3C>9bCo�mˈUI%̞E�_�Wu�X�G�"���To��O��VP�a�A�*b�"4প��-��{����D�r�Q��f�f�!���r�DH�j)P���_�E���T��4�9�̩����!|+��}��L���K��>7��gI�O� Ύc���>�q I�kػ�s����\w�w�}�EUTn�r��S����$��m���[�T�v����Sr��=�`���MO�%�oU��̔0��y�2E���[Y)��JU�o'���:���o�4}e 9����X	)Z5|`��w�^*��M���������0R91����;�{��_����
����t�,jt_��Y��A�0�a�B��r��+���L��l�1:Dm����12n�rg� �A�ۿ���|ퟩø�	>�$�M4I���XDp{��:::���/��@��{c��e�U�K�c�ۛίzk�v����9~�*�&���u�F�-$T�@t4�F�cd�BoGO^<tx%U�VI������3�%��2XX��Rnm�^��JM��Q��jȃR?u
f�)�K�KuB��#�����݄O�/++�}w�[�ρ�A�Ɖ��8�ǰ���Q�0��V����)E~��E�з����;��Z�0�M�`$�"�x�e�tu� �V���a�h�ذh��s���W���N%�о��*��p�c���G�H����Z ��"���'��}K�0�(%a�Z��uy@������
6�H��\_���?Tgdd��a���C8���p&�+�MX�[�׶��}��\���p	��[����= �=�!�,%�
4�ˣ8d^�5��ϛ�,���V���"��1�r��u��-F�R��{��Z܉X��*�Ճ����}�;�po���\I��g�)���������RUF��"��Bㆱ�è2��=�_C����Hs��,(BNz��Ek�4��ٲ�h�‐�J���.�y�꠼v���F>!���#����V��L��ԍXg���!숗�.��$��Hռ��H�	n�Xd�9�r���m�gЧΆY����;}Ō����-(D&��:�	U<Vg~��n���{χ�,v1�+�5��*�(,�0�/c� �!ܪa�5�Wb�{��,���%���.�{~���-i�ְ����m��xZ׽,��������_�V�[J�Q��rN%U����Z�)\o��R���ZC�>�9Y�����Ǉ��Mվ_���WK��ZQ'M�d�}?o0�?0��������ʻb��s����	XZ'ki."����Bw�tu��5��v7�H06�c2�4i7�q������3��m� �.<��<�;Й�����C�ɁZ�#FK�lP2Jv��Z?B��] ��k�(7�ɡbd�Bm��:k�Th$��8�L�)N�k�� �Ĳo��[������7_�&�qI`�g��ώ������j�F�'�K�4��Ƞǩe��22Pz�����|�O�RQ�G^�tčZpuD�$�̾�on�PL��2GG;8׶H�JGY@ ��4���4�;Mu\`�V�$:/�Ý4�f�J�=������Lk��d�5�uվ-�p��%�LN$5�E�U��bϯ�ӛزՆ�gӔ�J��;�ƶ�L#���m�j��!��o�$�_�Y����b?PT���8h`u�o�`�_bYJB�i�?�9.�\{�tw%�Zx^T��;7�(j�{�
S�Fo;$e'�$���I�QOi�q��]i/Lmmj��RgZ������k�b|7���KLz�m���)�.�ڂ�w俿H6�K�y���x@ZC
��A��,Z������^#c�;J���*|:>,j��	�3�Q��EUMr�0/�}�9�z�ϳ�$>>���Ϸ<El�0��*�x `Ƹ���l�UY��@�c��*��岾��3�-����(Ki��1A��z����G=oG�T�2�Cs��g�P �<xS���|N<�
!L]��oV��V��<��)ϨO��a���m�]�� r�'�F?��!�8���~FHXQ=} �s��]d�,�c
ך>�I�i��990Q�V��t���[�.XwSV�$[^��8g5Gdn�*��_6��)�Sx��B!���L)���S6q������"�>�v�vc��)����
z�����f}��&O(�@���J^��4����d����vҏ�u����k*b)�u��elD����ăhO��㙚�b�����̕����:�Z�(��R�&����g�Է��T-�P�9���F�[��qf�	��ᰂ�p�
�ж��$�;A���ˇ�=�U;ǗMc����uהX�\*5���I;#J�2�z(�i#IQb�]C5lQ���k>�k�g��(iFҹC����
��pN�7Y���Em���70xM)�; L�^HM[t2�1M�K +Q�C����Z�E4^(��̦��1s�?-&��	2/��F2�M�<0�A���&	������wu�y磌�R�!��q}-�IC2O�'���tW�z�Q/neU"����p��2�T=���Vŭdwk9��>@��(I{?X6�5��OF�kD?21[���� ,���RRx
u�2]���Y�y�$�v����XI���*��|\³^�V��Aӏ-�e�IjJ�o�ȿ�)���5lv_�ax�VV
�Jߊ��$�$1@"�p�{OѸo��T��4�O�^\uHT�5�T�{��<-~��X����vkP@\�e�:�ފ�v�b��o ߺ�>2�ٌj2��d��ET��Q��'�$�������px�(�(&I���M0�ǅw��Z}��kJw�p�m6@��X�+��J���8&�X��:�%e�0u�{�Vk!�`ySоt���]�9�=��+_�u���"Ҡ
�0�ˉ�[�sK,6n�	7�8�a֗���~�i�1��Nw�~�}����Gף�Չaz���ݢ��O�Sfޅ�L��B��2%J�c*�(U)u|�N��_�m�1>pb-s�@�Iuz�4���~sm߶��afs���\#���Rm�w��M<J�K��/s��qB8�E!r2��,�a��}ȑ��1� �*!?v�ܙr��	p5�))�c��$�|���'U�V��Ҵp��Ju�tYOO���K$�u
��c���Wf��*����'�I).
�`jW�APS`L�%�dXK��[�U�b#^�P�}���M���t�{��1화��As�F.�ݓ ��������|K�kb�#��m���=���K����]�c�_�mX�^��0%mz ��L���r���x.w�J<�c݅�b���22Z��?��19�YQ�[��f$�`��I�����!��}&���]�Y-�:a�beͯ�����|Qnfj||��b��x�f��h��Ԥ98��Ql��zmzg>������#�ǅʱ�â2�eg���چ��|ô|���2������m/U�s>�޺��a8�t����^/��vwc��������GyOi<~��D��k�Y��n�.��j�؋�5[|/��zL�.3�\㊇�#�΁�,��o�q}�3���}x�0M�	�O���n��[���ɺv�yU��>"�B���YhÈ������_	��C�ċ�#sg\�_���Y�L�w��44��%�QV��o�In��j��T�\;6����2�7���ސ��O݂zρE6�wۖU� �������F�=�m�XŐ��Գ^�͸t�$S�VN��o6����D����a�=ϹMJf�|y�0�k�W��;�/�^����T)�����x����#�toESB�.�$���X��A�4��#dɾ��)c���Dcߗ1L7KY#��F�6c��}0��=�=��k���~�����>�s�	�\~�Ϛ!�� �}�O���R��dyQfz���]�'��LW���5�gE}�=����&U$aJK�\��\�K�!�X�&X�����?iI�T.��J��ϒA�űI޹.H����}Vo$���w����o5��,=�W'�+4,�A(�~=ۏ�͢���������߸ʊ���[�^�����]rFs��s��>��t5�2��F�Ks��0>q�,��Q�Eӽ��}]�c��Y{w�"z[8ո�?/�=�����V��piN�# �:x�������b�'�7ƿ}K�G�}^a�2$)��Χv���
���c9��D�jC2�/x��2�Z�ܪ���1��nt�w����OrΧc�9=��oz��E���4$�Z�3$t�w�E\!���M�� ��1uB��ϟ��3zRb=��ʜs��ejR	�3�1ua5s�.�M]:|�|�k"A�+��Y�2*��� �p;ZϚv!��� ��+�q�ݙo���ʯ�ҋ�(���sھ�̴l���<������os�Q�酊/���� Q�UtU�绯�7�Z�+��#[g_��S��ٺ�;�jMr~J����
r�W+�����ޒt�|{��ٖs�أ�:�����1�����k3��eU�d.~�3A�N�ִ���Â̞O�C3�g��q����ГNp�0���'>0��"��ᥒ}4������pâ�!��X3ʱ�2�>1�/�K���4�|b"Z�G��d���7��|Ce��-�U+�N،����{��_�E��~*O�c3���>z6POeM��AU��x��V�OY5Ŵ�z���BH~���2$%����ů8r�ɲG�(*+q�$ܡ��q������E���p�8V:hT��P�~�=,��忦�,��Sy�U�,Ob���aMaP�N~-g���W
���I拷Iʔ��PR�|�cI6kP�nv��;]r�*���z5L�Ny�#2	9+C/j~O���1�4�E�O�֨�v&�*�������潘�x/.f�<=E�N�Ȧƹ����5Z:Q#�턬������/a�'e�i��iOY��Q9�%^�������)��O7�Kxϸ�hqNq^�����n�H�4���5���ϗ)xC@�_�"��R>2z���Z4�A��`SE��Ňg��.khE���͕G^�O|O��60�'^�V���v���$��Ii!� ��v%0�1�W��2��©b1����&�9�<3��S�z�����R*�7�x��ܖn
�bWex��=��U32�\�5�o�W������(2ĕ�}�^��n�։٥�	J��\�
�lno,5��!��z�m�����TA����%Ӗ�
�o�>$퇈d�J�����������9U��cV*�U�������	��WZ1�1�{���C�)�%&��f�n�®g��ӽTPn?�CF'��kEҎ�wFX'�v9n>�i����������MP`-?˅��H�-B>z�.���;C�g��C�~^o����K�7A��|F�%�.͍�>��@���6�9P�D���y��^��(
PW�DM|m8y����-�~�D6���'��@P8E�K��ceޜU��A%���v��/�z���8?������D�N�g�H�����������R��޷�������ߗw��,��p���m���vx�N2�s�M1=Z�j.�J�>z�+>��<�x���:ZQ<|� ��ۄYj���j!�ϙ����u{��`Ǘ�f�b޼�����퍼���;�ʯ�L.Ȭ,Cվ�yժ�ɩ�V�E���c�=�=���;U�-W���K�?�`?��#�P�z�տS�IK-�V����T�c����� �4�"o���!�Rh?oί��tN�٥`YژVf�!e=�N���'�n��KJ��#s<
*>+TÎ�W���e���KS7�~��2�^�\\���Y���U�%���0M0����CdШ/^�����xE��?�������y/r�ŖcrIa��?х���,��
��eX���WϦ���+�<�_��LձX��ޅ����?�Q.��ڿ}�JqԻ��O*�Iȅ9�������`m�M��h0��'b�����G�\ș$��8~�J��*(0vM��y臙��#�K~�0�gKs���m�B�7H�{>�����u?	᭸����f���#��_��\�G�<��˅�s0r�=X:����#3�9T�g0�,e�'�_�H�`(GG �z�f�3b������r#�@yiҥe��]����(�
;r'%W�{�~� %�J��/߹P�R&���^�S{C�V��W���pE�����z�a��m̓��s�f�P`�N�y&���ax�c$6p���ܷ9HCߓ$K��d�K�Z���������Vw�%�>��Y�e� �%��X��ޥ�6���z� ��41߸��݄^����W�,�[~�s��3ٷz�*'��{�8+S�0~�
�Y�FK;ާ)�!��I1{��hM
��q���c��`p3.}�R]4IYf��YK���
��ER.���X�7=�S�J���
m:�~���\�|?H�1  ��%��o-	�DF�Zp�:{�3R\6�L\�f��] =J�=Jrқ7��w�I8��qC�_$�RP@)v��X�������]�^G��$E��<���|��H��b2
��y�}xZ�Ύ0r�nډ��ö��S���r�J��j��: ���\PD��/O�1�F>D��uϒ�������H���]v�
�ݦk�����ң��
����⇡��L%=i�����GA y�t�����n*B����9� ��mc/��6+��f_��������kν�d��' ��b���_��p�^�,zB���\���*�d�c<�D���5�KS�־���4/t�{`�l�8k��ci�(BCv Z�
ɀ_����R��ZL���腀�x��#Z�ׄ[h��h�f����ܿ���rL�:��Rw9���c�[!�lWq2.T�>�j{Rl�ͻ�HP�Z(>�a�i�v�F+���<��r�n��u��5�9v�I,:��1{d��rj��ndj��r�-���o�s�� ��o�v:m���Q�r���nhB��9������5J�{
x�?��E��� �	�:�+W�zד�%��j`��@��YYT��..~�d�qáb���0Q�E�9qԅ}�5��D�y��.Ҹ�#H&�9	%������B4ib�:=Ĝ�ӈ�<����t,�\�Sȵ���xuҼL�۱J�� �R�z���<�3��-	�Eq�������H�ǌ�\SD\��X��7���2X�VQ��x������w-'����R�0�)ڸ$�SkB9��`�A�0�:�����D�]O�.7���S>�X�/P�nC]jn=�����ɵ���ɿ��3X�I�U� 8}�X�v�e7��#@设�+��;19�ۊ��tM꙯�l�i� ��S���,ڀV�*�����jkn>��ي$���xY�2����AE��E\Y���!������f�����j�!��IB��}�u�ލ;�\7����Աw)��rJ�-pf�1C0�1i$��[ik	�������F��	:fS2}e�{��AX,lݙ�����_�]�Ox>���
H��qs����c?�q��x+�9�
)z��ӟ$�?�y���A�F��N��CWɋ�Uy/�է���&��v~�f(
��	g��W���j��3N3X0�G���Dn.�SB�B�?�����M���e���@D	4=���� �({/�x�I4A���~9��>-k~���:�B;���K��5��^�tS�S�`�%*H�;Q���$�<Y��ʙ#?�6��衚�Y��r��^�kE0ךlu�?���ޗ�8�,4�u>͟�������e��@�/��,7���8�2�� ��dLC��V�p}L��X�I u�4�O��ۯ̗��|k�����ЏK���j=�W/�@%��		��<#�&��!�uS�Ŗ���o̊6$���kf�ܐ���|����]�j��$>���!��9n4���b�;�k�+ �s����F�[O,"�eM�@��V���Q�@�R횦�� z�9�'*p��`~��rfL�]ٰ��ռI1����F�+e �
\�w�ڃqN_?���RB��9O&H���ƀ�Ύr�⋔3K�u���Ę�B�&��V���,>Zq���T��駓-�
�C�'*f:�z��x�O}0M��x��U�h� ���D6`ј��O��D$�J�h�9>��aJ���,K��)���x�s��yh�A\s�㉷^E�W���␡6��9�-�^F��2ʋ�<�i)lÈ�����8���!.�f�T�ςe�x��c���F�}[�U�"�Y除�YW�+�t3�G���v��i {9,{ι����o�s�h����!Q1�.KX��1(\�&
?�n���o�<�i����Փ�Jn�ǅ0,7؄�N1W0�u�P
�aP}�����?�KRf��픢���]'rD���j�Z��?֪��k�r���+m&*��Y�� �nf�:L�g����[�}�����h񉷻�#�g�Jd���s����ꇉ�V��[�˪p<A0��o'�����\���g�Y��$�~�*�F&1ut���� o+���jfu;`���ݬQ�������9%{H�<F��6�l�3+wً1_@V�"��r��-0e��{ιx�۔���EJe���cR?S�c�7�]��ʀ#�M���LZH�LE�L���`�A��6&]���ߦ�ʆ�����T��8Yx��xGx�8 ���5����!R�	D�d^� ۞�c���|c����]��K�d\跥���G�]����
�8OX� ��A�k�R�����c��!����U�R�x���h'v��G.��L�C_B��7��0���� ���*����,�P���]�+��w:��s�i��K�S��C�$��rE��^�U*��]�o[��|���Ǵ�*#�����aG�J�'8�岁2�^WӃ�J�����k�eE5zi�U�t�U��*x:	V�#��[���
ڧ�$�0�y
y�ַl]�Xw�V�Q����?�G�:Y<8!��S��m�f�p�� �yDԘAeI���枙�|4�{�P8�x�R���7o�ϳ*zGlF�4��d��虗-:;f[<h���@�|�<~|��Z)��ڤM�Q���"����<�5gU�����\]������ʢ]���Y�g�@k~d��nvveS���]l[���~e@� �4���DVU}a��5��&)�!��`C��	�%�ρ}��g��H{���+���0��+i�B�D�)f��
b���!�!
D���6gw�B�(�R�|���6%.��5����UF���_4X3�&����O������]�Gi����A��d9�vw��r��z_'�g1R����]�1���n���"�:�=F�}���5?i���s��O���l�{���=6.IqV�ٟ@0�:��IT��2�ww/���2=�5J"�c�T�k�Z�����a�A����qZ�Ni����[Y��tI�199��ix�o��7w�U_��\���ѝ7|t4��t:��]�-�}�q�O����3g��봥����/Z=;	q4!I�_�8F1��l�ؘ?���׬��9�l�<������+D��/�+m��ʯč@�>�r�a�^�-����y+<�q�'�'(�cq�:�D�PJa���y�`�r�����s�i���,�S-k��X����{*\�.?�}G@�RAOe��g���d���A��)�BZ�*};��V&���R��؈l>���x����˞D Z�m�C�Wy��\�Z�\�Z�^}6U�N5�����wp�uPa{�:<���g{��;q��	0��?��Z�AlO��=D��)?MS���LR{�~mB�����@���L�����d�v� ��A����S����I�Ei:��W2�β��姰7y�/�� f�ݡ�i*Y|h�"��]�� ���۪w������5<�^��|�]��sύI��,S"�y�HZ��,z��D�պk��y�]���!��L�jZ5���J*�&/� #0:�g6w'�wy&�ѓb��5�7sy��8�u5!�v���K�����u�'��J�2�������҂��7>.8f|�Ͽ�s;��m����W��@+:`��k�~�lX�L�і��჈U��ҥb��2�M/��i�㓕��͸��%����T)�fmUsCy��jmk�TA�4+x~���e--U��<�l�4�O�u�����b�廔�A:��rd�[$ة�ؕ[�2�r���hta�g<7i9q��T��Z���h[�]���=M�Uv6���2fha�HE�M��y�M9ޔ��_.D���8Uj�w����O�&A�� j���9��ު���n-Ҷ"Ezk���N|�p)��$�rnW�E�|3���~�w��U��MY	C�9�_n�9�[�X�J���|>g�.V�Z%��6"�6�s�EׅU�w��$jq�,�t:� ��8��1q<.�jд�jh�n6���&��l���(��8�9����8���u����̬�L���L?������U^��ټ���DD�����K�5�*>Z�vuf՜��W��E��4Ld������|��M?�f|^�AB�_6���9F=,$�=h��m�H��RVMt��54�\��_���.���'L-2/���͙bUf!�/���ȅ*��#_~�& �0t�(�����7@Q�wK�#IW�a���׿�n�v�ru�}LD�o���)Skw0����!:���I�Pm�Y�x�̹�v.H@����[X����+�vi�;��E��v��=���Ɏ�u��ۉ�u���&qrɊ�@�v�=�a��jhͅ�RmZ�e���}οó��Y=h?ߜ� ��"hU��3E�*2��"��|ҰC'����YR�d8��ޟ8��C�U�u,��?��M���k��^����P,i���Yu����S���Nf��4.�zS�,���N��m�Y D�,̇���s��� �E��A�P'ZlZ��I0�������\Ȅ(��d�X�z#�Ͱ���ĿŽ`4Y����#E���{55�R��zY���[�J➿@�Nv;�Ԑ�y[���~��.>�,`��D�UUԸ�ǬէO�1ԇ�<�d�ݕ��\�q�����T�XEO ������DW�.co�wֱ�yJ?�;s���*ѯ/r��T���Ͼ�����X��<D�@�J�T	5�M��H=��i�Ȋ�_]F�'+9M�$�x��UUk�Մ�\���ߥ���/�	 i�����p�]i�S��z�n��+�0/c�W{��e��n�	Q�ꋔ�낥W�����nM����g����BO�,��ή���iM���&�z���:VcS�+߆7�N��}�
�Mg70]�-�ﷺ{�X��2b�̢��I:�Ĝ�}��Fi���¸��װN8u�oT�W���_8��lH�׵9!�?������DGZ��o��g��7��i! �@o�Z��%�\�ʻG:�EhH�Hl&�6!����=P�0$�˷O�\�+�q򈦘<�uSLC%�E�����F9U�@'�1w�q)~z+���7x̥���k��vאU#&���${����ⓛ�|�i$���SG��7�v.�p����q��Xk*��c�$�O̝�ٲ����Q��-�By{���_t2}]^�7��	ߚz��_\j��=j݈�#�������Niq��V�������ס ���]$���B�k��P�(���6<��p�����>	[p�-u��d��nn���݋������W��R��#=ཌ��S4K��"�v��E�^A��f�
��m�X�4�W/ h������;����� ܤ�t����6��/�	&����/J�R��wi�j�����9��!�ꘈ�'E�)��"_�?�����!$*x���bN{2���V�ur�&�C#>y�r����,+�0���E���;��~��]����ϔZ�.� r���|���"��L�5��WL���5>��,|���4=�tY�~����Ö���Y���7�W�ߖ�V�����]�F::�bL����nށƥ���v���n7�'d�1�F��"Q�$X���,rp��}a�$B��e�����
��+�T{�X�q`!Q] 斦���]�����,c*O�N�сϚd��g���H��҉}�*Y����̌�ѣӮB�xC��MV��&
�l�
����K�I�U�?t�]nP���J��AR\Do�qf�xp�q5x�d�k^� m"��q���zZ'�w��[o�m�*���o�Q�q~���2����y ���@������	d��m���.z�G'Rp��O�-������	h���&�}�� 0��%I�	�j�&#���sN�=�X,s��i .�)"㗇�7����%�(��i�e�Eg"9TFA��E����=��l��U��6��Q���5R���K���N��>��a��d��6����|g�i���v苧�i���*�g�L	�g'��`�~l�)s�|<|�o�۫��,���8/�v�@9����#�ΈЏ�@�~�q�ǰY�i��̉ZN_��Kc{�	���˼�S��B�؁��:[�?R@��Iyr66<�΀���H4��P#^8@��x��|}�̌g�����T~)�:���s����;�D�b�O�m-$�=�>,��r��Z�玪�a+Z�瘠'7*�S�[�H~%j�o��}r�+�°)��:�r���hx�)_�2������U��l�a����y�%��aO�b��Y3��
����x��y�� �4V��2�cj������(Dˋ�?�f����g��Y$�:��eWߑ�~���i��_��W5ե]�*IX~�9���-ڤ��0�^�[�`P���L�l��G�]����L֧)�Iqr����L ��)2}��c��!�&ʵ�]�����-Z�z뺻���ؒ��U�eT��-��pݱhpC�B�o)�+�W��[��-��3�?*i_X��\>VnTs��_  ���+) ����t��°<��k����p��l|�~�D��C͖[�  vz#��ed�]M�a`e�jD�p��뇩j��2�a�Vq���6b�PL�s4���7o�@wh�ȷ*[��G%�u�#����.	=�}J�XU"�ov��ā$��[)g��TQ�X܊��:d���ѠV��X�Msar䃽'C'Ƭꦺ6<��A%���-s��	�Y��a����ؙN{��E���O�4�ܧ1Y�p9�c�u�%�R�|��&�զ���W��׽�E﮼��(���	�2�������yft�!��3�G�mW*����ߔ�TU������~���c��|`��N�����5Sl�_JL�wm�Xf����lkk3-q�[a������8���I�� �#�G��)����h��C�DY<�?I�V]��ٻ{6���9V7����$����{�]L�&]fJ�hψj��Je=�V��A��v�4W#*����uP!����V(V�zm>���G�ؽQ(Tm�enS�5�,���hyg��zd!A˟���շ����$1I��@��ė�Y�����Fh*��$=D�bg����̞�4b*�#�J�Q_pK@�5�[K�vhf��O���'R�F���@����|b��X.���6��L�y���a�^^�/^���0�J��ʛ�"��itO��$�o6��% ��gv�x�-�Q��&ʔ�(����b#�/'��CTҝ�֎�+����u�߇��3��w��O��>�B�D	�����wB��=v�萾�3�Σfs��Kl�V(,� ����门�qu��1t�1�ux�*{��5��X�B�p�h����5�����0#���/���ԫD��?{;���\�R���W	��;�m�/�
��[-'+K��=)(�C�G�r~��]���_3v�U�1YQ��*���:ni\֟U��מv��j��]	C�j���.���~��j�K)����/�P���'��C��{f���wYШ� �=���]����UV�F�����!������eO��4n�.�<�{�O�[���D+��j�iO{I����0��p��U��_I[}=��4��dWu�8�V����t�O�+��%���KU��<0}P	��X���Bf�Z�n����L��)4�K[�`��3m��
�eȂ�e�
sH� V�}�B�/�M���{��!�*ꆬa��zb�"7�q��'�n,%�ڬՠ|%x��SJ~wu��mvA�8��)�N�@����:JJL�\�O����T�E@���2q���O!���&9`�6-.E�6s���}��3�6�1�8��d`[� 7[�s�n��	{N�'aT�;:.���:�+�*��yF �h/ԓ"�;S�}�?�2Y������L�o��bC�3b�˴�sV���=&YU��=��8�_��q�)b�z����z\(a�'M��D�.�"}ݫ�w�����`|E��P�\f�6 �&�%�o����?_�~��,tI��W��jm�8~�픍��ջ��@��OV4/D���\ ��Ehv�]��*H��P�!�^�¸��Eoa��&��?�xC$��WV�͹�r� �),�?WsY��#��]�v�&��ļG�F�X�\!�Nl�R�w0r���Uh}�����O��tzz�,�!��c�/�լ�8�%�ކ$�L�G�)���}A-w@&���7�Ȧ�l����٫Հ��?��������h�Gӆ\����?b���+_Mj��@6fǬ�a�$�Po�#���d�ݲ)��/��l�ɝ�O1]}ZN�ZV�1{}�`w_;�ߦ-�,�̨��iw�NF�o�~�l��R{��D���H��̭"��uX�ҫ�ЛFװ0<H��ȶ�]>z�
���j��2�ۨ�y%�u��R��¤�<��R><�A?z� ��ߢ��r�u�b`�;��B04�I�A�+��a��'���3��y �ֵ�-��Ū��Q��(6�qz�][�*�����\����{�k����>!������]\I���r��MJ������tN�h��x���b�4�+�FKx�S��,%�M�_�1vm�]
++��]޻���"�#�O�sC���U�U���b��i��<�v���b�+�N�>��a�K��ij��N��z�dg��f*������?BFy<� ���m�I��@k#1����P{*���R�����e
z�˾,W�Z�G���>��9��򾠏�b�5�a��o���G���Q�);�f�\�"eu)Ucˣ����ن}%�|�6��}�L�)|23]Up���i�2_�uU��k�&G�) �D���F��=�|�>M�k&�P}�YXE������.�CӯsoO!}�u�-�c�����1c�����5�"��*���@��޹����A�}���]������\v�����9��N�i�֩*L��p� RH@`i���!).bn5y��w샹W3��7�9c$XPw�o2C\�MI�]g��PX��0e�:J7[�x�,��,C.��6�\ґe����مAʄ`��^I�6�{��l� ����	��ȝ��߫n��ڍy6��D ��+6GC�S-�'����^��G� �p)��M�[���)�BJ���n	|�~�.��t՗�j�qm��)�>hSd�� �4��رQ���i�8��ɉ0�+_/%��22��O�b:���I��7���Q%�/h^��u�(Eζm��٥���O�˶x(=~��x�tY���.������������'~}׋ ;�U�g7�K����P0��3�Xߛ|w���gh�L����ď�#!�t����Qt�O��������1��Ha%^�o��f��g�l�y���(Q�b��/����������\��x�A��;`����>1ː���>�,}�1�t���Z{��뗕��yj4��&����TJ�1N�^�-�I� �ׁ��)��#
�����r���� �Q���ӂK���eb�� ��  0����x���̞��?����=i�t�mڠ{�֦�E���TC?(Z���j�S���P-�7vC~Q}��6���-T��N,�O�_R���.�8���xO��Y� �W�W���L�@��A��j<�ā�V�P���F�1P����P9�s�z�j��n�vé���g}�F�;_У�QD�^~��S��څ2���o�O���1G)ڛ>����ȭxO�X�<:�hz2:���]K<6?���A5���������D��D� � t�!l�{"wk]3������f��w�#�sr��̾��m���M�H��%�cZ1+�7�X����g��D�����h�L��1���!X���t������ ɯHEa)���-����B{�E��m��F�����o �SB�5e���o��[��o|Ȭ�I	vf˃���cc��A!U(�p�^��@�Ö��C�t'5����Q3�U�۽c���G��e~�&ml�Qpsb����J�hf$n��Z�L͵�f������Owa�?������0l;�}��L��b�O�����%�{�
TN˙#����(�<�?r�]�LU]m��40�k�1NY�/?n��j1<H���jQ�s=�u{!�>D;e9/az��L�,Hn��މ	�,�ns�^�޲��mÕ��yEhD/��H��@i@`�G�$n"���ښj�ѹ�@�<dzI'�0��"0�i�/A�0��|a�7��#<�6A#���>
�K��a�p���S,�H��m��,��bA��� e�y5ڪa)�\?`�ڤV{zx,a���[{�ɤ�������bv���Gg�MĘ�̋�����ۄȑ���ꎼݪ�l��Z��c$��ݱ�֧m���Z,b�����sx�[��̯V� �;�5װA�M�Û%�Fd�A�����NA�H���8�g
����bqnN�� ؂��rT�B�O�(�z1*=�y6�80��}p;S#�=���B/�@1�+���d���"K�f���Sҿo\~8�HK��g�sv��d-}2����@�|y�N��'��E44�l���?c�����K $2^ nwj�����/��x��r�~6�!�`y=�̀�?l *_�_3΃�__����(>�6gVU\�K��2a �3�j�e?�i�����`6��'�x�6�r6+���EW�o�d����j�$�4D�2S�[����|f� .���7�2*�Vt�쟽%�e��@���6 
g]�9
]J��������q�a��NM�����Ksﬔxj�c�Ŀ�+Z��ڀ�W���;e1�4�S�K�K�-��9y��w8l�s�4m�YnP��}	��^l�j���fS����Z�Mj6�3�0�j;��bY��wL� ����NB������\��:�:��#]�m����@�l�9*ө�\s՟W��Q�#�S7�G�n�s4�� 4|:�����hmd���")�fo�D��?goO��p"6�V#���}��Х0@z�Ϥ�{'�������U�.�S�vw���[)�7ܟ���������5_�NNjGW�:�����S�Z�0�m�odE���˹�t�G�����kx롲�i�d��V**/S}��p���Ҋ�Mz/��N�f��a�T�tb�M�}�0?bfBy���!\֞҃�r�~DA�N|Ed�vE��~��PY�i��_����;�f�U�k��,^D`(i�[i�O��G2%�Wy��y�P���Q���{��	2;�!z�����7:�/.Ø3�8��_��)��EZ�S3���hVt&���}z��O^���E.L������:�Q{��ѵ(��yD:ʓAtf��g���DZY�%#.Q��;�#��ZnnzC:�����&E��,@� "�O�~[�Y�d��\or=q�:~�S�#�U����5�4/2'T�_�33��5�$L�m�\��.y�z�=sx��No�D6� F��%aX4����}ޡ���P<]Iz?]��`�s�;n���H@�v����omC�	��ɘ�q�R'�d��Y�O7�����"0ŹC܂&%C��l�@��]���	^�$�S�q�[���p^M�`�}��K���B���^�� ,��SE���}��VP�*�Z�R�LKC��;/�'�}��ku����__k��n��12�����%;�N�����w�`�P\��gKǮ����'S�`F��$��;��P�\�=
�F�F+�z,������@Q���{�`T�L���?XĻ=��p$�Kٕ�}p���6�=˯�������4�h��Jx�'?H�=�q�5�%ΐ�)5�HF�з��|�@���L������"��p��^+��U��@[]ƙ%�Ot(1��Hz;�x_l�#R�m5x\"���(���X��Y��y"�3ۀ���/6.�����5�I�u�h��!�)^��ڙ��!R���ys� Z���]�xң1�:�,�CH� נ"��q�K��T��
��!{�L6C�����69�~���^����+��.��?�e����tTϐq[C�m�3}��vβzʐߏ}z� g�^=��r���I)S��鬮,D)��Y�)-{ʌ�~��1B��:��t��Zޖ���{.��ݱ�11|�X�6
tO��@�_��ۯ@�r�kИ�s��/���!:� T+b'����_�whs�}�!h��R����$?h�{eR�b4�Fd'�����r�C`/hМ"�v�%ғ�
�:���m?��d��&�`���%a?�}�Un�9�o����߉?r9i.����m�\qρx�:�VM߾I� :}]x,�ZV�H;�e��,����X n�
.��ͼGH~�-�k��y��*}��k{�i��ˮ�AJ)p\��7��[����Ҥ��� ��N���Ӆ��y:���[�m�wCX]���B��.�=#��͢��J|��Қ!Y�^���&\�k
��-��X^BZ��+(�`�m�E;��G�
��c��S����I��FDۓ���z��;�0��_���.O�Z;#���9�5�0I"|��|�b������8�lޢE)��r/�7�|b�o����,y����3�b�f��q�' 9���i���y	��XKc����(^�#���y���&��|h�X(��q���	�/X��(:S� �<+m*<h�?n�Z�����r�7�a�]XN��t�EC�2�@O�����֤�?����<l`�t�=v�}�����e��)��F������p#\����ܮYQt��Z`�`�m~��ψy��Rz����S�к����.f�7
�Q+� �
�Ƨ*��ð���^0n�pJw0��e+���	�M�&�;�\�Ε�ܒ�y;���^�_��:=�K�#@��<����)h���i�r
o�~�C�6ϩ��`x��(}F���@l�e�eq*j)����h�yk��)%l�͓�}��t6�<�Y]
�nZ-��}�Y-�i�6FQy�X�����8vmq�&��v��8e����`��.$�����.&��ZM3(��a�C�>9Ȑ��E2H.7����L��#������`�_�)���m{��pw����p��;����V
��T�5���}�C~B�,��&`)������S���v���T(���sN\Q}k�@e����Ǐ��̑g�vԱ8��QtF�#�H�`��n&�g�:���pG�ԑk��͋��zR͝�T��7�N���W�vAB�?��-��H�Tjq.�Lϼ��_߹��6�"����oA�lx�]4�H"9Y[c�}�c��ボ�P�h���2r�h�����M�׽ǅC�����q��/�fzV���GS��Hۈ?���9>c�u�*�y�@4`��~X-5���f���8�w���Ķ�vL�k�OA�w�f9<;��+{�m,�� q9���'-\�۴�1w�T�NtGߜ�@���=�;��ifpϿ=��s�����^	D�S�a'33C/3���F��,%*��^ƚ�%�Q���[��K{�fI�'�ؙ�^!�[3�T]O�@%�F��%;ٝ���)���"���냞��]A��w>jU��N���v��~vI���L�،������Tg�7�����#+SP�Vd�:�=0wL,�̬Q]��;�50���d�p��H#-�������R�ک]�RZ�.jf.�H$鱱>��-A��G|m���Z�;�-:Cf���%�np5�3@��jA;����oO�m�*NgY�(�F�^
�9�����s�$�
�#e[�?��Ra���Y<vsB�L�}��W^F(I����?�%E���D4��,y����SV��?���\q���'�� ���e��v��@2|d"�p�ccS������zjjj�,��K%W��k7�Ϗ��ֳ����2۞��u�D0*Jl]x߂��ơt1� ��ڟVې�-��7�������?��ܨ2�4�ɋ��hd�̋N9.S-�nr!�ӹ-i����i:)%�	ʰ���M�
y�lݼ<:�<P!���ڗE�~g�O�k]FM��dۨrq;��gZ�F)��
���ڲ#��}cv�s�N�XǤ^��ɥ0�'(��(�����JY*ju-r?�U������I|�]��"9Sxc̐%Y�����
�rI���'Jto#�n<o.��y8O���b��}%�X�����$0��߫,Gb����
q��c�I=���`*tO��&�	�X��K�ֻ�a�{�u��Tc[X� ��m�G�S��n_l��_a�$�V>�.se)ӊ,�6/��ՉX#�u_�_W�q{��pf�zƚ̊r�ԟ�=��>�9��y�3=}��t7ͣS
�'����"�L���w�pb���UɅ\��Dכ��(ăD��k
�k��-D �_�YG�:��4L�����l�ۯ���]�e�;��Uz�S����'+�!b_�ԭ+P�{pY=W�j�ꖮ�������R[��tO��7vJ�ͭO�$����^�u.�3?^:�mě)[?�>������$�o|g˽ݒ=���j0P���q��
��4;n#~�h%���2([�Zw�w�G�����^�K�R�%:t��gW�4���O��O}MMf���-X���YE����%ڬ�J��;�=\[n<Y�
�1���<���-wp7ï����K�=xw�s0E���G��[�_�ty@�5�{[2��M륀�}Ѷp����K�@�����fU�].���]/%��RK%��N44�ͅw�sv6��[��C�>��BݼׅL����������;)Pi55�$k#���I.�&�wY.�=�� ^Y\�K: �\�u�
O�lƾ��ܝ�|�C>��4���j����Xo�	t�<f`wC�m*�� z�7;ڻ��2�D���)��`6O�R�L�*j������8M�����u���ڲ_}�V�\�?q�{ӗ�M�V��J�J�t�5�4/��E-�mEJ�X�<��|�ŭ�j�"L� w?�rH+��s��[W�=��38._?#9oI���a
9�s�j�k�Η�!�g�{F�f?�O�����>�́��
�ܷ�|*&C�� <0�Y�˹ŗ�~��\�{����*�/�ᶃ��?�l�;Ky�8B�i6��i'�~<'����_�{P�'���t��%������S<��'~��ƨ���w�+�S�mCI�M�o� �����R���m*Sp����@Mf�h��kAE�.��� ҄`�AAP��K﨔 !eW#iJD�F��"UzU�5���~_��yo޼;���3��9�w~����c�uxߡ����ޡ����{�@���j�,G6_A�}H��\�8x�T�ǰ�G�umn?�8�ʽ�Xy<�5�߶RZ��Ri|k�����BV�]\�0&
�#pi�/���|?Dq�b�/��H`J���j3*� G�]�q��0��Y�
��5F�ֆ��:��W@�Z����[����""���H\�Y�T��H�`������t�6&4\�u�3�3b ��z奋�l�g8t�~�{C�V'
 ��m�O'C����t��J�nYS����] ^"�q)�4�H~ e�@ޡI�+�� E*BY��,�D��	W�;����1���]Ǭ�w���F����ڿ�?���m0(�-�C!�bh�X�t�2� r�5EYa ��ß�,K�����`�+����� �"�ҨT�Y�X��c�Ӷ�;�����,t��i��C����޳`��!��w��iJ�H�n���yx�[����C�@�n�>����g�|t�b��D\�^�I=�d
�Ko �PT\�
(0+NQ�1f7L�QF`��D�R���޷A�ؾ���a���?��!�8�u[2MX�T2s���d���`����D��%%��5k!�M�Ï sM�z}FR��̕��eǵ|��C��i��ل��(�W=f9�:�U�) ��V��^>^Ul�V�8_�[>b�hY)���C$�2o|���|t;\�W��t�\'�qb�Z
��w���P�� ��-�h���Z��R���t��Y	Oˌ��9���d>=�˹�"G0�����7�c�\}K,M������*̽Q�R8��v�EE{�Z�Fnk�)���ݼ�S�gH�S���&ӝŚ�^�n�v�����CX�|�N��A���*q�����*�Jj��^R{�čY��㍟�f�m���n\�?��y�(�d��Q�i�g��i�9��;��=ʍ�j���Ȟ Y�y	���qz�,$sH"�x�)��ܷǩF2�A؊�j�v�E���e�CD;���某�h%�vr��F7�ފ=G���&zO�����|�V�(E��1��*�`�[6��>��a���^a)�E�y�g��K��)������.�^�l�*���Z���䌛���������ʒ��3|�+�>oo������w������%�N$5�$��]�L ��E���-
%�*�S��� ׉6�OÇs��YB���Uѳ�-��'��A9|��KZ�Z�׿u��]�
%�7�������9J���[�zv<��	S�Ǆ�ߣ��ĘAN1�[��̨��A��\ۙ�������*�w7I��~wj鶙�E�fnoظ�X������XǯVә��u�U������f�����^�S~�4��O@�H��7W�#PM6�J��^@�k�N�Ǝ���,G�Z<�?��=v�~F�{����Qk�n�{lw�mxU�g�\?ˏ���۝�NZOK���S�;�`�b,܂/�q!d���Y�4-���$�ob����b�63V��K��{�փ&C	$ww�������s2�Z� �}l?B��?�n�=lZ��F��r%;?@o����[̰q3k����@���V�|Sr� :��5Q��@�#P���D*'���m�ƾ�)e�b^�wj	ZE���B�6�8���פK�9���R#v� �����cK���[�f/��>"���L����z-��#gn�6)8B�8��2D<����X�����~9h��;�d9�Ŷ��<�x`sʵ]n��f`1ҪL����\.V�YI0�w�]h�k9���i�A��3�ٽ8@�c7>��oח+���H Ԑ�aO���Kf��)�k5�$û���V�egb���y(DX32pTw�a�܅-N���o�J�<��ݐ06y��
��}1�v$�o�&Y��+�;�Ln��p��Ţ!3	Q���3M8֡1��b�Ӑ�J�i�B��g��ѻ_������{����m�t��XG���]��th�Y���&��k� ��҇�O�K����{<a�L��۟'�¼�S�ma��e�5D���]\�?}��z�`d�֭!r�q{�/�+A� 	@ (b������SD��cT�+A5R�w$��ڼ-���"7��ɱ��<��(&�>�?O����T5B�膎P�;� 1����#@��[Q�4{��Zh����C�mf�_��_�=.���2�(Y������~���/M����q���C�6o���ţ
I� �]�=�	zy�Rѩ((;Ϧ���w�o���p�{���u�\�\\���M�0�j����#3Y����.���[Y��u�u@�ƕ^��A���I�#�S���D�l��ǧ�PG?u1Ì���c�[Ua�2�����������Zr9��!��Q�u:\o@�,�s�>�ƴ@�_�0<R�v>��Ḷ�)���ńK�:�y�xs�H���v׀�W� �C]�K�%�dm3cg�ou�(<�_���,���PBaᅭ�H">�X�#ʧ�lQ��j@$��hc�rv�=-"���g��t��IDy��s\n���` �M=f?���F9gsDMa��ݵ�9�8_C|����l��'�9�pn���+���+��)J�:��ryO�1GIXUл`�QH�5F�&P�T��>`"
d(�u��A��#�,Z�}��m�:���i~U)���?<$x+6���~��ԘG�q��b(��*��KhmzX�<Uz?�S%�(���r<�v�k�=?�i��=�T�����V�����O�d%��HL8*=���� 9hy��+�0^�X��M%_~�G;��.^Ґ���?y�VKy��@zL�xL_^�cw!k�A��Ϙ]z����&���]�K�[5W�uc�ki���C�<����y�����X�NEi�#�.j��|���v���V���Mʏ*��f������wt��`���Z��^cT���Q�����S�Ǽ$vl9���E�g��#Ϩm˶�\86�z�=�D��X0OM�̀R{���{%��U���-c�8i����L΃��JSӂq-���h)pM֦�ƿ���M�oms�;+|��X�a����'��hxgQ�\9�]�� 'TʼS�d`�����7�;��*�3g�.4KN�<��p�Ja�RHF�?�6�7U7vV�������mSbV�V*�㇃��OOM�h�� ��"/�Cg[*�}���=w�\;���B�uJGuYC�	��Zh�Q-_��q�������"m?j�o�Ցjm��ӝ?��㾋V� ] l;�1��
7[3�I
TKk%N��Fn�X����G��脝{0�U �R@�矸~�.7���lՓS���K�ns������*lpoO͑�Z����G���Tk�AM�&{��v���M3p��Å�ǂZ���v��+��WF��震4�	z�� �A���
��ng܃��P��ҍ�٥q��<_R��>%�ր��$�(�$��p9?ɯ�����-r��3�`�JQ5R<듩���	0����A��Q��^��r����&��U0���!Ӑ<��������|�Q�������旹�>�j(1��+K�~���<��K~��SO���p���/f�����I8�����͡�"����; �:[�]yX�������9K�q
x��u뎨�9�P ����[@��n�Y�@�P��q�KRpQ����%����z_' �#�~�Ti& �����M���Zz��L6��?O+C��mG�g��TB	��8��}Ѭ�.��ƾ5�յ�$�/���)���������ު���dzoΡٲ�i����Z�Rv_�����эDT�}	�%#tyVcA�,x���ٍ	��<��0��(�pz��L����d�b�B��'?��F��Ò��ҭ��׍���s�7&S�C�ƀ�0��z&�4��cGδ �������ߒ>���Һ)�<���������q����U��$�����圷>ǩ+qK���um�;#��K	���?�zN�b�|�Xn���QrW��ax*�ކ`�p��.��Yn_���%�|UeU�ij̵E�(8=N���q�Co��u����J|S�I���L�����7b�B�4��v���D:)gy%�js�m���29]�@��U�x�鯅�����k�LzƷ��{*�9C�s�k�[ ����Ť��n�s�վ��<�{��*��򍛤���uu����9��& �nuЬ��|$�_ l5��c"]���ZT����:6��4e��M�+u�!p!y兖�ܦ#��O�{��Amt��*�yQ{In����@�^�4JN��,�T����ު�j���Z�� џ��q�DZ���+�)��"�v}XyD[g���]!�v���7r0����Cܭ�"��;�ծf>��P5 �O9��R��M��G�s��pY�>My�gL0���ƷS[�q�H�Є�,P�\mT�7w�C�E��:�`EBr;��a��N_�|��,�9ReI�Z���I�Ifn<F���.7�I�ۧcꮛ�3۬�̫�T3�C��P,���ؕYt��᚛x�T�J'�lW���tv����ZE3{˽��Ty�	���,��M�n�k���l9\'g#�gJ�.ׅim�`�+�A�z߱�^Nu�Yz9$��Pw�M�b�w�d�ne�T#�m,���:��-�	(�ʚЎF��]��H/�i����@>c׆�ޟK�Zz\vm���3t�o�E��Ƌ�z]��C)�F�,:�Ұ���~���q��	��T�ۆ�j�ə�E�ȝU���)Xh��v#W��!m�wb��E�<'�DQi�o���+CCI�=�B�Л�&U�i:�2x�\Y"DA(z�Nf�$u�	ښ	��������: �l�Q�<ڞ�\3��0�|~����ZռY����ɍ���VT�ϵ�~~�Ck���K������=�7��&�`�E�3C(k;
 ���=����3���+r�m�T��]�3`�tj�������~^��̷���y7xMZi;�+�C�eA�W��i����r{�#I\}X��{ɜԇ�X� �G���c��}DV����Da����6�^�a溺*��o���Ǥ*�tv��9J�͗�f���e���«�	lM�.���u�آ6�[6jༀW���RSX���[&ݚU�dA�uBɥ$<�
��2���V�����$��|0y��j��
���.lZ&�I��[z��<�fO˙z�[}�I9�ܳo���'�w�'��Öc�����m�t;ס3C����i͖r��΢2]D���!P�	�����o�Ik���B�ˊ#��߲
g�7�r��Q"�՜'����4/rڋ�����4�
xx�RZm7�6���]�p��I�7w�6�rO�#��[�ZC\<�[��bs�@��,o�`=|��B�~�
Ji�Ra�@�܄�w�zf�,x��k�ly\+���o�ʨ��>W�^D���������7ŵ۫8ԅ�r-�bl����b��uE�z�9�F3��c�[���p�t{|e�}/��E�HIϳ�)I��ߞ+{��۝�IY8z��w�`���7Pi#���ћ�]q����fX���'�~��eRnW��b��2��@�U�{{�#ZBT��ـ�􄀨{~2:��uq{!$��h:���D5��6"�,�T��T�]�OO��X�F5&����yc$�����}�[W&f<~��+?W�?��K¸�n�����B�}��O��k�.כu�%��ĸ�?_E:�;�(�� �/����2����N�J�)^�6�/����F�Kwr���Q���*G6�����Q��g�dE gf��l�X�j������sm��)����n��_Vؽ��^e��p���>9�J���s�����gs��`���&�`lS����/�8�mV�b��_c�E�xd��Mgg@�@**�����;	��_����"z�V�h	�
��9�ă��;�T"0[xי	�����Aw?�g>bT���~��/�}~����;߱wˁf�\oSS��_�zU��� /�@>��יc�C���H�U�kB�^co�<�AE�Y��'�Λ��,�z�ri�H������C�6/���D�̻?��_1�F�dz�-,� ��P��*��������M���c�^K���L���^6 T-um�JF�F�w�}�4oI�����u��b�����h��ӡ��]vlMU�vou'����2����rY =uLa�戄q���W��������!�(H(�<���A�GB;b�� ����	�)�'�c�7�����)�����&����6�6�	�x>���^�؟ն��sH������E��]&� �����y��=��;�5��_��d^�N�ߎ�_�8Y�1���#�j�i��/S ?+Ӿ���&�⮖JΒH�,��T
�����?�C;_�(��,��B51�����h񸊘�c�nr��<�O&ƭ	��3�J*�� �E����-���zYP�ԋv�m�N'�tr�L�-��<j��n��v���$�mz���0V{f��k	D�-�m��c����E�B �:Ɍ�7��K'���KC!&#������?�d����AЇ�3`�~"��h/���*r����z1�1�TWo�hj��g�t���(pg5�p�bY�7��խ|<!�E����jb��j1��;zbt�&��"r�3|�33EBoݺLZ6*���gl@�&�g�i�{�V�#�s���`��N�u.q�Y��2C��S� �*�g�s{^02:;�h&�`k�/�r��'���#�>�2�#e�;��w"�s�Y�� d�2�`3�q8c�@U7�y@3py��8�$˭��h�!�A�Q�S�-7~�I�}�����B�B�}�����\J�����%ʻ�)�y����E9�&�{���p���ĵ�c��� s3�c�p�Á��q���R�R9c�Z�����+�
�vQt@�'u��$�B_Q��2O�h��ԟf�ɞ���z��W7�h��~�����j?��H�d���m����!�J="��Z�� :)0���7�l;�0��@�
�p�e�_ ȟ(I$�{]jmrI�M��L"\�Ǉ\��3v* ?vy"9�=Ma�y�������c�e�D~KcG��#f/P+�^H�h� �_ڼ�O����p��b��!�m�<x�+���un��fG��ˋ�7�-��X~�hc1هB���~���.���E��c�p��f��9��^���Xu�:3�E
pF�{��p�ߥ�YA"�����.��uk���-[SGZ�6��3�h�*��������6�WbX %� ���[l��-�&Z���QZ.3�`�iUN���w�I�^��X�X���|w���AE�s�K���i�3�K��k��d��K�J���bKH���c/���W�
'߇������쟇BM���y�πެ�r�5�X���	�:��2������?D��ʕ�*��5R݉��Y �F�}��7gLj?�$�\^��4�)��9d�w[_b`s ��~aRk��(�|��S�%�0s6������C�;�t��������|Mh��B�-7Px��C�vY�@\ה($��J�e[��S)����~R廨ʧ�"���]�c	������'S�F��H���7N���G�x��Esk-��![�|�Y�8�n)hTY���{>�ak4��G�`�)���F&�l^NW|�S�J��> �%1$l=I�M�h\��ˈM�a���
��S�B@�PgC)��Nd����-I8㼔��D�:�v��Er��V��-_�h�V ����﬘�%��@��ڨ([r�p6�5�mr���MR�����R������sz^!#U�������`��a�~�XV��T'�`yz��G���^�
�j';:��8�=S�o,E�r��-̔:�������<��'�]���&���b�,Ԃ%W�+h�U#)��cf��V#Z|<�t�Ư������Ϭ'���+)p�4/l롻��j������c��W7V��Qo��ۢF�c�2r�`Q�/�f���L�s��r�q����~�h2LVUY	K�j�f�Ne�ƚ ���zFi�o�zV�N^?�+�$���J䴾B�^G;�0��t��T@A?{�9�� 쿸X��>�Rl��Z��4+ǿ6{]��pD����'d�.�5���3ڱ�j}|�\��n�ys�8v��V�� Z��8���e&���pp�Em���'��_�A�+�c�NO�F�Tȍ����*&G�����C�頾QN�	+z��--��F'���D��7M�v��6^Cz�Wl<��Z*���8m�O��y�K�g/���
�?�S7{� y�;#�Ժ׸�p⁨��_����O��{�,�S/�5{��8j-O��5��ӡ1�^��P��;ݍ��g��>�1}��1��J�Xt�7`?�x�o����4FD�qg�	�O=��i���`?a�QV�y_|QC�Eջ�Vv�u�^P�鹲z7Crd�2���񈪛�}���w�y���� (��60��[`m�yW�������ms�ػ��4�~I-��=���3x��*<1�٬P�n"Ǡ�ݳ��%[nW7	-����l(�a�t��,�H��V��35%�EàFa����..�vD��Q�I�LKn����"�}'����T����f ��0��%�>�oz[Ɨ���\����j������g4m�Q#�&g��f�L��)-[��d@$,_��z{D�J��v	`����{�����Ȗ��� xY��f"͝�6K$�\D���u5c�f}	�P:�mQ��Z�j6�_30�ӡ∕�u��TZ�ַT����
P��ע��%Vq�����߱������[��
*�����=�3�R��NK�}�^�h��W� �]��m^ќ?���Z����\�V�R�Z�s�-��!��l�X>(Lֱ8�DLDc�T�P�.�a�<�f��INn�!�D_�l�[��[ AU��|����Pn/�:���H�����/�N�#;�E��F�d��|	�@�����h��Z2K�^��T���R4�Y	n���]/�?���r`��[��<��Ht�q6��o���%	�^�2cj��捈�+y ��*1�,��Ъe�V(�K��j����&Y�T��B�8ȧ0ק&�[�Z\p^PQD�9��Ŗ�M���/�lz9�v ���L�<�t��#�LI�B��5���!T��t*�BڹR�R���#�h��kZ��k��#OK�yN��Y A��/{��� �S�X���)�ﹷ��ܬ�o*���"Of ��k���
�6�n��8}Iy�(�^����C��D�;<�>��I^@��i`���$�5���OxnL�z
H��o12��� �&B��c��Vf�9��{V�T�w�^-A8y���^���8�բ��ia�
��������Xօnw�]L�t��Mj�U����8�G��r�bX'>�������7�q ������I3gE*4�M�2;w�U�uC�y���}���3��qy�Z����&�Iݮ8��]4Xx$J�l���S�Z^�q��I�^&�6J��ή��Y��L������i%i�����AX���8o
����`h�ZE0�+wT���a^�뫿�~a��J���Rﳡn��_ݨ%� HJG���t�s�l��#sM��A�u�0)K�X��6��´�aw��'�)����s�s_s� ��~:�M�4+V��?�������-��Ϣ.#;��d���(�к�Z� ��wqL�}e/o��/!ǡ����~/%���H��a+��o
�Do�-B�k�$�y�_���C?"��o&��ڔ/���_���Po��b�6�� ��};!S�ũϹ̫�hk&h�~��PZ��#��"+D�&x&� � HQ��3-r`ޫX���W�$��yƉ�&��d�p�u��IH��Rϗ�h	F�\���s4�J�}��'03��@1d����|���|ݬhv��#8'��
��(�}���P(9*�>P��`\�z&� �w}e�:3.��X��5�K�X�{*�C�{�x�N�W-FMF��o.{��V���L�N�U�XoJ��U+�qG�ndx\JK�V����H�ܿ��6� ~ ����t���3~�;�B���J]^S���55�5%�޹��*l��U�"��^��z�Z�tא�CݨEՆ�F��8Y]\�pk>��~�����F�9Oe]����ɹL0�x�ܧ�U(@�@�.g�]�-X�@
�:P�E�����?sq�m{E{f~Gm�_���3/�:8�k4�S�N�_{��ZJ��z@	��TX�-��h�\r�7e(`c,![�������H�78�Aί�p��{:�s�>�5���0$����w��}'�Ԥu�\!_M�j5&��!� ϱ7R�s����0��ot����]�֣�\��p"��� �'�D�Ng>Qԧ'�~l�6�B���﵂龜mA��h��k�2�Ǚ��jQ����a<s�Ũ��&�H���������W����3�ȍ�E������[	y�)���~t��s�l��l�]-,xSQp�ި~9; �++�m۫p�G ���y�m�#�Q�HHP�i�d	Q(�n(�EЏ�OD6$F�E����~���R�s�I���J�z̀���ڐ��1R��lK.�{F.���Ԕ���6鲊�?GZ6fƧ4[їU�_*%o��4��U�H^ڥ�z5�MC��}�;1���ŚM��:!��ͩF�yK�c�d��-��R_U0����2~�Q@k�#<��}�fSMUHxs�1=Dx�e_r��lQ���K�ƢBBl��ф�)�$���,��/�J�FW�^6������W���`[`�&u=W�\6�&�Qpx*�Ulr25Y��I@��I�������t6G踒K��h�yqP�j�]�	�]�3��.z��+^���J��{�Ho�?]̃�b�+v�\V"Mݜ��ѴT�N�lv�� �dx��YaL�M~8�Jw~��G�̍VL���r*�M��r�6�,��d��M5�q�L�M�c��3��@9[b4рz!Ea�-���W��}`���Qf����Ⱥ��x�?���E~��u���˸���c���C6��Ja��^�	�J��۞�?|�w������9����&�N�[PEJ��7P�0���Y�[���o��d���0����g(+�h���_΍��(�dA�F��7�}C�n�GY�9dEəEr(�s���r���6Vr�K}�mF��wg��kL2�<B���Go�
�J�̕��وn���Vq0�r�ne-�Kz_��m�g��愝|u�KF��kAV�m�\��YV�B*܎re5˶�%߳�V�4J��Q��Τ�+9���6K��Y�͒��o��L�m���y�M�MY��AnE�D�k��w<�k�-Ϛ��n�V�׮�NvK�jx�Je�$���W0��}탵ɡ+D�;~��v��,~���Gv�A�S�(�	�iw��G�U����
�z�`�!�g����1(^Y�\�u�a*���]dV��p�=[x0/�W�RY�gnL�<��^�M��)�ӛ7i��V}.�!�a5���}�lS�;��)} -]R��~Gyˋ|��R� �y~�p�}}3,zʘ��t��r��DE�
r�ס�9�P��m�䇅G�zj`+9Td�?�Å�غ�5�6���ԕy��f�viPS�4�}�`��E��R�Ej��<��\�e��l���)�J�}���R�`��K� ^������jecl�8�2'	|�B�)��s� �n6�h��~*��콚zl��G�X-#�������������,��C�;�ġ=���'1dMqna���Y��3�s�t�O���w^��x�����Y�<#v,�%��s��WL��J�j�z��j׆/�Sfр)<
�7@N�������ZHҞߎ}fv��NRv#*�F I�0M�g�J���\E���2��Eg�2������sOȇ�+H�ý���S]�؝����6��Q-h�N�BҌ�������I�M0~�a�s��^2Z�(�W��t���J�m�r���fQnj~v�׸�ӵb^���TOSQ��Dt� ����m)In��t��s,p:{jO���l�5���̳�L�޴]�ö�M�v�>(��K�z"
�U��{Q|���e��H�����_�����d�?�d�e)�ܢ��)ɣ��b���]snv���h<���4fR���uj�����8}7I�g��*i"D�H��?�ɕ)���3=���lh�e;Cu��4m�H�r<����ƀ��#��S��'��T���C�mc�|Co�3n�$�sw��.��k#��x<.��h��e�φ�^���+w�õ,����cW��5mJ�i��Jxݓ�ya��w~om�jl��|q�CG>fn�I��t������K׏�%��*�M��X$ұe��G��oW�3����Ty<����~�5J���q���1�?i�T�AUE!tJ�k�ude���$.��;����q3����vQ^ �'E��Ez��&��N�&�rm!m����5v V��	�)��5Ɠ����?Q#�;�^�x,�<$���E�e��a3G4p��<꣋~4�
�z�k�sf:y��YL�ԈCg�d���#0��My�i��t��F���k�Q�N��"�tc��N�+�P�i�w�@EѽU�c����W�N�J��zg�%�&�{�'�� ^ަ��-��Eŝ��-�KTU����6s�G#mx��2 ai���Q7��[{#T�G�KtYt���iojx�N���y�?(O}�w���/�1�1�I��W�ѯ�Z�i������,Ĳ7
�W��>��߈�|��LR�����>�
]��c��ΩZ�HSR����BwS?�O��S�ّ��!,pт']�x�!,�#�D����}+i~Y��Βq�N�&P��Q�׎��� u�ٗ�)��?�~����@/�(M�/�u�v�Tv�?T�<BW�"�c�7s��1���(��G�y������o�+Kr�/>��KwG��(}� h�X��H_z������T$��7�X^�xޥڮOw5�t�����,]�T1ѡ����-�-TY�� ~h�,��Ѥـ�,�A\n�1�2�~@�*��%�P�Ł���\�pzij�7����Mu���u�<�pf�f�v.���
q:
:/Q�ȁH�E����s�e
H���8����3M} �L2uk�6ߍ��H��H)n7p��f�w�����.Nii�ﲙ{���g�8���%��3K5�x��Cm�K/]Q��@��J�:��!z�ӄ��G�(NS����^u��0� i��@�SZ��R/�s�
���7��|���h���M�߰�
�ǟ�^&u����N�@�0=��ӷ�;lǙ��PM���_ʩ�]���Q�!QQj���v*��Q@�eTqD��8l�*g������h��l@���x���5zᡧU8I�%G��:�w�GLN�ݖ)��T�E�Rj_��|���c�3O��MNǟ+��~��|0�@����D�0D#�)K���V���fX�S0L��Vv��KU�e"�/vQ�8w��KV�Έ��&�L�?�Gb���3-��]�Q�g;�KL��q�(�(�i����ڞ�������Y��29����û��A �������Ϭ��7A�&u�oѼ�GLa����������ߑyձ�A�y�)릏�8ʒO�J�Q�Ǝ�] �����թ!B���}M�]��^ZI:�=@O�3�)/g��M�����`4,Y��lӨt�nBc�����C�����?���0�s�}r/aS�� \��	j����Lw()
�߬��e�ţ�
�N���\����d_����wg���pI���(S<"�9�{R����X6�WR��	˼hO�sh1��4�G�U��M���3D��98vZ�r���<u��2N�HWx��"i���4�y�c
�_qَN���������;���T�z�F��q�(f���d������Oe��	�L_��/�Vy�w�vH�歯o�^�s��֦�å#ػ4y�I*���ӾT)|S��cK7�e�R�ڎ��9����O��\�b��&7���E�Y|���w f��z<�tn�0���AN�hǠ�� �=U�MRfɧ�EEMA*��rIz�å�ٵ�T_�*PU�T�m��zk;(��+��.[�A���e��O-����U�ӳ'�O�������j�pݕ����*�u�m��lC<mB�A��xe�$�C�aMܸ�3��U�ܟ�)�>�so���?�'X�V�+��Z%qM���s��lu����0Ov�����
���y6/g2�o�U�hqE��s�¢I��� �:���Ն4�R&�\O�N��3�yD>�jV-g��6L�|����5$���(3������~H�]�L\�\����w������LIIab_���s�_M�_��ܗ���������A�DW���OiEΜ��'��u���hq(Z����{�������Wqs�[]��g��_H�x��:j{�Ez�5!�6��Rԯ�<ˠwu�֥��h5iL�h��gJ�^k�U�O�oH�P�4!SE��)��w�>�n�� ��#^���@,O[�?G�'>��P�-�1ku��6��&lB�%�E!LJ�����Pa�Q�?�?��:�-���7<�7�R��f�E��d��.�}~Mj���U�P{=;Z3� {$�ͤ�܁���X-7��Wm(��0ZS�r6�n�CkȪ�2R?S�f�4?O� ��_$�����a��3�zz�㐇'L�8���EБ	�`�e3�� J��+W�����6M�ڳ�����k�N��|��Fs�^D����"��C".��q��Ϟ�q�ʞ9������\��=�E	�g[�
�����]_�V$��eѿ}i!��:7K��Xj$��qB�R�:�[����O��فKUß1�Sm����MYp�J��p�l j�����܊�É�Mz�X�Զ5�~��D�e g_�u�������N��P'����k8`���?��z����?sAd����B}�xl�.{KD��^�\��"%ʒ3�|%�YӠ���bKJ93$��OV� ������nkɿ�r��fy4�N���R�~����pIW���c&�7�
�곡�<|3ca~�PM�
�nz��(Aw�G�ߪZh	A	#�f_��B	�xh�W��r�a�������^�r�/�Lyp����&��?F�迿�Yݮ%�Z ��Nqm�tQ�#���'�~g��Dֲ���uS���ك?V~�  �?�3��U������/�w���������9i�G<��z�ո�y̓�~��c�#�^��_���i�-� �"�8�<Z����ܾ�����2���v�)�}��=�#7s���ȸ���Ť�il?l���]�� �r�wa��7}xo���* *.��s�N)���v��W�p��$�����/�r������M��NK���ߙ�JW����Ɨ֖S��ca�r���Nq*	 �K�
��e��
N0����Q��6�&$�.� C����k������O�·���Rƹ��K�����)QՖwէS<�K�k�ʛR
�v�J���9r�!��E��V��I�|�@"�ن�1�wBz�.xhG��dZ���cW�e rO7Q<�x_�F��I��Ley��@0(⦚�˗A���Z����ڏ�?|:f!�����G���'l.���9a(1�G��x�J�q��L��5�!�P� �ͲNH���ف��1�?}�񡱿	k����6*ª�)��o�S d�LL����fi}���]�K�@��4>����B\��M���(��y�D�gmB@��<�2̡[��U��*��`���ǳ�xo���o��FZTF�;N�����6O��e;;���� ��5VdI�s�r�Q) �	������T$Rk�߾�cC���0��"_�g!rA�;��A"�o6W��=�#Cc��JR���ykW��B�/��G���R:��w||�W��U�˷�E�'7;�/D����rz��`�߄�C��vf�b��ݥ�&ߩg�J�B��v��]�L�&�1bv`��/jք<�4}��pqc��T�)I�l������^u�$�r��ed�`�,����:vzW�I�Н>�W/_%6�"Щ+�ا�v�1�;oW����e
����A�RC�x�d���v@g=�j{��=v:`}�Az[ڗO�~i������3 �m�nH����W��Eq6N.s��,����-�iƋ�+��~�D�!��F�c��>��@AN���$��66��UT�8���ͬN�'���Ҏ� �(�vִ��.���? ���|p��/��a�ۦ��YY`2)���/�	5ɝ� f�������ӿ�����"�mZ�
�ޏ�.eK@IE��d�ľ��rY��^�i����]=���^c������ǰ
.�v���F.��p#�����gt������9��7l�NO�[��e~؅nHm�13��)�@��M=�S��m}������$U��R�Y��b@Oj�ڙ����~�;��q� �u~68�������i�o����oܻ������ܛ.@�ӌo
�\[Q�Q�JXٛ�^й�%�G�l
N1a׮C6v8�i����y�|�������E���E�|�F�EF/��7�<��ow�Q���t��!g�"�o㲿P��4�>t��u 5L|\��!�m�*v�	�O� I���Y+A��+Qr���e;+q��k��Mk��$(��o(d2�� �A�f�ٮQ�g�
]t~���b�§�]0���WE�߱�Q�<A�E����.� �Nvq���` |��������##����@�A�6%1 t �������'w���	� �@�VD���y�R=�H���K�=&�;�^�n�.�S_��%���{�y3�+ʘ|T�#���-0na}���~�-@wF�	�L|� ��M���2l���:5�]�W�e��K��}�C��Cru`$���z:������~
�=/�)��r2��2��x�h�t�;� ���x��5�*��\�Ose�$���Ǟ�� �<�sbqG�	F�ɕ,~��\N:�w�3�	�;���;���|x����/��o^*��f��V��N�Ƙ���	 ��	{J�j�SH��Oȧ�m�{����Z�c�xJ��O�_Ew��쫡�Ɔc�/^�}�����ӵߛ�Uq�:C.3�����A�\�ځ����*q�lU����$죈�������L�>�Ǹ�`˾�2�R�De�-k��8wz�8ƀ�V�l*�͏ ;�Pv��I���}�rSX�KoW��P���Kc��[�n��@S��}��'��`T��Ӯ�X�2XY���ad�{��F�� n����K^"~�b��j�/rۼ��\&4n,J��؍{{.]+{Љ ��o랴���%ȺG��F@+(WY�ӯ%�Ł>�ޞe�э�_e0��C$�C����7��F��~���1d��K�͖�Q�� �!zE�蜝���|�����6b];�]W4����?Gd�� t�-FE�	t��U�r�B���d����l]F�Sb��j���Xp���,+:�!IC.Ȁq�L��~��S��8`j��~� ]WnO&�B#�>��sY:�N>��� �((�н���F\St���EC{kk��	��I�{5��h�Zֳ=:��()��$��ܒc�>������	���'�["�PDc�>H/�����B0G���c{ɜ|��~�c ��4�)ū>M$&?�����/4����2t6�e��>���|���B�e��rf�=wZ�����\��h�b5{�Όww}:��*A�l��`�X�|�j-ɢ�x�nƥ�~��܎����pEA��IF��}{0�� \6�8��A�H*KU�t�`f���E|!;�^F\���/U����Yϛ�:Ƶ&GA���I�TT�΂G�99}>���>�q���k����;k������B�O(t�l}y<������n��n��H�,���5(��}m����WeʖK�*;YʾO�f'������Gx��}<���3����y�g�xfn�*�-i����O�d��d�9t�ŭvB���S7��L�\������m�%˶�*�[�r�̶�JW.p'ik��7���b��������Su�
������G�K� ������ь�ڬ�O�pg/n"]�)X,vj쨍�C��V��8�{x��N��o��>|�a�$�����8tY8R\�W0o$��r��cp�&Msl��_Vh�=�rT�z����2{Ƌ�p��+Z�!��+��RS@�����6�A��7ݐD$�b#����4ǚIn��_�������ۘ�vW�\N����KE��[u�iƏwH���k_M�l�h�a�k�]���TnG��f��+�؎���"뜶�Q�U�����ü t#K��?tˆ|.Qm�[8��s ��+C��VkvUnb�$w��Y��=UA$�[GۀP?��J�
TDٽ����KJ���'�NU괧��iQ����@-p�����I���4#~޳Y>��|e/?��=�aoI�s�.�a?�苾�N-�w���t�;6��s*�����0�W:6d�J��{�:��h|��'�)o�s�H��k��\�|�&�V<�l��/B]y?�Tae���8���0�.��#��؆�O;,NB�������B�;�?�gO�a��N?�n;��`\go���ʒm��s3�5�.K�f���u��m�����lz��5��"��Y7t���p��ħ�Kb�e�Gm(��/}��"�芍t���e����o�~��d�CP �+�8�n,K80j���n�o�tz��T4�����̹l2�+�➞�|�{�g�&)�q���a��v�d�a���D/ǿ��G
�f̷�I�f����ݪ��Py���������w��|����:������:�rfT�����?|,u������쩺?I���@0Z4���"
�iQ� �tC�i[���Z�1x�� M�捙L>݀�t`�^�lL���*$
�.
�W-�6��Yoa֙Y��EZ%[Xr=�̣�;l���΍�X�b
ȃ;�-	�_�oԎ�?��]�Bq :�����6l��̥�I^ݦ�K�J-%D��m4PB7�[��O����x�>0>s�ze�L�F]��&�$�䓀O6egd�ob!��*� E��b�7	}3�����P(��(e���NC��Ҫ\ƨ���ͭ"�.�¨` ��᠊*���LAy��?-EK$��YC��R�m����^�v�
,�y�$؜�P \RUxUȧ6��b�5�rk�ĸ�B�����;�j�=2[�c+�j��J�a9���D�5��P�}������MA�_BF� y���
i��	�&P�P�pڵi�%t��nhftg=j?݇I��H�� ����ݚгqG䵝ə0F3��մ7
6#W��@~p2_1�EY�6[�1���֮.yn�m��Գ,�����_"������4���e����,o+m��ϥ��kf�71�mL߷��ߛϪb�`!Ty�U_������j�w��n��u��d+yZ�H��	Wu}5}��E���;����X�_�y�j��J��~<�@�?����_��Ɇ��['M�Ic�C��0o��Z�<���f����w/@$I�������o�إ����E��̆D�f�R����;DME^���l���P_Y�?��W��P}��ۺd�Do��x`q;!n����ڄ�KC�o��q�~��)�6�W�pi�� �k�	�(�P��Udppr��U����Fw��:�k�/l�XX���M���_���n�Y�����v �v���a��;��y�-�`ڍȬ��*��[������5N�C|{��A���߸*�n!9Ԍ��`�;�6{}�!ea���ŏ<�8L���U���@��뇫Ng����j]��Q�q3��B� �77�0��#��V.e�@���Ϫ�[xD��'vG�����4;?{N�=���(�e�H�r����G����UzE����me�/��������ќhrǙD,�V(�m[�f
[��o��r�Դ�O0����C�(����6ow��@�yU�:Q�*�)�(;7�ޫ>��31<3#�b$m�3T��)K�����c>�����$���8k���9]�6��mx�;�����#�UT�l��{2J���<�+�ױ�W�/�6��M���|D���(Eo�
��1x-��]�E��K5/�wR�q%E��$��ӆ")C��贴�K+i:q�"�i\��&O�����m�+��/)J���'��+X�Eҿx��k�Fڔ�`����c ��2�R��t4����������$�a�@h�RQ7���Q��۟�y$g�OkK8ľU<_��ZX �0Lp����[R[���ړR3�&�C�'��U�eo�2�:�]��=>���B묬�,�1���Zl��ui��~�6Ȑvg�ٌ��,�"C�C���������
������_I��3�(�K�f O�	�&���W�AŃ؇�6���q���g&�����2��辰�[CB��r�IwxA"|w�֟sfd�Y��v�����aS�3gzk����x������
����F>��/`W&�b������{�Z���p�ܚ�i9ޕ#_��Tg���I �u���܏x6�ȣ,��Bb�3wވ;p <WCS�H~b����݌xR�rj�C���4��]�bM0d_Z�Zfgwr��xǖ-s���£���]@[�ob�'+�;tl�8w$�Z�͎�8�o6����!�z� �+��� ;Y� �A3�Z����q�!���v����ғ�"o�I��Ԋl�_7nؕ��s���	�Kٍ"�*\R]�E�S=̩�;�O�&�V.��b���\|��U���t��g�ݕ��D3^��9�FK�`9�Hڕ���h�L�P�ڷ_<vf�w�9�ʜ�Mqv�F��k������T�Nt1��;<�Pi�����I�Tx����
'�!�M6_���Lq����\sw�*�U�f�'�N���{�Ivk5Jo-|�]�F5��+\ý��T������-7�m�n2`e�(SX�E(8��?ޑ�bN��c���ħ�)f�~�����4Yd�.��~���-󔊷|-��K�*}(���ii�*R�nK�̎Ō�������jt)u]��.;V��0r�*Բ��U�9��t�io����2����v@4���S�M>g���4=�˴�j
���霦A�j/a�A�	y'���	�����	�B�r�5~J%�J���A�j�#�%�yR=`���j�Z��j�Iu/fi%��z�͉(��0A��N(��ve���'�#. =��sٺF�C#\L�}V�a6�xp���i��=ɱ �i���X��&`�lOt��^Xt�m��Y���8�����o?�n�<=(dm�@<���`e�Ӛ�gZ7���	}�ϟs���&�ff���/|N��G�Y�0�5�|q>�ȱ������V��dH7Ӡ8ˤ��-���E� �E%�{'����t���W��g"S�=i|��O�<&��O���ə��_���AD]V�R�����,����Yd���?��ؗ~ �P^+�A��?- �-���7���mM�HS1�@��y^;0�ce������޽4�!!�-��gẰҍ�N�};;B�}	��Q\*�g���W����'��W�a;sx�2�-�P}׍��RNK����C8LS���ꜙb���!��J�� �e��2t2WS�����旁�bsCv�[Z��ȥ�X���ٟ���n�H|!�x�*_�
�]Ö�q�_P�(i�������$,�<"�~/!K��բ�_�_����C�}�\�ۺ9��wT�M�5�����@�W�N��B���=e;p�<�S�0z�,�o�5����bQ�v�|�s�]A�?��U�-�2)��\iѫh�\��N��z�UA벅������瓴M� C���g@?X?ه��~
N�.V��fy�k8���'T8˳���0w�*{�u,~gC�C��w�9s�G
d�
�g�T�d�g9��DG����ò�C���\?�Q=hь��c����0w����Y��z�a�kh<]턾�N�; 6���[��ނt�f0����(����󌤇v1�03[&�]���E��9���Ho҆\���h���V�f˕�����x7)�)��y��u$��ts�Ɨ��FQ�v�6�ً�\o='�̼�/�l��Z
>]ݧn]8|W]b��J&���)�kwp���sK6�6���V�R:Ս�cdT�'����D��6�9Oy`�� �]���%�����Y��N�W�h��ogh�9		���2��Nn�R��O�fQ������kz�Ef"ŷ��Rh�U��K *�d���М�X��#�����j.���7J.�	�k:Z�O'��?h/T'�����S��>.8�8AZYF��,��T@�N猙����h��G���OLd�Ep��N]�A�ҕ��z`KX�;՝2�K�nR�pNhK�E�>��4�	�۸�Ӽ��_9���ci?vO�j׉��z����u� c?�HP%�f�{_�&�!\����̽���9��^Z��O欧9��Q2Ni���W:�9o�OT���s�����wꝫψP�<�M�`�*`�|c�@�n���be6h��9xVV�L\;��r&�n�B�ŅN���g�@��5X�n@��ST��&$���>.��9||^�S�6,�"�[y|5{�s�gƝ��q�Wq4�ͦ��0��T�,�?յ{_־U�)�[*4�����v�e\�H�5Q���߶#&75YCF� K�J�bG)ׁh��Z�,�i:��u
�\
C�*%xP"����iۯ���>��#a���pw�����7y܎XM�h}����=?���uѷ�/�@����5�w� �Շ��dq���~��6?�̛eǽ�g_7ˏ�ׯ���8�^Y�B"S���8^y�4�� +q
�L�X䑜�s)0L�G$W)5���3w< pn��:����gq�-ݳ}䪾�51mr�>�Wc��!��1mS$��`=��������(�V
f&'�k'0ѢT�sj|��|}�"���?�B�v�/[�=	{������6�h���b'wIY��wnI�f�#IX`��i��`���O�X~�ܵ��lF�,��-�3A����8%~����F�~��������I7��`���+�m�j��#�R �t��:��V��Kf��L��3��A�9���Iv�r�_݀�*k�j:���"�J�5�����j#v�F%Kp����؈��Vڽ�Cê��IW�Y��q;P��7���>H�'I�A�~[V
���84��-%i�MTbpL������~��mu�MS�մ�������Gj���8��/l�GZ��S1�g�_Z�4�0�LC�'�o@]¾J��
x�w<�os��!'��?��斖$����NؤFn��ɭ�p�V�@���'nD�oЧ{ߏ�07/8	[��M��0�X�����f���	Yr�h a>l��F8�*.�mw&���-hcC�������;�X��T��pd
����<��\È?�-yݝSg�N��=�`D+����"y�{����ok��7��W��t��m�c���I�|ŷ8��i�R��&**{����I��_yf�6�r��:�ف3�ގ�Q����3i�i0Z�1�L[7�� ��D�;gT"�W
�)���'�}�@A���7n��Gv�1��B�
�F���N���b���_�B�NG5L�C�p娾�5%u����O_��
�����QO-O� �9�����/�^�mf�'����M�M���3��Cg�\d��OX�9��Í��#�����V6�tU�j�����9�T��V3|(�Ǡ�q��Hwg7q&ŧ��D����Q;�+pSgSc��f�}}�⁢�ax4P�,��P�C(��'>�C8�T�$�k��	�F~��@9�4/(��A��8w����7n;�ZB�����z�v�!��Iz�t�Lr?���$H�A�/�|�2��s�F|�Z��Sz��4`Dc�������'��i^_mj��Xs8�/�m�-Q��drZ�XC�9>#5"g-Hq������W(9p�W���z�4����P�9�
n���x���T�%1ZC!�Ձ�/yӗ0�O8�n�}>����1B�ڦ�|�� ���Ž��{�iG�c4��|��FAW���|<�ǹ_u���C����45�Oݗ��LM��}8�A���rQ���0������"\Nr!�k���k�绛��M�*�c��X��䗞�+"�zfeqf2_���bnN�\�tOgh�pM�������J�HB᪷�z���0��9x���`:�k�~݋y�����+k���sx����n�ب�֤�;��$$�oi�vWD)��6/�j�
�Ҹ'�R��!g�"�A	uk;�i[�#*א<�9q�)�L�>��DCx�֨��b�{/��e��dN��s0�UB��6�>���Z���OQ�m���>3%'��u��H�%
p���r�m�oi5�˾�A�0���;M��)�����sh��mN�2��?��ćиó6��נ���<��-� \���[����|P�@�޸w�?e�7d�(pղ������p+��;a\�P����y�����㲻�� ��0�� �m?��+�g�)�V���a����V�f8tr�s�����:�Wt��gՁ�}A���2#��+?��{��ni��cQk"݂�(Tv @���16`����`�.���y�qvl|,�ߤ�rŌ9�U��:��|��/����`|4��a�I{��V0=�x.�J_�c��.�Y�+��A��i ��1���v@�xTbG�m��Q�7�v��z��8���F�Yl�b1`��t�}�AX�Wb%Լ�C0���[ڥXjb"_�{3���R�����ZX"=X��K�s5��PP@�0ҋ���
_�s��W(��f�ὴ�X�q>O�~�!g�0m�swSn�}vAf�l��} ��z����%���Q��;i&Qv�߿�H���A�G}|�Z����_���<��\�>��:
�Z:�)̲�0B�t�N�V���.ˎ��z�ͯc5���l%m�,�&��3E`��,7���Cx:��Iǘp /_π���F�/G�]��WRv]�k�[Zvd���d���g�,G\�`�c+��P���m�5&Q&穳ީ<}�]xX�>�tW�,��j]�!D��_}L�R`��殂��%��f�����kï��$�ēL4�y{�-�.�'���?�+}�;6-hU���q��ب'��Xl%��D\8L����vj�9�+�*R�X�w@ t������ؤ��չ��JeZ��
�\rf/Zx0�:�{�w�<c��PREǉ�{4ܷ��N��g����|�j l)���Pc��L��f����\2��q�L�WK�����Pg�9
x�����BJ�n�6簗 ��xU%([G�`�Ţz���6�&�g"�nv��I��<]��_O�J�-S�QfY�l�/�
K\;�%H:��U+�QD�͈n�>��t�ll��f\U�};P�Z�W+�,��8�4�nT��As/�ݾ�O�g{ǁgv,n�g�u�����	Tp��������R:*�<.]�,Wy��b�f�o7�?����9��iu�b��W�otQ�.���e�>�(���4������k��F�m�-��Kx��Y��9���vBUrOiN��VZ��x��������S!c���8�_�M��#�}Dx̯t[V.H�����Y�n�]q�����M�k��H���Z��������d;%9P-�((�ܾ;|����\q�>���,�ȫ���>-}4 �,r~:�
K���$�f����80mѶXv_nH�nv6$���x����.�+q�j��j�J��A;���Y�	
����`�`Sf>��ǆb�Kۤ�6o39�kɦ	X��)*ui.�/�o5���b�b��C�jь�<����/�K�?�+�ރ%���=�B5�9�T��4㐴7[hK���8k6Po׊�� wٱ��1ut�.�S0���Rz�3^Ld��1�q���#v�-�7/�����g��e.v�U3�R�;`��"�-��cu�ͮ��WT�$����Lw�6������]�YZI�����i�z�݊)v���Y-W	�o�����$:Ty�b�;4Y�~}� Ň� ���9��~�ߡ��Jͱq*6�h�̞���>���1�����$ԓ+4�|��h��\����2���C�è�>�MП5�ּ�D�QÂȔ��2gA��Ǡ�^���g��"�q�]_��j�%@��3�����O%@��J��Z�W�t���@���F�~{�U��'،컡@u���UY���0����"}�z���v�-v��&�x-z>��(?�����ˊid7����c�e�,��)�L�,�������Lj��U��#l)�UIX�n�H��	p���#���p]��*RP�u-���'���(����QCE������	>����!�w�.=��im�����Uq���ń_�v��2��w�7�#[%��G�5�P'n9� z��F0�=-�p�����a�f4z���\��\�q>Z�d��sJ���D�2�,���+��)�F��{VBGM�,'P�� F�8K!�ޡ���3i����d�+hA5�U��F�s'�,�l�����y����\?h�IB@-x���8�[��\�?;D��HnH�ҜoܧZ�N���B�R��:�E����4`P�����{�Ê.ptdp��v��o����'43��a�*9;t�r$-���ޥ{����y}��=Q�V�D��{]�u�w���3�T�r��@���ipX�}�����
[�6�.��YQ�S�S��H��f=��kϽC3;:-�t����]��:CI�55�N��pw�A����o��'a�;u�����ǝ!��w8�#1��#W�&-���0�B��܃�:C_U�r�~p�~Y�Ǌ�6TU q��+u���\�/�$�j�sBW���Q�Tj�}#�b>����\@�T�X}g��on�"-�&t���~����� �
@[;w�ӷ�'{�"%-a��������*p�u��I`�|�P��ޞ�U�l>HT
��F���������ˎ�͇&z��V0;�G���19~o��jB�;�a3F�!@��h�p�TTû��|�6����	���W�O�J,;p �Ȥ�������iP?���.�y`'G���:���m��_���wf�-\��t�Dd������Jߒ>�(7���`m�d;x�Ր\��ww�kQs��9�B<*�oڧ�/ -�Ai��N����z�s�m>��$k���?��=��N�� u׶�<���s���g��ڟ*Jӎ"��@s�`���6�YU��2B>9�W��������eg�A�h�d��v����l���>`�ׯ[��+	T�z^��~���d�5.��^�3^��V`{0Y�x3�jXw�I:(�^B̥q uo��4l�E�����$f_!$��?(z�t��|���A~���C az�^[#NʳMz>�v�<�܃���\����o�&/��{�Δ�q� 
]{B���#a"�|7���\W�Z���E��	A �<b������P��M��
|ba�P����ǖ�60��w���̤�ױ��F} ����f<b��
&����#S&@*�h:�	����6ý�6�1�*#���v�$���\��Rҏ�<T͊�MQN4�e:�e�A�B� �����FA���!:�3��CCcAOq8��4�geDu��\��E;e��c��	p�����Vo;�T�KDЇ�n�]y�Q��|��j4����#̭�tª"�SQ�a���w��zq0^ǘD)va�`���P�k���9�^ܘ�Fa�N�/��N���p�:S�q�
�1�pvw��e
��0N\��J�7l��v�\k�MfƲn7�4 Ǯ�͈�b�n��6�g�uX�7��鯒'��o>>�n� R[���
C��ם��y]����x��Y����u����E��g�f��+�c� ��_���/d�T�Z�J֜�6���;�;�;ave��7�+�@��Y�~��� �m�)2qUK ���=��:�+�İ-�8p�uLH7/��y�Шo�H��$N��dK'*'���#��y��{hWPw!~�
�c�`��#S\��+j�QN;-���H���1Em�
��3Ǟ�r[�V~u�̽_�vxG�\�3P������⍝TT���V*lʦ�G�a�o�9(��:�*:��
B�;��Gq��<�Sț]~���i��*���s�*q�j�[u��D�8�v������$�n�S�*�Ӻ=٣��ȧ��^}��
�q¸/��H����p�_KkO�*)Q@��1�&�L�W{����x1�J���\���	8T���~���L�0�N+ḇ��z勴G�mXPj�Z�<�(v���*GB�p��ud�����H������������x�A���0�iO{
ļ,.�D��|���@�J��R�/���N�i�Nf�Ò��hgnk���a�*�-�!�.�wd9i/T�e�@oA\8d�ċ�������H��.�]�UI�Σj��8�6E�1ĕ�ۊF�#K���U��a[͝���"oow��5.�Dg���4�>�W�t��sƖnD�\^.YD�[�F�!���^	Q���n�cs���$�GÄ�9=�+��|��$���7�gȴ�l�m]ֻ($�T×�w:�����}D�2�_���`�V:NN�/��F�2{ˌ�e��5���4�15��o�)}1��qtI!K�ݐ�;9�F:\c�@����|�1b܍����Q{��:y�}0B��X\Q�!�s��By8�,J�����%i��g�aR=Uj PrKQ��srt�e�r��H���p62�'^�,�q��N�Ve�EStz}�ACZ�k=g������K�����u�]��w7~V�;��و�o�N�"�k�ŭ�����ŜR��/h�ן�t{i�5������<a���ow�W�j\��{�����{�ޏ�g���"���".�.��A_�b�x��'"c�����G�lQT_i�u[�k:�Ql.�i���־}�JL�������FA�d��Gt�B�y95��l�p�ڪc��l�?��;�ޕ"��_]L�6��V-qw��%4������>�79Zo�����o�T��	u9��FQ���>�yi=$�ӠT�ɻ�q'����ҍ�T��!{'6E��U�ዾ�_���M��Җ9��U-�~���ǳ��j�(�1���������j�\�9�[�D�vh�)�o�G�bg�E:�I���uF�h3��j�	�o��%���@�:6ZĔD�f�궡�S�_Õ�ܦ�8�۞���z����"43��e�^@\'�b#������o0З[/t`�8�U ����z��ߴ��A��l~M]�1�>*RaK������ƇG�rw��A~=�8wa�+J�S�2%a+�*̓�'�L:P���n�A�2�(����G5Eik�� ҭ�&�Y������yl�b�U*]HlYJgqX��XW�<�%�)��Os�*)��z�Y�V�|���z�K�F��LB�r0b]�%��/�~`��+�NƇ��+���U%9>�ư�4�Ң�8�Y�=��]"@�X�Y����N�_�/��ԝ����~F*��6;�qpАȰ�D��z}�������������P�E�n^��
~�ӏ$�A���$�?{��֌xL����cל���جSRq9\���8�Jd֐�H
u5�q���N��G��Լ�8'D<�fA�=�b<ͱ��a�^�}��jb������Z��.M9B�c>��_�F2_�uM��'fQy+���.,m��6�ġ���Y��<����rTm���XU\6ΰ�*���1�g��<%%�kv�4���������~���k}���e��%�����/�t�5���O��π�|�_�>W�VEpq��9���F\��UO�&<`��B�Ȅ�Ԙb���_�tt?���O�!�Ƙ�9�N���a[&7�_�Wj;�9���k�h�0U�̾�j��f��&޿��8�Oc2���*���1p������O�{�b��w23��R�������U��K��l��G��Γ���Ջ�(<}2G��pj/^��SAh��U+������d+0���!z�u�o,T�z��r�;����L��᜖c�o ֔.�^��]|�>s��̬��⭝l�;Nւ���^�o��e+�!l(�x��11��L�'$�nj�׸2zV�F�����ꮝ׀��A�b�fo6_F�d#��U��wie5Ե)=�7��AW�.7譔��D!�`��CcW���B�&����|}0���X��Eɐ�H5��Z�48���W�H@D��[s�;{K�T�k&:HX%�
^����=c���N#,� `, �}�gb�tԔ�O�m�z ,8<����Cf6�)A~;l��F����6�2�͏��q/�x`���^e�j��a�%o�~h�TyVJj?��6zN�2��S5�!ș��m�w����=��	T�q>oUo�����W�OG�8�����xi�d��gIgR�S������ٿ��ԊZ���ls���x?d��Js��v��j��z�Q���ո��>���n��@I!䃹��/-h�|s��BB�U�;��~��9h^�b�w5�p�w���NG�RX��1`��EeǇ��DD���kP	��}K��Ց8N���ͥ�+�a�����kp�4�0u�[�=o�'�����98�a����\��C�}���4 �z$J Z;j�������������Yo��H8}����5��c�k��������9QI������K�"�s�<sA�E�x�X�>��"[�v4��t+My=�����\/&�GL'�f�����{�`����N6Tg�|A��B#���:c�)@Y`��� xYŬ��D$��(���jk�j���¤�l#}�ʠ���D�|O��^�c�( �����a�d��KR�Q&H��9�������{���u�E��Ѿ�V��.B[���f&���5���_�U��S}�4�D�T�ߋ�_;Z�W'�s���C�rz�?����
= ��J@�e�w2Q]=���'Rs�u+8I�Ѩk��*	�D
�T5qfT1�(���|��Ϸr�ěO V�S�$����ːf&xr��;h|�i��q����I�utt�iF���Z�5O�XQ����� �	#� �I<5(r���@��'��h](�}yV��֜v��[�������^m#�1�b�x�?}a�E'�5�q�-@�Dob>��
̷�7e�F�F����ݜ!Ȧ	��O��p�DP�1���:��~�:�]Za�ʹ��J�v�KF+��d:��D�����eiK�E?��?T3�`$H��՝���"�P�jY��h����8�����)kk�g�V�u�e�_*��3����޼���=i)m���a�-442�Lb=��Hŝ�}��+ (����H��H�������sz��S�p�C9��DDXg5��m���n�Y��QK��%�����jͿAj��B�{_>fo�N�T��ֆ����գ��8�S۟���5���&�^���d �V
=J��n�/qUg#���uk����Y�夐O���ȥzN�\]��(����_c�@+xP�V��ޫv8w�7���?�땇�d䯙�h���%���uiQ}�
5�?�7u(e����;ź]��L����1�w�B�;y'�~p����8�'��l �j�)������4vl?�	X((,m�Z����^�_~��*e��a0��+ P�������H����̚}G|�`@���GN�t-�/T�N4�g"
;�L��z�����	� P�-�H���}B��-�\�_Sc`>����h饹*�A3����9&��i������A�y[&0��a�
(�'S;��ّ�g �f �8���p0���	 5�T5D%��c�� �.A�J��e'�Sl��*��P��D��R��wʅ�`��Å5��� �"䌾}�����#<��G�� Cuʳ	)�$ul="%��c-�>,��q�۫~����!�I�2��O�!��Z'�*������%�66�H1!�$����Nx�u��}���k�'䋎���e/ �x�k�}� �@=����Ϛ��m���ƣ�k�����w>x��L��|��!�VD�V�#."�OcŖ	t��	�j�(m�|l��������$t��Ӝ9�'
�k��]bOt�>F/,��ҁf����'��2�zB����!0]��;��:{����y��ȌXq��ola�������9χ�4��x/�}!�����K��)����l��0�r�]|��P�*�]���+6�G���)(���a�2��	}��<�3��j�ל���|$E?̻���R����N��f-�{Vᷖ⸛��ɞ�:5Edx�E� !��D�%�lo/c��*}���Ed�S-�j�#
���UB�j\O~>��h���#�ʤ]U��[��@)�[`u��&Ӏ��������%��2�ŗ"R��נK����Τ�G�;ckr��⇎G�Gn �<��R���P�������ݠ�B�f�7C�����cƑh�(🜐���0�x�,ܰJ(�Dj�����5{�.�
@�(�Jl�0hHlX�,G4��蕵�����2��>��|4���)_�-.��+v:Z��-ǲ����(�/�
�d*�Eǎ������Is�^����ʬ�h�k�G���!�R���i�V"������Zdf�:�j)���:��y�q-Lw�DR�]�щk�?s3Wʁ���lMN�\����%�Ʈ>+&7���g.87k�-֖Xn���B���|m�/>��ӻ��� \�J���������ŕUuX�=��-�����)o�47���-o�1.g9P�x��3�9�b�}��V<;S�i~�.�LH���~%�շO��K�a뮯�L���̅���A�G��"�+1�+����KQ����V��nv>�^^@����n2M]��6�@���he����d�"�G�_�T�]9J�߆7�����ʺ�om���|j��F;�=Ԍ�JR��|���g���
5hk�+h�$g�IOI��z�\m��BF���t�|��P��]�K`�4D@�i
h����ŷ��$���G 2��J����TC �Π�ů�6t�>�^3���*K�#������_�্/�_�l���r�K����@Y�,��3��#D�l�L��g�Ǧ!�.�r�a��Ϡh���J�����8���L��k�T��3P��sZ�I�%D�BTJ����.�_������5c)�8{�{��a[��9���Aƅ�^h��XGd�܏B��o�J���xg@	ՠ7wEl8}+!<����s�oױ�'�}0l�N�ޔv���s�}'������ׯ�G�ry
 ��@���c���x˱�;��_US��LhE�f{u����;�q��w��}�7��������<�d�ڏ��7�Y
�)�N+��7�B)i�6��-�J^�7c�?���Y��Ƣq��
tK
��[� )Ն�)(S�8Oq��?kkB�9��2dh� ��*d1�Gԕn�^��g�)d�	hL@�5y��%�J��}���l&ps�� {��D=�IGN91y�T_�s�n-�q��R��SNF���(�](+�:PB���n��[J'a3�|1y)ׁ]U�M���,���fN���a##�<����7�ȕ���\?I9�|_U�/�9io �9������]ƥ���q�� Z���ӭa>%]���'���W��DGw
�� 2�����;���ʛ8w�ٿeJN-&��9C��-$t�,G\�sy�¯\K�^��F���<+3�t_��҅Z�_紈%�7	n怖GHg6���|��}����T����7Փ�r,��� mx����m�D	Rk�i���w>��2 �����t�sv����_��@���J]��
r����.�}]������~�[��I�<_8�H����'�M����~'��a���c�L�����=�"H=^��������f��Ùr���p4�(ed:t��d�u�Zߪ���]8�Ԯ�G7��1������;���@�/0 ������XQE�fm+ÅZ�E�#?�\��k�������&��̔��9O}�Qt���%,�+��2'6�ش��ާ��Z�_�����K����?>AK�)�qL��vQ
��</Z"��G:�j"q�UhBB�C%వgmc� :����L�1./jh0�p�o����R/i��!C&�(���*�]Qk�~��9A���九,e=�z	�����c�oP���`g_*��j����. (*d��3�V�I���SE?%����!��9�\��x�p1_-�3����Ocf�}��J���@��>��
���zg J����� ��C`4��t#�gг�e@����l9 F% ]' ��!1�+ݑn�3�e�^�����x?�a��9E~�(d˩�RH�G3>hb��?�]Z��m1��3��薻�f$�A�dW�2�0	-�]�ۉ���rA���"��5��P�t�������Xd�F5 �b;*�(6�@��{l�����	E� >4�˰5���n����V�f���"Nd�����1�[J��E����z�R�X���ۏ�p�/�,�Y�K�Q��3�z@�z�)zL��?�U��}a������2}��u5���˚�#���[n9N���7,r�y��� G�?���U��CS�߷ �M��.��&Z�D��[k<o��п1	�.�W�~m\^~�r��܎9ԧ�T?�x@B�HB����\��@#A��Yz<A����?���s���ޤ�ѵ��{�a�)�띒��=��y�OfKo=����[�S��A�*�6��;x���j@�.cc���rd�1�s��'���ݬLFF��8�vn;�A�������	�x'������.x�w����|�%�K]a��4�D��.�oJ�)��K���ne��������չp�\�R�Y�/
��^ ���|�?��,�l���1T�VP��,�	,�q��M)�d3Ǫ'���S�P��;���V
{@#���wCV-�_����kOC[[��B�p�PՓg���w�Ԏ��X2��r<�������t�����,6Y��oCm���I����f�^E���o�=�
�UxW����A���eOKr���$Ȝ�ﳴp��S�T�?V���9ZC\���;α渐m?SP�"{��?f�]�;�.%�9��Od`q�zH@���Z�2���H�hk�����5� S�"^K���hiG��C�6�
+��I�Ѵ�_��1�(�yCY'���3�a,��(G�ɘR����+(�?����DI��}�jcO���U͖yF��-��������ݥ�����)��̗��և���Wg�r�JHL��󵘹�g��J����Wu�I���?�������qt���T+���\������zr��%�y~���z�]v��x��煋�!CbL���r�;B�����x��<-��`Д���L5��s�������4��w�6O6rRvR�(�\�M��[K\񺤦�Y�Jq��s�Vz S#�r����I�*JIu�`��E�6s�X�"Q�f��֯]t�����o8ui�r�:��oI}%��%�������Ck����o~�OW��7���21��5�0��<<ĭ���ґF����x�w���7��V��9�|w�~z!�������u� }a��h�A_��vG]��+�B�/j�Wc����7M�&#%Q�w���f�m����1'W�s׾�jz%E5M��Mq�/]J�>/ȵ��@=O��0�UU�ڥ;܉�oI���M���t��V��gYOTy�w����nńgؿ���U���=dh���_HjU�C\^��z�P����'����lĪKr�!���CCk����k���@)�PD�\t#���݈tI#���f�����A��\�{?~���w�������<���,Ŭ�� ��E6j#��%E���m7�8"O��;گ+�Q:��Ȫ2�6Df�R�����^gS�O�U6�����f3�m)zfr)�=�;JT�sƉ�>���N�F��h�o�t�B���	���1�s���Q����|T�(A:�K��Y�F�r���1�8���Q��`���[���<�#�҄��G*/C}���qS6*h���`���2nP�Z��O�V�c"��NOSF��
H�?�:[�Npt����4M�5�+Xu
(H.�Qr|�Y��ĉ��V�`���bPg�������?�y��ؤ�Vs��B\���%nw��6�(x�[���B�TF��`�?g�
^Έ�,���3%3("���J���Kuf���,o�#���Ģ��r4��oq�%}[�#�+�����|�M�F�4�Թ|T�a����/8�&��7`-���x}J.�}�h�����؃���f��)q�{�}���*ܐzPǜ��3�R�p�C�)��-Ng�?��~Mu69�4�oFfP������[�A�}�&�?�6$����s��|�n���\�W��������sx���A9FI���6(���R�?{_��/��\�ӂD�nA?_ؤ��/�����fGZ|ޔ�uf��ݏ�f����"�El�۳�t�k���@q��'e��E�s�B����$&,���g}�xٌlI{�����JM����C���u�1I���|�:J5�ɧf>>���ļ�����}y��DGǳ��\Eai*"�����֕!d_�~�?k!�P�\_��?o��lz�	-w7�ٜ�-��t�;tj��� j�<���Hu��b�����jW�����@+H<މt3_�Fw��'I��?Cq�M۵A�||X6�-V���C$��2���{��VJq�N�<_6pq��
n??��Ζy���ks�>�.5�S��L<=5
|���ж�[1�bcU��"�����^��3������W�T���]�w[C7Jmo,q��	��-GQ�f�)n�]�J��OW���W�K��ҡ��Wa������U�^A�6�h�ѹ�	8������i��.Eףd9���i?���țN�i�l��'SJĝ::)���i�,�N8�TXp���,�����=��_��N�'���1�3�(�A��;�16���D�c���_O|�K��t���b��6#��\]�i�T�&���9t��Z'[���p�o�UO.����[���J})؋���3�bv�q�!~��-�x��G�	��c�h7Z��Z���`|�=c�D��F1Xeǹ�>��&�&�ưh�6�x1�\Z��gvj7�k�]�$�H'\���\:�M���������Eޤx��*гDe��f�g�����f����g��7�u�6�J����
	�Ƭ�I�R�"�d����w"��]-U��g���e�֊�C�"I�Tg��m���zn��r�H��qsfQ�au;Sh~�:�=��HF:�<�	}���E����\h�Q���%��ų[��z6x�_G�qjv/�;-�	
8O����∬�".��y~;Q�m3��t�a8u�.m��Ԯ�gD\ `��A�Vmvw�~�,�r`<�ct	L�9�8B�o6����p��}�5F?��$����㽵�6I�DF�(/�����wW����3�̈K�?���D5�G���f��2剢+&?�yu�d���փ^�ꅑ�G�E'w���/E��LB:��~k�q��(�L]�M��t]�g�j�S̈́�1�4w��[}Pl�L�T�J*��l��Rӊu�@B3ЪQ��^�t��u,��O5�M$n�2x����'��1J��R$��ur��r�U�M-SO����M��&ے�O���l��@���"2"���Np���ǐ��
޾�ǵ�0����wv�#�V%������=v�9�Y�y�j���*�p�?T΂շ��/���*	��R����"���?�C-}F��)A��Jo���L�b>{�wCd?E���j��f��K��pY�8�C�"��px�wT <)b���OuU�s��Q����e�TՔ�J�%m����)�P�h���Е$0>�?\��|m�&���s)�BE����86�Sf���j��А�1���c�$ؿ��F���e?1 >P�=Ղ�[f��>&z߷l����|��q뿐�Ro��ȷ"t����G��ݔ��ϷX����>����.����.����.����aߠ���w�?�@Ng! ������	��������ƪ����0K�Jcc�[��p�s���-�2�@ �L!�r��+11���a�/5W��,����Ё�
��ƗHV�ժ�vt��
**Lvm꒒�����6�9
��ʬ��Ȼ\ll{�M�%d�����k�Z��K���Yt�E����zVm���;?G�T5���\�Z{���h~y9�����]�lR����G��", @BK+��8��s$G(�t��Ѩ��P�DY~>d1�:AK��U�K.��U�U}$�
ӂ�g��<��<v|nn����i5���p�@�9�Z���+�-�cUFa�����h�G�͒*,���P-�ِDR�c��6׋��t}�:�P��W)��\�"m��c�u����3�e�E����^��Ơ$ats�\K���R�V[50FPz��6�����'��'�y%�$H����||d3���o����l;�#=%���G������\/�����|ae~[��f���%fl��N�qu�Z��@ꡡ>{�"��o��b�z�"t(M�m�~��e<�ネ���IK���|ڛ�s�oL����V�������tW�z�+�o�;�gԢz�Rv	W^�Au�t}CN��`��֡!N�]$��Q�R>����U-r~�`22����!&��kc~n#ô��-��C;��*�7f���ӭ(&~�o���)1��Ɠ��,�w���./�Q�7�	�����밌q�#�����Qf�a�˅�V��v�#������_L����^GD�Q���Cϖ��f{�b�+$��1<�����Ĳ5$��"�z``��(t;�>��
)���MF8�Џ�n�O�%�\Lk��	ߌ��k���TV#!�"q��Z���-�ðlE�<BX�Sc�jվZ}�M|��z��XnC�-��Y�՚�ݫ��Ý��a��PQ֙~�	�o�!͌*iN{
�!!��q��ߣ���-�u�X���%��
���'�		����Uvo����!��ټ{'Eʃ�N+۶�k�s|I�)��'��\#����k��}K���Dڼ����ڃI$,%�s>��qI�������@xnm|���\hO��1�?���,@4I�%44QT��Vq��%�Ҝ�l��q�
5�!�4�,`�IxO��y��jf�c��5&����'y���l>x����#�S�<!�3��LR�����褽x�H]�
���Nۗ�DH���G�9�
���Zh����uv�~,�A-�he�bHoc/\,õdڇɭ8��y�	M�Ί͏E+�.9 �0�$��$�c<'���-0~ga\�	���<��k$$�m�؛�8"��=]KEY�����qh����<1>N���;��Vhh(�R|�1��8��շ����7G1M�E4G1Ȧ��l���\uj��G�5��z��z�� ����%6�'M~�煼��v�����q���ut(��~,�~�&K��j}}}���� 
�t7������^hJ���F
�YWV�Z��	�������lَe��6)��0~�HcSӠ����x������?��ʃ��S�����/ۜ���?�ۿ�Z�[)�hɔ�^�?YX�ґ81�\�"������+	��=X_��lh�O��_�ǱO9�����rՏ����7/$ۊ>?:��p��i��@w?����T����N,	���'*_Y!s��������<��Y��3�?aD#+))Y4���!�h}Y��i��'V�;}�矍��!L�8/�bG��A��Ǐfg��1Ȃ***�MLccc�-,����ero<+/+�ECC�[����F��)��r2�z/�����&�Ze�6��>�(&�Sv8%x�$i�4Q�4}�N,����O[������-X���'�� �_���,�[�㑱��|%D�1
FY��p���x���U�(��񱱥e���h
a�4=l����H6ICMS�n���̹.�vHݕ"sK1d���G�S��-چ������;�q�P(�fp<���y��ő?������z�$))	}p������O�~ϲ�	`*6�;^	��V-��<��C��T���@�E��6
��c$2U���%���+{�;:O����Δ���x���=>nC	���q�����������3�����S&��^(������JE��)9��=�+:��y� gE��/�Qu��j������"G��*vyg�|���hp��:k������B���������=�LyO�1�����j���%�h@[���3b���n������$����*+E߽k�Ȯ�2Ih��`bbj��t���CĘ^қ�����RP���5r<1A&��� U��Z��������߿����Ϸ�sIn���2��Z�i��yxxL�aP���@�sc8=_�S33B�ǡ�>���)I399顷	�J�+��}�VQ/��Xd�7�@�"�#��Ǥ��5�Q ��s{���bw���i��술弹����n8�HԷoߪ<��+Pwf���WFT�+��o^ y�Y�x:�~�^�v�:>���
���������pp��LYM���-������r���g��{��E�^��JF�qWS���� Lv��ήA�������A fOK���!�kE�.��t���D��*�;.f�)����|�(��h���'�㍝��t����/�η~�^�ALBB��~�^�L0%�`}����+�8�-�����m����,)�dS�s�#���_��Z�98n�8�0�H���O�'��.kXvL����{����f����nVۚu�z9���'���;+wm��G��A�A?���H��v����n[��5bg�2�o�G�!Y}x&����r�j�����.S���8-;����+�k~&h�^XWOOO,�A�ĳ��������%���^Wf�<�Y�?9�������=o�O+-ewqqI������v`���_Td�R�����MѷQ��G~֌���8[��.:�Z��oً��3
o��#A2vWx%/8%�N|@�UY/�LWYSj��Шit5e ?��\Xr��[wF����A��c�3w{��`�X륟�2���5���|@�hz� }s����.p�����lSѿhʓ�IF�a��ؙ�L��zzz�c`����w`��,��okk�HIK�{�7��1�x��]^�<YI�����V
�H�*��{����������R���6HJG�٘��)C�NcCf��uz�l���7����8���3��M�y-���Y�Hn^#22rZc�@B��R������%)�v�f#'�L��o*:��:+U9�!Qe�쭬
P�P8=dX�܎�DAAIol�i�Y���6�����g��J��	�:#mO�?��ZR��.d�qJ�������+͍�Q__����Ӈ� =��'O4���Pvh_[��[�<i�N��Ǹ<�٬��7��RY����`�pQ��*Kǥ������Đ���\[��_����6�a#�Tu�!���OZ$paD�d�p��3���CҪG�)Y�,sin�dhd��`��5ⴟ���ψ�
�I�Yr��Z��Pv�?P?�0Ր���{j�7&+���nn����]3P���}u��t�w��zO:�n|�Λ�a+�iMNM��2�7555�l��Q��(�IK3H���&�c�_&��W�XKқ'�n��6���4����4c�X�� 8�^��J�������{z�ޒ�.��,ܮ�H�&:�Mȁ@�\s�H�0�78�B��xp?���P��/q Fd9R��[�չ�(cb��@�YE؍ɇ[�9?��h��S���W�YoCA���!���NT�{��N�S��;��,���.Z[�[��K��ᥘ��p= �ON:~��T�%�r1J���. e����2���˙��$]zH��+.���t;���c##�߿?�?~,,*�ANS�Y Bm��>i	�y��\ `'v�qi<$�/4���Ru׾)�����G���}������S���q�G���;yڻ��4ȆΥ^~Y����s:�`6�%�~Yu����B"�@�����хiG�Ң:�j�$�+C��A[���ggg_;l�کT��x�*�+j6�������x���IQO��>�k�gӌ�t�\w���8��$�5�Ud	T���<h}��Q���r92�V��>���:��ڿ#ȍ���|���F,��N���r�蘘��)�5�ܗP.��F==����_�-���og��#=�@���jrp�,w���ea�o��E6{��"�j��?��Òn�&_�r��W�l���B���@H��w���ӸQ.---τ����������̵r�����K�\I��_�l<$���z��7W|b(H�nkru{��@}���.� �H���p��n���v�N���z���KGkQ>�$��ܐ�)���%��\_53*� .� ��$}��'�� ��ϝ�ʷt�M>;�J�47����XѦ�t��c��ՃM9o��@M?����w`�f�˫B�z��ug �Aٍסk�z��H��`"m�g�2�h����~`Lv�;��u�@�4X����r I����;�'�nv穵�S��Ĵ��e�5� ����慔j3�Yt�R.����"���sZ��o��ܸE��7׀�$$&����_$ƫ�O@��4��1�`mOO�=���=�Eב�s��%���(A��;:�h�XJ%999 �b7�����s.$[ۉ2AY儎ix�����z��sr8}4�P����,�1.$�Ԥ�l�O%��"�:.�~w�H	��u>_w:��=c�����pM�Rk����E�NUi��ޚ4R���ζ<�O~`V(G������\(䗗]�H7���%Owy�9�l�9�N{�S]�F�xf���)�g���4�[%�%&ݑ�K�ŐJpV�Y
�J��ڳ�g�g�%|��m2��S��H�Y����o�5���2�\Cv���D-���؋j�2n';H�Ж�g�D�����3&�p���!G�^I�2�ׯ�|��L�IMEv�iN�yi]�o��.��HpEEŦ/ �Z6��3��� ���������>̶��A �=��C������V�40K�蘙������U��}��GGG7W[K.�	�otG��c�'�Ǝ�C��������݊�0����K���8��� q�a8��{�:!��3���9�zi�cq򣮎T$�Mb=ڱؼ������Lv���-�_k�p3� ��� Ʃb��yGY^锡�#:VVQ]]J�)���/��57~������wS�睋a��All��;IF��>a��ؓ�!�[4��Ett(���t��}��c��������'0 `�YU�ͬ�|��@/3�c%%�b��w3.��@���P?kp �mo��f��ؿ�XH3��B�p[a��H�r�Ӄ}R���H^B$e��P���8V�j��ao�+�'^y	Q��N�q� ���FH PMK�7�D�լ�u7~���?�܏�٩$���h��&C���?���W��Կ@����G&;X�:2b��y��w���S��eݼf:�ߡ���X�^Y]L��]f�P��Ibjj�56?Ӡ�({(pvV۩�bo����R��b�m�⷏(����"��EQYy���p��e ����S�'x�^{��['m����	���nV�o�p����v�P�mm����ѱ������^g�p�0�w֘�Yc�����zr����aFv�(=�'C>>>ՙ4��ǧ���:e�Vf@`�;�I��e-��rź-������P����ʆ���~�O�3lo|/����P���l,M�\%�*��\���jn^^DRܮ���I��ྏ��!�HU��Z�����,���x���z����R�f݁}rv&���Q՜�|Z�_��"������m*g!⏀�w�4��>`,���92ǘ�$�GUU���,fl\�{�ʴ��^����	866�@�3I��9w���C�TQ�_��^ZZ���}�g�&$!imjB����i�n_/�9�����UO���	Y[]e���G��}�z��
�����G�Sd{D��z�T�
]儧Ň��R+W�������b�]�!.>~ZII$J![���du������A-�V���M-���o�u'�?��������cv�668�lP򪄸X�YϠ��� �j�)�[ή.������N�DEDx��8�˓RP��||n��f4�O`��xubqQ^J�;��G��'�oٽ�Z��h=�7���&'}��W^N��Z�m�1?e���Vr���AV?..����b/�~�~ʢ�P�>2�1)���N�
66<�����륨]"t�q`?��x�F��tt䪃����/6S\=$*-�{�I~YS�Y�m5)~�c���B �ڞ�j�i����q�d�U�������C�U�*̴|�+��P:�hݎ[QI)����A�k��yyh,*K|���-d�g���@��#���]�A��R4Yjjj�+����!����v�a�n���wVx�7����M�����&�n`���ʚ��~���;�Ӫo!j�o��ިEZ��Ԭ�`y*DO#�\kk�`�B�܎��%+�j*��3��~O������I;]JD2�(R��WNɫ��GGG�=O��\��I��E��Fks�%�4X�0��L4{�ik謡adD$��\"�dj�

:yo�s�"��'�7< �N�3�;
��%�����C"*��֌���8�����$�(��?�y@�*��QQ>55�kv5 �)�؏�"���q9֏�\���'��M�]$P�,%de>�v���d"�Z�u������-�����wl����X�!Guq�i	%K�O\�4��;s[���2�r*u~�K~�1������]��'�;�%4��iƅ���OXL����.���y��Q��+̆��Q'�h7�Z������5��ԿM�&y�28�K�9 @L���q�`59��7J&��{���$��ށ�"�UW����\l�Y�����R���@�����{�N��U6�����de='mGd�Ӝ���� tMט<����\���^$�HF�W�EY~Q&,Iiix2��פ�ޅ����_�P�z�p_�p仳Ѹ�O�-0�	�� ߜ���z��LMǯ�{VWa�Sw��9������Io���[`�x���nJ���F����"e��2��ϰ <���V�X8�ÍVJK��ԃZ�=���|�p� ��ΤS�w:�v���ʛ��Y#��h��f�C��Rϗ����Q�L�+���]�O��=,�z �3,O>~t:8[����%��k�:�VU���/�*Ef��+�+�(*�[a�Is;c�E��؍�/������mN���?�҃=~ힹ�P�"����r���/GI	*�S�������(*�v
==}s_O��Fzlpڻ��!!�I1z��g�M���Q��ee�F$?y.!���)@�]�o�Ci:���&�/$���넅9�ͻ	�q[����!��j��t�����ձ������$��'�P��B����x&zkO�2T�d����Kr��0�
(��)
�Ʉ/%������iن~�w�շ㿼���3XX�F94��ڀ���� �0<�.�i��r�'?;;�u�@o����U��z����Tt\kTl��fAN��TTJLܤ��`�lB*�">��" t��"�#���ߧ���m2V«k��E��I&�Fvff�^��*>"����߭�E���w|/��t�9�?�"�"��ьATǅ|/�8L���K ��de�����?�:j0�C�o���P!:�7��Lp&?�^�7И�^���8���,�/�+���G�y��� O�:
��/�q� /^#�f332����A�����L_�����o�;�u(h|�t2�1��вa73`F�א=
�-�HK.�V�]�\�]Y�3�p����΁�^�4о ����K++z@�����F,�o���R��J��AH�hEޜ�����ݽ�\ġ�&&�3�6/���y�ƪZ3H�}!T���@�!U�c���{�D���x��ІGG�rs�Ƥ�S(��8�k������y��ꕘ��s�n/��yiq���	s�f�A��@ڋ�ⓒ�̟G\O�><J�b�H������<�%6jSIII�Q?9�h��Q~��-��Ю��OH�NO�g�gF.�g|�n��X,(�"����x�A��û�;L8�����wN�ML�͵ciBU��0:�2@�-��͠��)\�U�39�u��oԄy��w�bUmm庄A��*���E,8�}2'�I�ig��Z�B�rwD\������]]�e�[���(r<�q$S{2�DC��aVRE�x�@�w���ۀ1������%%��=o��O>fҭo�*�&(P&*�m�8!��^��&(x�����A��H���҇���ts����E�D�`�����歚�9Z�(�y��l��VSS���������(���ԝR)�8Ԓ�o������U>Y]]��R���\;"�������ǫ��u��f�4J6��(}����o�	��y#���ӺRC�b7N�]�4��@Z�02�m�K}��>�X�O��!_6J���A�t���766t��8B��gTp���~Kא7����}�,��ۀ�Zm	!n�//-}�� ��-�̅T ��6O�,�Bv�Z`;��x�V�E c�`��z�C�u��`�0�Z[2�k��B�#�7��.Z��"_���y8rX�nfn'����׷��r�|�������W�{�����<jt?VC���>Q��l��s7����������v�u�9�yed��06��8��-�99��z��Xw?~L�¢LI	@01�4�����
m�f"d 5���m�c;��W��C����o�#���)�4x�����rtt�e���$��Q�Ĉ�ls	��RL,rw��_���(b�|����7��==@�@�t?�|��=Lxw�?��M���g��Xcc�*.��6x ˜��Ѕ��� <X�FR??�R��o 4ʷ�VV d~VVƱ9SK��C��I�����dQ�oh(b}϶�����"�K^�o�m�;x
���5**]�eJ$%--
hU���f/u��H?jim�I�C�-' 	}8�R/��u���:/��J�A]�}U\n'��US�]7����@q��&y
�"53���1`QV�O����z������+w�w���%T��=��Tì��� �2=1h!��v T(�i9(�_�$G]]`��������/� x��zi�Bh����mT'�9�U>�$+S�7P
��`��o�C��9���?MT=���`��kޮ�R[�Fd=���:tKa'6ټ��d�b���T�O��up�����e����)@�Qk�ka�<@D��/M)g��P�D���s:�t����E��t�� T��
�J��pk:����ײn��E�\^Fx�G�d�y�ί��7@���J��#{�Ally�����3u��}������}�B~���@��sM�w�����z���@��xv�t ��Zd�5w��zba`h��5d!�u�-�xz㉴̏�>ߍ����g�X�����*������Q�z����T3B�z�z��(�Z3X%�BBTTA���/j4�V�D \�C ^IX��<�=���??a�|o����"�
����%�|�RymM1�p������z�s�TՈ��39��?m�4�Z{����@{�fjߥ��b�(q��d��%��"��_�8�8|�r��J)3(�����o����0:yα��s��K��D)��JWM-��OP�=3K�����=C�"..5��tɟ��J�?��W��ځ|��L������`�:/+S�������_GzLD�dk��>�9����;��������~��QC8�����H�<����f����a2b��6���(���D؈)�TY��L�D\��H�F�2��I��P�%�����!+�L��R �Q�U�z�*�E��ݺ�����|�~~�b����J :�>����"�7o$W�.�6�J���<][ۉ	/&jG;E_p�p�x����� ��z{{y��d����%*��U�-O_����`é����ٚ��@�Q�&ѹ��i�8�..� �4YTƧm,K�H��(!��Yp�b6�:��tZ���e���(�n�!ˏ��4�e��_gn� �����u��yfʭr=B�y�������y��Ey&\[|ܦ�
��Nq�H��쑠1����t&�>��ϟ?�=á�_RZ
��Cj��Y��`f�z���v�v/$ M0o�eފ�SUG$/Onr���F�Q`E��6~����V�USSCG�1��>��ty�6>�����3555�<1���)��F�Ё����-J��? [�����)uKC�����X���"M��tQ*�_W��+�Þ@������WUS����1��� ����K�[ºt�30�~�{�D5#�A�����l�X�y�o��	cc���Z�ݡV���6�b򈁛�{5؞n��/^�H	ޙu9V��˹j������T+�����	sU����#�!a��jC]��}���EC�:MA-1� �\O�}�u�G���dde�>7��C�pq�@��ֲ֝�Y��U�.��
ׇp�{xǿ�Xp���Z6e5��Ym±��D�uxu������#���hC%aGº�����8S�TB�[Wr�=:���Ti�D�����;�qT�����
���¾.�US!P�� ʋ{2���zӗ��a=!!!����m:����^���z0g�\�x��na>hN����K���/��_�
��W������W�j�@���J����Y�Tt���Y$��;�hh�JJ�BȀ���eggzs��A��TtL���3\�Jf!Ê�m����Z]���i�(���9��;����t�9��>�('��u����꼞�/ �$f���=��z��=Rb%!��`N>a�����@`^���K/Q���"�rƐ�G���sI	9�@���J%���xv�!4��b�T�2㥇@,nag2���r���6�Y�?+�����>�,�aKx��L�;���I��/ �j\w�0�f���S�/e����Ӛ��~�����5l�5Pk0�`~�g���{r����?@�SNN�_�X��@�:��7���o�UϷb��*�|��>L�lN#DM��RƂ�fd�_	9y����=�|��ja`d�WU�j"�	fI-򅶼�~ƚ�G�����̳����?B١���g�I7@�l����zq�p-�z
�����`��p�=����:��V�	q���"��#^�9��m��E�M�ň�]ja�
��>�J��<��۷��wl-n(�y�&me��0*��Ǎ �?�8�>V�v؞Ωr���@ԙ�5( `�,9�se����.�:ff%J�gy�/���um��I=���y3�!`I.�=z�������� шCE@��AA����yRؤ'��׋�@�������YY��E�c���X{����7��l�����pm�u"�o��#��RC�6:l��UѺ�Ǐ�����2��@����	Yo�����r�Dv]�{����;����x����j�A���v��@�f��{�xS��А\�� �E(1N�H���.	:C�n���Fp��y�5�}��>p+�	w���8���~Y�������'� T�@����fc,�x��}�n�s�����>��NA���^VWz��k�TXZ:55�����P��Nryp��}�j�@���Z҄�yh$sk~��%�	�� ���B�z;�bg��	����qrUS����&_qi�{F}����;j` ��<|�Y�kxun.��~����`_&�9W9$�3�?����y*=Q�@��m�3C�!{�%��I2�I<���*
Z����+�22s���� �*2O�������WtC�(N�ܬ�#UZ�}�^@�=�)\f��r��OX���wT�8������{�S[t��ti��6����5k�Q�KH�@ ��D���|&\�Pˊ��
h�(�	���7WA����u�#�>�����f�l7I	z�� T%6 ���m*���hd��r����,"2����rӄ�<%66���\_aA>:ɘi9vc7����:1�u��&Њ���G?A9��6�N^~�J�(|�=�n��˗r������w;R��z���> ��C|kC]]}�4h$�=��1o��T�Rޗ�=���J��`������:U�''�QL �=�����b�<l��|�?�<;^�ffTi_��_-.�`��� �ٖ�D���3`-�It���Rbj�犡�T.q
��r��QSzVV���$��ً��'"X��d�t�b�_@م���ql�ݷO#lFx� ��\y 
?

B=��1#�M�����p�e�1�+�Ҋ�х�����x�_o�k��Vp2���x�yi�Og�)i��@]�vR�2L{�A��+-p>�	n��;���Z
����O�=�`�L��KJJ
�N�O
����9cZ�<���s��	d�ǿg} ��)C�)JČ�+��mu�*��2MUyt���0�?g�ſ����E�	���^�<���(�{~>:�i���iM�͙<�i�j���x����ۢ�Rk$8�O�WB1��OE�ZPE�t��{�k!��ԏ�|EJ�Q��Qz��{h$�����$�>������;��耴�����iI�����"@O�Ԕ����'ȗ���f\�Kh�,)�	�!ʊ_BIBE�k��} �'�u)��	s�r [�ro���ޚ�*��	�=umm�����w��fZ[��� ����㵊�Fw�(�x�'Zv����x����$�/�GFF�N�KL�s���{ ��-�WN�t:q�p��
��ɯ��ZÍ����æ����PC�5���||dp8\w�N-E��/��.Okڑk��DwX�7o�0�Pհ���EgǻelҌ���~�X����"!1�������|��w���P��o�����$�fP遝�[/�	�~�^��a�L�h8�d���	6�<���W漴�(��[.&OGN�[ ��ME`뚲Z���x���<x���nQAAA.��c֌��_0�VI�'u8ܜ%�,ېO��H����0(�����_�^s ���sI��z��x&�f:��Ƞ� 0�𲆬���k4��S��
��NWO.���~;����>Ej�����(N$��\2{H0}��Ë��^��~c�wCU��;;;#��h4�����{����h輸4���j�AL^3�����p33�݋+�0U�^x�E���}�7"�7���+�M��\~æ)�.��s��[_�Nw��w��	�bG�Ƶ<|���/�����)��?�Ϲ�-���:mV�T���M#:%L:3:��c��E����n��A��lo���Ę��22�i+�}N���Dt��~�?�©f~a��D��������E���wO��wXӏc�y�t=�����3:&F���k,�c8}���@Z&7:�<^2����hB5ϭ$�s��u/�W�<_��ښ=b<(�����ᑑ���(][
�S$Td�>9���*H���N6^�C�ӏ��������	�//D\$�����-#�@;'4��{JNM-p}���]o�v�Y{���$���{��u�3��.��N��o��-�p[q4YbccK9���ꇈ,2��ސb� ��2�
X�;Ӂ��J�S����R�������)����c�a��^##JU3�-��dZ���QS�1�����&Ɵ\������	�^py���* ��	+�V��)��/d��A_W������K*��nZ���r�-�|��4Wۮ&aݥ���|~�4.��{/dm�gI�v���־�?*凗߾�a		AZ�Ŝs.m8�۴��������c!�S�k�&������De����Lp��p��?���~�P�ٙ33���N��N��>77*e��	�e�8�LGg��V1H���;����sk���_�^t4.�y_鮫g,zzz7����\ZLY4��� uww���#y�� �a�S猱Ќ�B�4�%W�"u�j}�#�¼k�b�.����i�����}�`Q�mt=<���<�F�$WT8	�(����HQ?{�{S��Ӱq�!H7)�"�x�����ǭ4/��-4d+�$P��4��#�j�oII�>n�ȿ���jMk���c�a)��:��ȃ_$7Onz(O�%�;5^�s;7~���l6.._��W��F?K܎��A�"y5��5���OS�����뤾�j��m��j�_����2�dM�EG0��5{9&�#7o��p'aHKK�2�`x,�]D��ɓ�?Z~����Ƿ��ZV&B����;0�Q~AA�1�͓n�lCCC�:�+���w�E��#>Isr��70������mn��KF�Ή�>	���Q��ځG{p��u�%�H��;�%��E��ԓ�`JJJ��\<F��%��Ή-?M���
dBK;ȳ��|* Ⓔ���TJ;;;�Gtu�JfdR�����%$"j��d �ch;��������y��(�v��㏀�cy�3�]�������T<P��UU��j��=��-�/""R�Pf�	�W�i�] ������+7��\d���M���0l����kb�Q4l�zB"��ji���������/^�+��)�GL)�mƻ��0�"U��#���f⫘�M_Z^E��-�0g�	�.--u���!��LF !v �B|�jz� ����gp$��֗��*s��O��4,�6< Ff��CB�)�*:�ZQI)'�����%-;%))	�����H9:��ڋ�U{0
d��uڍռqQ��CFO�����?��=6@�U��oE\p~֞?7�)IA|p/,q���_ �s����$$#���?4\PU�۾*JK7HI#�J�t#R���������K���p��n.�����ctu�=�>�{��6���(?!�Ȫ�X�Z�v�T?�v׵}����Ā|�D�\h�ˠй?�<e����@*��h���"G�����5��g�^e��1�h\Jj*��D 3a���
�	/ٟb �=���l��F����CY�=��
1d�@�Q�I�*=.nn��4>�aI�T�Oe���d��ie7[���{��1��j6++Tx����~?�F����kKy�o�'���<�dڃ�o�D�/����-1�.e�?��ȀI075��V����ݵ�^T�`u�[l�G�5՛�=�j����!5x;�=��u �K2�V?e���v����5P��*�LrRܸO��ǥyns�wq�FQQQMO/� b�?H*$$$V�IQ�b����+�#_�Ȳ�pe��g��0��ŏ����i;Wd��^���5�����p�kVo�"d��-I���������FG5��Z?���0����f�4ZorXwx$�a��C���4b�E�n��
�H4O�TQf��ly[�����
����8V�ԇ��Gȗ%`:���E�7e[PZo�26����Le�w����rk0��9�G��75E--�))+�x�↬4T�W�,�X��'~�:�a�J����#x�'���RWW��7o�n�Gl�tt�����z�Q	�7=���j����V
P�����п=� P[��gdt���:^��m�տ�gP�P������$�9���K�Y�x��]ͦ�A��`���3�G�������Ԑ��Mi[�"*�I���y�~���}���XN��꺒3�G~��<R5�[�Q3�}z6\�g�`��f����K6�w�+����n��IY}�b��W����6��ũ����DEc���|�B�������3�cޟ��p�Y6]�������$:�O�>@�66�+++賓����GU�����_N�ۥP2z�\I���%���h�X��[n�[nt<<π�W�ބI�/..�쟺������gAc06��p�+��}["�7�vr�%(yttD�j��<p,D�-\%�1���E�Y�Ik�r�A�Esomm-�~J)V�$Z(�5$��J_?�[L,ȩ ����^�L8���3��Ȉ]/���D^K�&r;�[��,A�̞��69��A!�R�<���I��-�;8\��&�T6�?w���dW��f&(AsVC����j�똸8s{{LoooR��3O�X93�qp"�`�#�1W8⡴�����L~ޗU.r�xxx��� �cB/�s������p�<�G��ݟU�`,�&ҷ���J��I�;��pv%K^�=��`��᫷oɶ����|�T�1Y��$i��v�~�s��"7�}�Ӈ͝��*�DZ�E˄IW9 �mmmM�Ξߏu.�v�+{�2d%��7wf��	�B;�:��^瑃ܮ��RVV6��j� 
����Ps����,��F�y����xVu(�G^�:��~���_�A�ɖ���:� N���G��j�#,8��!��v"L��^�~��ʚ;��(�3m����qT��l����ކq��܍��N`TQ����a���;
�U��b���������dѹ���ݥ�8]��y:�L�o@tQoU�@v���F����`h---z�g�X;;;^���*���+5�ה�H�.��7�r!�x�y3��e��C��a�����a��\݁߆��1�J?�����o�"E ���������5ɨ��:�x9��^��������.t��"�?U����;>9і�^�&�\`~��&(*�W�Ẍ́����ˡPP-�ˠ�����D�n�S�x�P��I  ���)�<l����~v>��{���=�ݩ��*�K$\MMM�)�}-��`:��w`V��n&��p�df���q>��|�H���R�������zY���J_ד{6WW�l=l(���� g���{bI$���_h�6t0>���)�^��n��01;.w�/�F�מ�`�.LYRZ�dE� x��
���ykK��8�#�v�ڴ��bw�N�#4�WP��j}ccY]]d��;A��>	�m|h����9���}"�81h�?[6��n��>Gn�OJz�U�������$������O�*82r3�0�9klK8����
�TKoY�#�0�;1�0/���2��&��TP:� �fnF�Y����[l����S��RD'�$����G��k<����u��gMa���!hI��

��DLP� 0���0�y���='���uCq#�zƧ��>;;s�PW$Q�N�i��i5�;�J��'tB�C��(�V|/�edeß|2��&����k�T�.6�m�/hC��gR@��5�Gn>��<���DnY��~O@D$���M���w3BB�J��Xx^W0��A�C��������^�d�T@�@T����3��f�N���N�I�!�J���q�%o|!��g~���d��f�d��U�����W������3��O�$nB*�@S��J��DYp�=IJ|ɛT��7�p�z�,��B�G����>(�m}���)lll�V�n�&��:���� |�@<������Ƶ��"\pxE	�|�D������ʣQC��XX$����mǨ�1���@�1[��������:L�����-~T`;�]+Mzik*���WKV�0���`�r~v1�ȶ�����d]c�x�:�i;���;-�#B�#T{�����m�����-^��7q&��XL�%�u_�#RLD�I�i������{�b����)���H��4�g�����T� ���.��=���}_���=9�ʢ؝�z�T1~~��"���������5L���xAH�ڜ��{д�<���?qdp�H�+�C��Hx4��F`S;�U����;�t�H��*;�휁��9ƛ7m� W�i�x�J��V��WԪ~02��5v��]�3I���[_�i�2(��������$p�M8���\v�K,y�$'��ǆ7���{�)
�qKdqq��%����}\�;�TZ�;~6��<Ƞ �m_�b�O)��#��l��ɟ?��&��[|k�A�� =��m�G�l�יm��8��{��vt"�xY�����p�#�`�����]Ҿ~���&m_������'-���5Q�����k�y��D�Ӻ$��ْ�/��+���h��X8-",(��ʭ�w%D�3Ӓ����ş*�'� �YXXd�3su����؊���y�E}�&!"2����҉Y�L�t���J����qsq5�p����J�ʬ�"��n#���Cx��e�����<����a�3�-4Cy�%&����ݘ�un���a�&���������E��P�ʺ���y_�2uiok��kx��M��5;��e���#�d��O�8�9�h.��ք�-�t��}ɛ��p�	' �UwO1�C����ʓ�`��47t]�<֕�����t����ɍ��D�1�K��(��A�ֶ���r���S�v��,?lS���έ�TXqw���+q�2��O���a.�hY�GVG���?~�hbd���S�c��(���.�X�gr���V_[{���f�����}Ȍ�r7�w�<��Cq�9��~�ךW�G�s���R,y��������ɥ����򨙾P���z	*�u�7�Қ��^���!��D�{�
z�z@Wc�Ax����H��S��أX,������8�R �,q��e�vO�\5w���^M�����_�� =�t��yyCy��ػw��**(�F�E�m�/cR������G�3�M1m��Eb�'k��A��R��º�����.\W��A����is]Q�%���`��ߤÇOt������VB�����ә��E�y��]�F�<=�tfa,���
������]�l~�C]���S���KA?䑫Ȁ��{�
7,2��$�x�?_ X��Ȍ$"&v��6��s-��~���eu-�d��{i'q�'���H5g�dR���U�Hhl�ML$����	��sh,1!!��@��[��b͢ʟ�U؆/(��=��v�d���/��~�ՠщ�b���[�j̡�o`��xo9R'�\.j�"?�72F �7�����E����=��l�f�ð�`�����IiCg���� |�;�QW���̏_<y�=�ۚ��WY�M':8܇poD睂����ʣ�S7�rB�bhQ�u�d��dd������¹[9M�)50j�0\>H �P�X�vU����f&*&�g8ȏ������ ���=���V񷢸�� ���G��!��spp��Po�Di�7E���� �����VWA�G�t�a�d��"��-���0�����_�Ze��W�-��'���S)G��G@���#�QB^g�xb���B"�
����ڻ����}�{�I�pr���Vu�y��+�tn�K�rQH<�X�?����/K��Jx�6a�+�+��@	tc�#_m��:9P���.ox��τߪ�}�$;;;?�۹F��a�pQI�;�6��7/v�z�d�b��=[s����z�����0�Z!�����)�G���%��Î�a�ɵ-]��Z�ih�Yk���
j98���2lcf� ���2!�Y�M�H0�VZ�E�奤��y���A���}��8����v��Cs�q�DU4�r�=�*���n�?_ER+���iL��?U��oۘ���f_�{QR���b�����w�r������[U�7�c�Q���sgd�l����΅~��%��~d�/(�}NG�RSS�QY[OȏwU[�����y[��}y�,���-n�� ��j�WQQ���,FGղ��-%922*���E���I�dIJ�aؾ6��\l��aH������|>�yE��g&�����A6�� g�(�`���i�u�u=�������!/����W���R�\����՟X5ʢ��Tj�,/�l���q�U s�'�C�yY������!*�D�#���mHH��6����^�[�=�p��N���@S�G�,�?�A��C�!�����6k�JVN�se��(
(��)��^���wE�2��B����>1�����0=���7W
��_��!��>>>�3���:��GO_�u򕃌`�||�p��l���1�c=9�۹]�������錿ԋ��'p�ih�*[�UUU���T��J*!�
>��x�e��kI*0�ԟ������Ioo��v���\��5%�����8�c�j
���K3�U�o(<z�H��0W/  �<~xkO�J��0�,,�����h��4��3Ԕ���zv\-�f]C���.bf����f�em-�����%����򖖖��h\{?���g1̸苃�<�s��u𝹹�i�����dip'B��UVc#Sr�@�h-�T��+h��� N�0~�L]t�h|8*�n������E�)h�rg���q�����W��������?���8 ��ݵ��)�:��x�k�Ve��C
`�M��3���G�=�c�o,�����Ur�)��@/N��ɗ{�W�������U�+!*ڢ�4Ր�`��|/��	n����[��/]�J�4����+:���xz�k�q2��J�1O�*_⭓��/F�}����-l�#�@feXQ�Z~م��r�������;�S��wO���CPAw�)�srr����6�gg�*����;�;��&���W���J���u�G�M�4���/���1���_�ѯ��3t6�nTV�W���<�k�����e�{�%��i)����-�j����_vDW�<�^h�����������K�'�7�7Q��>ZU�S�l5�� ��RuM�3Cz�>�`O4
}��xM���>0>E�����o���Ρ���X�̑?�Oǂ)���L�GZ03�P��1S5h���,-�\]G�p����:��͛li�jz�~��D�g��3��_�1T߳|����#�8��g'lbC�j�����յ�i���@���|��n;^XLjff�_���k0C����Fq��tu -)%o�����$6�E�(8/��g}��v�#�;
G�Uo����̋4�u����O���ݤ��)����*��	쟪��5�d�)�_�^Oo�S�	��كhȵ�ښr\����I�����s��**�La�_)))���X��<<�@���wl		gՋ�z�<F1g�yq���Oȶ���w�! �X׈���ǹ��z��+��?J|d;V���d���~�#�c�+�����m�K�C����%��{(��L֮	���j�g[���/��D_��>B����*�A*L�z{;ШM�K�G��YYy��r�Q��:je	�ijŌ��r����q����a�regF�����1E��z`jl��Tr�������p�7����Q�0V�����U�UY�9���פ^�Dz�N�ҲZ�F��W�l�i��fEH��P��v��^W}XSdN�0fE��^�M}G:b��y��_�'�1m8"����Ā)�ǄN�e*,�;�n����@UQlv�&���݂�W�P�n��0�o�%)��G�d��_DV̾[XP���v &&��2�9�v�z�u�)'�d0��m��v`���)5���V�԰X�p�[K��Rc_�E*~������ʡ��%���M�,�$��T�}Ђ�>>4�Q[?�:r!�t�]������w��6��xWS���sf���	'U���ł@��A��ׯ_�(tt.�=�|77��Œo�_m����)�j��t��K7G�~���\�l���K��V�	���ۍhD��֚(�5�\���Խ�c��c�����[^��<N�,���AiOc,�JNI�|��TaqwKR@Ψ!�� �=(�cʹ����T8N),,4FY@�!n>�j�"!��V|�M�f���P�6���Vd�@mʉ�{��Q�������[?%\<���׊T\�Dj�$ǜ���PaX�{>�\O4��VQNF����䤿�G�`�#�ϟ?����˒�֣&�dd�!h#��r6��ZZ(�}$l.y���:i�֍��o�vp��QQ�u�wI"\��5��>�l%q�r�w����n�L��Z���L�G��Þ��)p2��6�����A�w��^A$��oj
����50�<�
Y^6G���W���9Dd���rW�o�,h�������c�/.���{����I���g��1��Fk6�����
��:`�np�߬�i�DmǩwZ�s*�a�A.��틎�N��2j���Q*�~y[���X�8S��T�$ȑp��R�2/i��lDZ�W�&�Y��s�G��A6N�ҡ/�h���75��{ק����
��5�5TT`?%������}���a�W���"�MXDĤJ���l�f�n�	F������j�U��3Yi֩gZ3ۚ�-��[�	����_������Dɰ�c��"��,؞�� VuM<���ඳ�ϚkJ�}XEW�*,+�񱶶��{�۸���c��������&��ů�|�
�LLG&w��GM�g�6�;�y�p�D��QVF�c�|�ڇ}
"*��iU�0��i*��$ee���x�	]�1�ޞ������^���(U��I{9 �GDɵ{�g���vmo��?|ͭ�M�sꊷ3���N�^)�GE5N����S_����c 4)�k�������M5�$���+�b�IϤ-��gH|!9%e��AK�\���r#G�4�90��RF�6��:�#s-����-�m�>��V{fA�о���8��(U��}w��fI)���0�[x�s���E�/_ű:rX���᝝�.v�H��^r"��y~��ɰ���������[>Z�q������	U���|�|�����?�]��SP֗�����*�!�J/d:�׭Z<7R+�����Nӭ[����ik#�����;W^��{!P�j�����߿,��x���D��k����������ꩧ�-[-R<!~X���͹�A�N=�=����W��%#}]|�\3��zN��O����N����a-��g���/�ߠxxYoA��>��Ņl�mc٘��aE�<�D[;��S23����M�S�Z7��h���}�wI��@^|�(�>��z�E��KXx{�UI�
�è)��n"I�����ݏ'�Ţ��5D�Ҹ��3@̇�w[�-WFN<Ol,�����]<|a7?�I2U�&����&�ĩ322(.Ex��*VBp���*�u�g"�GY.�q��7���	�L9����:,,�WzW�є"z0�]�DbF��f�g�w�Z���~M���p�gD�JKq���Q@pp��QE��^;y��:�~*͝��vˏY0����҇��ez7Pb��T�g��'�m��7\�C�b�Ɨ�!8�!lo���u+m��Z�s^E����ߐT�Þ�`��|W_k.��>��\I�Gt��EG�g�)%ԏ���>���7��o�����'eT(�wm�����ZY�����A���_	0)��%�&;;R22���Q!L�ڄ��o�̓!Dm0eu�t������(8�D�`>���
2!	h(^U��[�+�3��FS�#��p=�}�[�o�ў�s�g!A��4�H� �s:�+`*:��2��$�7Ե��� ��@G���Җ11���U��B6t�����{|r��P��F��x�d�o��K�IH�Խ�#8?���2X~Xf>�2E�7h��<�]g%==+�����I���R����J%H���u-؋����&Jj�<港e�J�X�jq�6����61�b,�cn���|p7v���8�_+��t����v.i��.~!�a�<6�j��;㖳d���[(jl�����鏩��b��l�����B%ڥ��!吷�&;r�ލ+&���,~�<�X�!��6y����b3���n��ؤ�ސ�߰v53Z ��^�o�t��ْ��wgZ0�.��gv���3�[o��i
����{\j��#�F�w(c�C~��eT쐐��C%xZ�f�mAu>���j�Cnߨ�v��P
q�b�WW���>�k��W�R��������>/�#�7̙q��U���{ji�/^\ �~�����_���9�B�'�??xu��̼L�K-i�a���V���Ts��aģ�~��Wt �8����H��/� �NXI��*z�K�4���}o_7�bUw�㢢��h\�#j�~X=.�ZҢ�ݖ���ݰ���(v}�*3/�������/	"��E0'��6�c�X�����c'���5?���Sd	s���Yj>��e~�،b��A��4f�"����9.�ᐮ�vX�
r�WI�|��<c��='Q�ѐ6f�<���=��3���X�_䕃�N�ӡ�:lmVC'K�3N�L4�-�L&,,,��;:�/DB��=n���S��n���KHM������@FZ�ϛ]���J,<n6���Xr`榸�l�%ѥ���4�����X��c��7�r�Aq�#¥"F�E�Y�DLշ9�����F~`��z:hSU	u7
�QSsbRׯp��yG'@݊���vtT�ͨ�_���;���&�Uq�nOr&	����g+��R9Zs+������d�m�D�7U�$�*)+�����Ω}e "]p�]x{�{��6�����kk'�|^�TVJzbk�W��_����5�79Q�*3��(h��A�˫��9랗��m;Y/޵]�fҙ�>{Ȕ��l��z��e�ZZ��焁����V׎��DR��Ƌ�ˁ�nY99nq�O�06]˓7���Q�,H�M�*�E8�Z�@����77G�����[[kj�T���s���Ԑ�Z/�B�em������s��C1��Z��S#��n�e_�H/��%��1�t)ZFL:�O4���}��X�zŐ�<(�P���[*��%�\[���Q
��#��@HG��=�YJ2i�������5��+%%�5�TLM^G�����G�fW>�T�#��zxof�a��I������G�\�h
�h��&�ж},]Z�Υ�q?	��B�+ .�Cڨ���0&(7>�J�P��VI���� ���z���=��6������y���p&_=�C�@�pE~�J�M����Н������Z\�c�j[>nn����&GgkR�����}���2R'�2# "B��� �&6>��������l�4)[79�x��NEwx���7կ_/w��C̔�	���U���~W[EV��ϙ3���Tcn}w�%%�Yb������be��Q/�́؉�%Xj)�;���y�G�M�>0��||�������Ю����4\\\AoR9H?���?�������aq���9���ZI���*K��F��ҕ����כ	T�q��!�	!m����FFF?���n����褰*�J�5ũq��I�(z`��K������9Þ�9����s9܌����:::�pv1�ǔ��]h3p(ڣ�����T_K�<eB���/��e���R-�P=��9;+�7SO��]9�r�)<�J,
$��p~�Vc�F^^��3�3���?/Un/�E��?r�Ƭo��FPu��8�h�-�JA�����ndz:��IX:_=T����\R3:�Cf66iKK�����>	�P��T]� ��߀&F�GAڸ�E�Oa����a7́�k�
?��w��be �El��	��s��?m�JA��uXq�%A%�ma�I$~xCJW75��J�r��$7ҝ�D�N�4�N�I���X��qp���~�+v������aLF ƫ1^�Q���KsE�I1�I��j����$f.�Æ��q�TZZ*���"-��ȋ�����)-ljd�j8����d}�r�w9cۓ�(dx�u�q����D�{����,>`U�A�� � #�6�WZ��˗/ߪ����� � ��[��Th�khHFA��M/��MF8p���}�����P
�d�%�������-�\p���Wt	�n���_]����{s�#��;UQ�a�j쳵L�Ճٜ��qKJJ(<ѝ����[CM�߾]�?�
���
� k9/�����$$Į������׉����y#�����]`�e�)z4AoRM�5"]7�)	Y�K�7^;v-��}II�&H���	��Ļ�*v��k������%<�Ӎ���;� �1䊆��eA�+q|_H�5t��_ث��t��w�f��ݭ�~�}{��G8���ެ,
䩐����%AɎONr�6ra�负��B@Q������-9�H�+))���q�����K<�W�|f\D�ۣ:��D��x�_�A�9nw��^Y�=�&~w�&������m�j�[��a�(+"��9x�4����4٤�n[-ǵм��^��#/5`YRR�xyyi(������G�����J��� ���g��qQhkE*'��l+�>OeǨ��>}���n�)}ҵk�
~&�]\t���b�b���Ė�;ԏ���׮	X��O�9��+Ϡ�������&�ąVB��O��LL����A�<��p(?�X�s���Qy����7Dd�H�?�B'�wX& Ņ)#��c�VS=��ֶq��Gy^��抝�r 
S�����hM��vq�*�a��;�vBB¸O���ڱό9�ů	��L��sp|�H���	���2�50P76�3��w�����VV'O���@u8��PE�m�ػ�Ra�u�Ŋ�()-���JT���iEcc�?�� �@fǻۋ�6�W+�g^�����jj����W���i��6��Q,�M)��zm��V��r�b�AX{����Ʃ������ܔFLlR^3���_�0����/J2�לQU��a��wz&���G�w�����>�5�_�0�!��y�d�Đ����O����G(��~���YfC�0�s5���YY����Y[��ф���'iy<��U�л���_A~�n��H�>cJ\�C��1�Jv(O�g��,{ێ)�ˋ�?9N�wa�Zڷd8xi�ȀAh|�j��,!�"�Oumm7ww��m�l�Oj������<ϖ�9��o�w�yT6��b����U�È��f��p�yU�����y�G"gT�Rs�N=i3�-3sv�Y��
�3ss��k���nG�=�͞���#ќ0//@�䡸�YKa>���}���r�X,���_��݊�g��r!��_�41Y�A��Օ����_���y�Z�ݭ߽��9"Vl+82�1M"�X�!-8���}�_��׵����������\g9;8Hl�,xWu>�ts�oi�G����aI��KxuĆVX;���u�3;�Y���ڞ�g`�pT�-8Z�G�vD�.S$h���f�m @b�b���3��[����m���Uf� _X��f3Bg`��7Wj��~_	\|�z��~�̓@�;Ȯ�˨�����5����Å�i����Znp��*��\!6�'���H'��u0CW� �O�9(�ku����4�&&1�,{�N/��(͢o��b�UB�%�=�R��|�l���_�w�~_�����$�p0�z�e�E���Ϋ�Q� �#Qh62�%�4ՔVz"��8r鯮ȡ�z��O@<���z����>ɯ������"�"%��TTH����tSs�����w%+j�ql�y�Edb?������r��ZS�_⮟����Գ@�޴�[P,����-?qj�q��A��m��yc�b.���Ӿ_�Q<�a�Ů��V��))����.��>��lW�[^�Cr~��D�7@T,��}����`��WsI2��F5�#�C��$�ŋ�X6�*=7�|�Y0V*.��hw^^_�O�וj�0t%98��5�\��9��-O�:�NY{�����F�6θ1�866�a�nFMWW`%���Tg�$�D�[�f�5�4{��+C	�����R-�	?����z���%�{����`:I�='����I�L�T�����:ۜms[#`CCC=��*��� �>�2RQ���S^�WX��k� X�q
x��ظ�cf�/��k(3ƻUџ�(��Tzɢ�ݱ�e<�z� �z��O��-j+%�.�v���c�T�k�:|�<�(^Տܿ��0���"����p���^0�c��?8|X��Ҿ��͘�=Q8����^� n[�X��>(�,ָb��4�������<�����]W���&
�e��VV/q�YM梀�1i0�]K��/M8�,�D�869��7�E�(��z����G�T����k\���|���j��\{�wH!�w�� f3៿�����ŅB�cbHP)��q?��/�ѥ�ݔ�����xW���w���@ʓ.ȳ(j|�ۓY��'���ߎ��ntS�bR;�9��*Ɋuw��hIM��Yx��lnzu�g<^MR�z&y�pu��ߗ�'�L����򳼽(����[��UZ]��r�6*�v�G�c��K�e��a<�&��U��9���Oƒ�0�T�������s����n��h,��(� �a;M����(>��}�^#� ��Gσƙ�pQ`��׭��؜~��ڼ�	plu��YQ�;��࿪)S��Y�⒐�(%{���8ZY�9���>�ݙ*���M�H06?>����m;����h2�7stՅ��O������~��v����K��Ʀ�7�ܺ�,��bN����4��dD�\8����<fUǹ&�l[1���8a����,!� ��Gj9F��Ue��6ic��dr��s;N����l{X������%��2���	����&���vD�E<]z��0�u�ں�ұX޻�
��|�LW��Y��S�R!Q�t��a,��Ǉ3��5t|��}ǒX�"�p�{(#�EȊ$@9e�C�H�z±��^��Sz.~m>�#!�˨��Y�Й-���m6x��a"�Q�r�Bh��wb�����U�ߵ��B�Ѕ^὆�q@���U��{����Ӵ� 	�u�����4��§��Z��?=c���I�}�?�1��=..��������^�P�@|v�z�{|*���dΕ�D����߸��ɭq466�
��S���T�l��ip=��Cs�`c��Q��1 )�B�Ʃ*9�d����3-��M��9�T���My�CC�.�]�c��ia����}P�o�j�zqݷ�n5>��o�9������R�B�B�t����		����B��蜱�)�����lX�<��� ����H5f�V_�w:`�5r��G9%%���{-u�`��Ǆ<��­6x�wWp��5�k6_#^o+��KF������`��Vo����g ]C�q�����1�<�� ZORP�m&��j?�*��ݎ|�5D�Շ0���`���ŁN:'f�05��f����M*�������SXD��]A܈�����_!KĚdzIo��KA���R�~.j���фX�t$OF��\fG����@�-�u�I�p������||�W��@lc������t.���-��B�j���$�LL�^��-K��S욃%c�B�Q��
��U/��jI��]F����Gˁ�+� �;�R���Wı�+J�=	�EdqҸ�şU%��a�M����{7�sX2Rjk)�3�(ۮ�jSg�%,����~u-_��ЃA˗��}��}y�e���(�<����#�pY��e�s��M��N�mM��"���ܣ�d{�!���w�������H�'r���YD-��҇��;��NMSs���1یp��l��ݧ�Ka�,��N�4�R?��^ј�0���jP�����.Z�Ș�iլ��)��vþ��t�~?�|W��g �|��1-
9y���1�<�b�b9��v��O�f�MQ(_���m<�J�W�зriQj��O��Ed��rtA�8��v��z.�H�}�����C�K�������O�6/Xx0s0O^/�NLX��SB��a�K0*�������o��G��=��[�������b�?Y*p�s�r��mG������+�v���w�Ɲ+���$�f�ۑf����M ����>[|�A�B���RAÝ������v�V3�[��<nC�Nu)��m�rYi���c�:!�&乼`����W�+���C���y*p�A#-m>1ȶ����U��}0�+	�u3ː�d�����@ގ�sI�i�1������������+��^��f��}G����ZZ����P�K��wTBn`�MA�Gݝ�Z��]�����q
��ɓ��Hv����c���l�b_ڬ��:�����|n�嵯5bC�D�W�%�x�M����*p]I'u��g�**y�a/�����Z�����0��In�ž��t$ddմy�OQCV�5�P�Oֺ�t�ŋ�<w{�gl����5�,��&��@ )�
4�k�����{r���H cSE&_|k3pG�89+It#�{upYQQ_�gG����e�Le�h�i�c#��eF�D��K6L�ȣ?�Һ�~�[<��~-`"1l5b�~P�&�mkU�hg�g�S �2SSOq��$8n�2�v��x�⿬��`\�щ�$3A�t���3�	-
�a$��׹�������[9�<Z_�(����:X��[@�_�馕�}ɽԸ�5��Er�t>�ut�p��NNN>21�8纒��T}�F�)C��C��\�0��Q�%���Z�� H�W-L4ekeJ��2P&7�EH�4�#����a����>��ɬ��*�U�&�)�����8�
���{$mQQR�tozJ��9�"*�kI^U{�:�aB!�a�p/D�r+�=3���Ǖ����3�^����,�>���$`�M��b����+���T+__n>K��� �*a"�H���gAK��c�1�9X��雒�@8�Vuҗ��m�hjk���&d�ƈG����&ߊ���^��HF�ފo0kKR�W�޽��8����IM��WWD�EQt�?�������%��l�͍_�qkFK�<QOO�^�{��x�wKxn�#�/eIi'�y��ϱyN͌���B���	�j�ͥ�������*M�^-��N�|�rk�@�Әm���UK[��W����Ι���a������[� %��4�c��H�*�J�vU�5���hw7�,ȡ����ܜ|����U����罎(<�!ф�^{Ur	t�چ�o��)� �£�K�����mkD~���i���x�ﶷ�f��'��fM�������LJ^g��ࠢ�j[�\\�vjJ�9��w+��V�WU�D�Pӆo����������{��I3��f-��+�w&��L�IH���xYՕ1�?�|3�5��G�s!6��}Վ���0v��q��ꚭ�8����l�q��n�ZR���Ũ�<��I&܍�_vm��R�]5)T���*��ۜ���<h��s��{{\��G7��4�ex5���C��93j�m��/�����)��9��T&��ʐ�M��e����{)�As�]�Z!az�VRb>Um	��2�<��O+��2�G�������5�y`���u�%�U�$E�䜜��U�(j��$�ɐ4�K����K폂��`t��l�w�R�
\��x���i���J�#c��s�@W��!W�֓Ehy\��F�8(�6,�E2�Wrf�C��c���y#�)l��&/؋[ZD���>�Ge�^M[��b��r�E%(�R��Dc� ��]���b�K~x����S��� *�	�$Q�㱢R�s�p[{����R�ŋ�%$��.}zf���A��sGsN���Y�E��& ff�2�(���rߵ�f����y�n��?�߅��/��5�NqI��g�'��o� {{{���2�3�T*�^�y���%8���hZ��5�V�l�RQ�#�Gm`� k}�N����{h�j�׫y�\��5z�Q;泐'a��-�yT�TUፏ����ͼ=�:^#���
����*g�g)�S�oon
� ��l��`��M_�����
"Hwww�,��%��!����]��-�J#���{��}r]�Ù繟;�������]�wJp{��!~0�{a6`�0���m���q�H;s����x��6�_r�Md�ah�8FGE)����qTU�(.�wYm�����k\�ap۸]���9�{�+&�7f���5�h����i����,)�ۋ^k��R����i���NX$g����	�!��m�^��c�1��}dw~�zdOV��RHH�U�I��88�MM�)m�T} ��>ݼ��s~�>=�mњ���_׈���"��:�S���	�� �Ư�߳�����:�/�c���$���U�Yq���!�Җ)d����%4l7[e���u������@��ڑC&NwC�]LLLK����hn��7��B8cbv혙�k�{
������v��V�xQ�9	P�>�R;�?8`A�E�	�hv�'��(�5nw5j>��HK&�(2�[Ո�bLZ�l}m�MC�KR�(�� 3�b?���l o�Y�BS��K�7�����nN�U\�= �ӿ=��K�2�#?���:[,JkcuތP��f�tj�m���.�yz�!e;ꙃ�K}����j�zt������%�Z������N\\(�g0���.��h�8ت8(I�����C�6���0�3��b�y��J5�"�2{�
M4�("9rOScdd��s��n6�w���V
�)���%D�Y����kd�>`�Y����s�*U�2<�#��B��@�d$q��^�i��ʥ�����h��E�	�Vm�N>���@�%,,J�-�@���D�j���|�0{�>C�O"��gd�y�O�\	��;�������e4N9��21q�v��G����-{C��/m��������Q.��Y`u�x�Ӵ�(��o�h&���cc��|�3��Zg�ߋ��̤W����Fk3�
�|ii�𝽎��Q�[X 0F{��	-/���֩jڐ��6f�b�n76y0癫'����-YQ�����8�1�%���0���t�)0�ɾ�0R��חd�f��F��c�5�����]��/���C�fs~PI����?w�w�(Oۙ�ꡩ�}}�ł�� ������ɤb�H?'D�|��(�Sn��*3��q��Yc�#2*/|��Ѭ�tAj!��#�2��ɰ�_F��D��;�)�u�RQE_os*0�:jf�%��%]9��p��۷px<�3�����&C����ݡ�'����L���/���[���wx�G�]lN.��j&s`q"�|�l��h�5�-�^��,��t.f�K��֝�N��.f�`��<zzz���Pqqx>�������r���s��M�Ge�Mj�����v�� |yݧ�_i�6�ڐ����[��e6�L'*��b�~��9$N�ع�0Ѐ��Wf�
���U|�n���`�P�o�-
�R��x�Ƚl᷊V��z�G��g�
��G�Hn}/n�V���5N)�s���|D����׷&�{e���T��% :�������D�`����L���)HSJ��&��4-ߘ$Qo��>N�Ih�Po༶_k�~��ۃ�~2X${8,_������,�a{rv(��?bAu���a��.�~[��(V-�����RR��^�ݥ 9��QE�=�H�8m�CЏ�=�g�?�΄w�#455�(i��3Оɧ2���\o�;�e��K�)�ZS�h���(}����9f`�����0���b�e��v��L~ssj5}kF!�N�;�]��a$�Of�r�T�ukE�8j���TI�������>��N��y���
ו}��V�fW0���e��/O��9~���������(КU�Sk�Xg�H]f�d� �?�k����7�g`=�f$��Ņh�R<_o��m4=ž�c���>���do�\�3Q�+W§]�����Z�h1�SX@K�ꁛz��\�`�!={���>e�. -������5�����p��c��b&�s; �aaa{]Pă�Pg��o_�i�G�_\�z���Ej<� �a�.�<}p�A���ѵ��;�5ѭo��b��^V�'��!N�) �1�,��U�z/;��4��7
o����{��s�؝��ۯ�*�w/���E���c'M��w����m{�킞�&5���Kq��Y/�ئf��J�֜�c��N��m*o֘�[f��BRRZ'���A�z���G�j]�v�ج�B�o�ߒ�>��pqŷ|�geRi�{#]��|���tٖCB�rLŋ�'U�W(�x�5�~�x@��3`^�����@�Fܺ�s9��Ѐq'�3�\jcMEp���׆��S�`�t:S���P4��Q�?;B�3�@ǡ��� b�x�DRD�����]�����Bؤ����m����5�=�n*��3�g3QIUdU㑒�Pf�λ�n0����F�_R�Zme{�dz����Q��J����!MD(ۑ���D <��� H��&�=��_���zEȴL���嬍��5�����h᪠����$�:�#��Q�Ph�������C���{@�U+̓pD2�^����v̝���V����Su$�/냜�sT��8u�~�8�:�L�L�[,Qr�	5��8rL�ʁ�R~K4�fZ�;��Vٺ?�����w*���&k�ח��*��b��'�,�e��i;�bBaK�л�Ku=��I���S�lI�<l��k�TD�%2fO8�+�-y��Xە����G���,4.f��ei,C�v������H��v�5j
_�e��x��Ec��100x��z�	>w~��WDh�5	N�7�i���#��lrZ�����B�FVG�ߥ�lpqp'W~�E�0S�1�wZ�lcpA�'\|>=,��������h|��膻����뚃�j�)!8̿�6���Z��
*��'��7���L�>�߁=�?9��]F/�i��k_])���1�qk[[
�L�v�"������9>�<�݇^���i�������l��$�UID�րO&�;��b��B=�MMM����D��0v����e���c��h�'����:�3��5z�h]���U�:�V��&k�p�,����*+��<+qs/���#A㛰�C�w�uŏh�k>��H�x��?���r�quu����;�<�t�:P������%��7WC&q+s��VC*���3��k+�PUi�)��9���v�����"�ƃ�݆�i���2�f����~u$�m�\̺�;?��~K����µ�y؏�:p��H����QuO������j<|z��L��_���륍�6��R���r����D�!v=滠��ۯe�g�2F|�h��̾y��))&���RY""�^��HQ(ss�M�#vr�泇����FU�������p�<Y�AVG����g�a�Z���\�$��,�F�E�%�;�o�6:���o��SXU�����~��Q�?�p�����O��?B��D��7���-�*�x��M6{�����a�����a�������*����N�E^�;�>d��p2a�F}j[/c�&���<::*���>2�@����P1�+�ˢ4�q�d_밂�"��R�3��pV�E`.�&):�
����b�w�������8�`�H�/�����)���Qs.���G:�J��
;��4���B6��i����0	*Bv����r��۴�M��K����--�+l�-x�Y���
 b]�-���7���t0��=�n����>���PAa�3j�EN�h���?��tN����s����{�����u9yy�M8L75�Cob�x��BMw9���/�G��1p�K�b�2#�>>VS��ǭ	���r���SRz36�}h�7��v8�+��A����|�t�ds=�Ã䳾�H⟡���������l��Ќ.k�6TTD�[q��<j��,[9t�u$�CC�3q��Y����8��v�)��P�˰��OY�4ޱ�v��VVʍI��i���tǢ_3���Q�u�^2M7�Dyxx�_bnFM����ң>��}��vkz�|�
 ,�-͔�ZQmou��oUIS���E�?}_.C�t�7D$��˲��W�dw�ӭ� ���S [�mr)Nz�^	�gV;���U��}�sl����(�zA��� o�Po�P�k�A��������Xe��S岍����Y�0k�qdˎ�c���1� Z���5ǡ�k��u�x�#nE;��aC�~�(&|�K#-m*�#�_���r�����WvS9� �	eJ�M����E�)�MMb����s����H.�;s#����y$^q�@�9�
r7��ꍘp(7�t]q�v9wS�4��mث��Tw���%\eT�5��%��o>�?��.s�-rPC3�F[Vzѐ�˄7��kb�\Q����ؘ}�ԛ-g<�B���"�^\��Cso�|�4(b ^ݰ���jT����"4��Ν�&��g�+h�D�%�"pD�<�L��]S2ҹT�H����H�7�vy��*�H�㤊�]9oP�`�5ȍR�����Ҩ>f�.3�3���6� I�^Tқ-C�e:�<�(pz ��{Q�8g�ۈ�h���uPa�r=�9`YX�7����g�xW��:��R�eB���=����j+�z�HN��\~��>���L� 䰸��s����9��0���M�P��`B�r�ʶai0	Y��W)�#*#��D���Iʓ�<�W�9�5Ct�'��;k����;;����vhx�pm�@LV�C���<���
��blP~�}Ž����{l,��0���Չnm�V?�ƪ��R�zZ��!�T4�Va��j6��E����g���_ODNv{�t�S����zQ�g,�.�!A��U��e��5j�+F�Mޚ@����8��\���	1 �u��:��|�S��ad�wۏN&C�*^�4�b,��@�v�ȝi�ڌ"e�ͅ/���ȱ1��%���l�n��0k/;Ftd�5��%①�=��-��|�jȽ����j厃�z	��x�����
�e��\����Tfn��US�:A:J�(��:~��D 7�N��-���2ω��T�N��D8]O"	10Q�b��~{�EK��(W2�!���U�����_�%g����P�~_����w8o�FM��ޕk�������9�y�*K�n/�����<�6|���_��ϯ	�	��-� �~�p[
y�5�;%��Q�*CRx�g��?���	.}?�`�6��Oo���̺1b�J�x9�6N�	[��lTYn�5�-k�� F��_�+���@8�k_���p��n�Ø����KM!͡���K��⚦%�H���K�4|�.Y��,ML�;�jQ��2*�d�e[�L41�hj�`l�.1,'���4zl�ÿ�i�sP�!��6?o���p���5z����1n�4B��j��۫!@o
Mk<r��Y��6�陘��=�5/�mX��w\l�I��EeJ��픘J9��[�m�DP��O�-�����ts���핟i�(Ù$I8-v�l���{5T&�P
��"]v������9n�^�F)&���?+�G��?X]!�>��Vi���k�̢�B�edD>ή2$ ��$��-K��1�j����{#g�Kj���ʅ��LRS�7m�x~�c� �IՓ�6N&�sp�(B�(T��>��Rn?L���xG����65��7��bO��Bg�	�m~"n)b��|%�DDȸ�܁�,9՟G6��׶����	2`%���m-^�F�qn	�����'q�l��~�lE����!�.Y�2���pYn壩y�����x�䚈��	3I[ق�?(�)C�+��6�
Kc�U������oz���Դ~����x�4a�sŊ��E���0K>"�ҩE�:!�T�� ��T�{j>�z������M�{�_��	��ȠG0�AP22"�cs.h�s
�<1Td�Cl�#?6��+�1y�[ݓ�~��}���1�y��UOf]���W����>���W�G,k�C�Լ��.)<�s�B?X��<�e�H�4 ���FF����� O���X�0v���b�8�]�M�/UW�����o�j�7^}�K۪�\ZQ�{Kh�p����Uu��'�2�mzkL]G�Ӹ��m�D��d ��*�䏗^��S�����&`��Y�����i���<9,�>0����F)�]����mSI��k��m����m�L���dcg���@O�P(k@��� ���;W&��ݡO�9��ECz���Y���F��A^�k���z�U0J�?����6NvQ������M�b7�@L��+.�3����m�ђtҸ�㺦$<�SEtf�FpDU6�v�l*���e��-.����,�J�dPy,�h�Թ��k_N\�=&k�3�W9�χ���W�Bh�CWސ����3)����S�FoCKQ0�ǙgG��Ŧ���KJ��v�f�544�<�&�@�s{���NΦa��ww���1@tYc�	��yK�W�8]M��]� �tFlB]_x�A�[ʄ��m��px7�<��#��ɱ�X!n�Q%j���e���,b���dz�sA��ؗ1��|Rr��������O���1w��Pm�>n
�@�P�;"Ƣ��K�O�n%bۙ�?��\;s� �=��w�4���cat~�v�0X��C9�~�*�cN��ۢ�����b?��F�ֆ[s��z�X\ۧj �@уѢ�ބ��ޮ�o<����������=zbTpK̵�gϙc|\bK���(�W4]�ܥ%�NȪ��.t��&h/|�����q�\���%�}�.K{�۩)�����̪H���)��ǀ��]7r;m�t'jw��\f�u�`27�u�#��_"�&W��p�.�);���P~;Wm���U=HM7�l��GLl�Hђ�����v�n?'r�U�X��6��V��}9�Fkc����j�.ښ�+{Δ�w/�}$�;�����]x�����OK��]<6�
���8Aniw�m��0���8�f3��L���N���Sj��]b��Pl�6��g�L[z��u>��n���!=eXM�x
}���ଢ�Xe{k������z��&�D���c&]�^����f����n]������@���U��c����$�*�H��7�.n�,}�ē`�Ɣ}'��� �'M��9��= b1c��ym��K�*�ۓ	kgU�໥V�j[H�
v��+4�X����Z6)&�י�B1���)�m�7�y��Ŧ�e���_�=�j��v��P��y��UȽʹ?����3��*'[�IJ�]=^ǚ<E�U���Ԉ��=Fߔ�K���\������4���o�?��U�݈�[�E\��0�_�`��jEۘ����:�M0���"���n�@�)3�y4�����]�{M��^Eg]]]�馔��>��"�8D���۷k����_c����W>���ר���p����l������Հ(��ґ�k�%�O��(�"g���tt�
�%�}�y���>���\sv����X���*�@WĹ\�\{�Kɩ�bR��*(�rwoUcMO@鴦E�:���޷c���n��d�0��W��To[�-��V�kO�m��a_F���ϰ���Z���?,#��-�� ���8�̗=_6�ٱ}���t��;���+GGl*�N%�u�\r�A���Q����ݩyyN�t��Jδ"�
$�C�W�|�1IP�׽=����-�3�_�Ҵ���]Δ�d��4!�?�$V^iRʎsK�U�sy�hS�������mQ��)??��ɜ�G�V�̬��Z����}�,
SU�!�4�t�7�\j8D'ֵ�������iZà�S�
4(���onX���X���L��{�c��׷_Z�cG����&�'SDt���oM)��TA�1�&��B�����I?N��ޚ+���N\K!RF{M�:bviP�~��b��"�W����&��Ɓ�*׾�+S�簊0!����]hh���9A>�%5��zFh�Ju�ࠣ��3H��&%޹:��(.މ9��9�((qlĦM���2V��H���週�?�]��]5��x�R����o>a����5�]u|�uZLI��A����b`�{�&x�9�zjc�MW��J�F969I��ʹƔ^����Q.�t��I���I�W��	��p(M���T�� Z���m�4S0R�M6�U��y��;4#b�T�v�g,}���?�ih�m���!�-�����m����4��v7Ŵ(���8k0hy�z�z��U�<��fl�r�N����m1D kH��4��{)����v%��\r,һj-��4��l�>����]6dG�3��&�G�ݛ%P�N%�t��)}����"@e�O�o���ܭaΰ܀:E�E4ꅻ!�����<�S+���N����d.�^����W�a��C!f-�q�Pߒ��ʑ�i������D���������Ke(6n�:u-"H��� -M٠�#.Ȍ�߃�n��"�y�w��rX�����$}�QlNV�ӯ)�&��b�9lĹ��͓�ѡ��>�nJ����Jk�%�>`�|����#�k�����0�^�7�4Gc���n�f��ף ��>n�����
r{�P�R�n���1_}{=y���l`G�&�\�4�l�e��*��	�H!pړ�3	���4f��x'<�;���m��X�S>��։(U���l(\b�7�05������.�p]�����x\�Zz�&j*�j��a�ɑE�|Ä��#e���{f^�E�YUC�׏�xq�Q.��s&Bo�����hÈ��=`��gff� x<�9�r�E&3ͣ'Q׳�X���RF�~�b�??`��8�F&��>�[���-��;o�
Z�c�m��m��m#D%itW�s�C��7�O��P0���ѓ��M�5j�8H$������(**�g���'���S���I� �#�Ine�r�/�fZb�t7<M�TUE�Q�I�1竩�[����:��XhS���YE��O����9'�4'��+bAW�~�*��T
��Sn�i�5ay�(�]�6��}��0�����hx�4��.����L�X��� �^�[�拐޽��:�����ϟ�2>*q�%��zz�b��4�ѡ�$���ܝL��S �y�,��W��N�w���ƯA����)B�>B$6��K_sI)L�ٽ��6�G���*�ga�3hQG��s�֑�.�����	�?���ҕ���}��*Q�|u�N�+��FT�B�'rt��%���b�A�ovp4.�w���6-5���V"�^���+���y\,���N��O�<*8�ǻ�'�WA�������'z���n��}R[�f�Q
~4mcG ༰��XG�U٬,/�#Ϝ(���?�`4���1/N>V���!���)����k ϳ����F��-ボ�=VH?�ѻ0CP�MS�M5���rN���<\y����\?��9j�ޅnO@�k?�2h5�RR�R��+D� �<#c�i�x�_�a�}�
��=��:;����Ι�N�r����}A�;3ӗ;���x�A%$�)��T~�'#p�`1��!��4�����H�+�m;�@EK��0��z��!-�N��E�^��~�m���eiCF�ǵA��5ǧ8���%�/���U�g�XrK����SЕ��~�����9�^��~Kv�!ں�Y똘� +N_J��`����& P[G׵8�8��+��!�/�g����.�����c��x��^;�\�.�M=�&��U��j��6�I��w��]��3>�;GG%�i".rB��?��y�?���8����������B�^�䮜���}ݩo�S"�-aD�.���xiD�u#��}�t%fj��E�w6Ǥ��vC�e�����>%S	��Q-�}��� 4���=̦�&��#E�GOo!ff���%��yd}$$�d�a�	��WSS+>�����z$��Mz۳C�Q�[��6
��>t<��r���:zT�=
~~|]]����K��#�*=�����z�^����~�,3g�5���љ��������#'-a�ϰ=4g͚�1�f���JO�RT'�uu�nmQQ�;9=mfb�l�eT|j
?ˌ�-��Zg�,��5�MѰb����������Ŷ�\���'�z(�B�=��U�\'^��a�G'4L��CJJ��h��%��4V��)#�o͕�����r��_��{|���R�j�y�M��,��=�@}���Q�_�K�آR��6sg��A~كD�*��{m�٠�_�ib�����w�PD������_�Uڵ�pp�����_o�p���;~JW��� V3̎���*���:�NLJ��q��r�=�ӿZA��?H[O�VJ`��}l�[B"T-�Q����������̬���q�-�"u`�y}}�	i�����4jH�E��9G�<�6���
�������L���D�D�ĕ��闚���m�-�y��^ȑ}��������ǹ-y6��;��}�U}������=�q�TT�����Z�1�3�=ηo�W���***��8�*�:�{݂e��,��V�19��.�����{^�̲\ke%���9���K�Z�R...%=�htrjȑ�$w}��R��sOɖ��>�cJ_������D���!�bN;Q�!���2;$|DfY�^�볻�yˊ��Q���@���}5#�����B�R�༥%ƣ��y+�dZqDī��",h~��r0�&����@ꮻ���\E�9++kؚ#/e	6�@e�g<'�;(����L^S�h�g:5��I��"�z���c�����ׯ_'$&�J��:��K�)*Q,�	/�8��K���}ww�<�[G_�c����t�<�Oٹ7�HoG���p�6�ϴ��C�K�����==y8884�/|�����<�Ҿ"��%1.|�J���HO�Wq�OB⋫�˹�S=�35-�R4����ƒ������~l�1��auu�������~�Ϥ�z�6$^��ƙPF!/%��!P<RR^�􊷲�(��� O�'�ir�O<B��|��枭�����!k��`�II2�������ZXA
r>=���1����۱ �!�fM�
޺�Kǘ��/U}yxBU�̡<C��^%�r����;l��������III�n�(����t?�E�)
���k�q	��?$��1G�(@OT�;LQC�M\^^�y��MEM�cp�sL=�J7��R����`����4;�g6f�?��ЗO<�SR*R��������/�����@u��t`��1u����.҄��%z�q[f���[W��Q����6����z�Ij�˃�Mr��q���?�a6�SD�F"Hj��2��Kv�����r��os����=����Ҳ2���ǝ$�E��HQ'�4��rzF����gWyG�S^E�Q�N#'����?V���M��І�*At���_O���z��$��HffS��|�r7xH�ʫ��0���ޫ[��WA�7,w��4�=h��jV/u��Z_͏��B��<;���זz�p!�"B��m*::�P)FJ<d�i�(��p$�Et��d\㓐��)�--+So�:���~��ax�)�5���v���,����^���V�=<Mӳ�8�	w,�����e�4�[V�HAw?���#HG������g}+)9R��.ATֈ��NН�[�i+ ��V�����mRҀ?&{�!�8H!$��qH��k+�FSW��c/�DC�(�/��Q��<�J���] ȭX�p�Xp�in�*�R���;����԰d��)L�*9n�'�#��'?�*� �Y<����,��I6���U%ϦÈ(&T�>+MX[ė@�9���Y��WNjx�t��}� �o��Q�&V���]��]((��C����ݾ�#�W�<C���_̀�.�>��BY���m�@F/��Jx��VsXT䬨������^���eŨeG�6{G�f�c�
iUmma���[�Zs�5o!zz����鉉wF�����
[������ש991���+K� �)jzec����,�1�W��N�o�+|�<@�֑�dL��&^^��)��tY<H�7�{{���3��\�9�!!!���8 HI7�)g�J����U�����`����V������:3�6�(�xqF�K��3�TUQ1FQ��6Q��迻��??���	}����VN67C,��r��A^��/|^�S�+ ����6<;3cz�Lk��5���B�"Ґ{HG���a���������ZV��×dz���rf԰����X���a�'�k�KKK��~6�{�"�����Pt��p{��X��㸊w��a;�b���4��XT� ��ZΠ�����V0�����xƢ���}CR�����`�x�U�5{�T�����n�6�I�ݢT��Zfvv5�������S-�1N�z<����0�������Y5�k��S����
�����w<;1{�w�o0�---7o<.L%iM ��2t.���ބ���x��� ��d�MTTUɣC���Cj����YY���S���XR9ق�Kj�lG��Y�M�kfE
_�R�q�QЪ<`m;����a�eͲ�ﳷ��LL�Fl}PPPM_t���}�`@W��*�����"�	��ַ�>P��/ U��B�aԀ�M��䤉���1���8���	6��a�,u�����aO��J+N6����D�<J�ڿ.[����ԁ/>�V�עƾ��?�8�� ֕X �"����y�����i ��x���l�RU- ����%�;95OV��J�?��>\�h�gVVT��Pw�m���|�̠~+GϥX���ߟ��=�ǁ��j�yr�@d�6�z�F��ّaRu^�,,R0�Mώ���t����zG��������H�+cy%��?�����P\V�lE�N���X�vEEMflYzR �E�O�tX��"i�����12r�W�`�<����V�O��]Jq�p?VW3ihi1,�=�l�R�|ka0�����f.nQy�Hp�����\��/����GB�麱�<�����@@Iep�glY�{ ���xs��mڸ��L؟(����S��Kv#e�D+���+q��wy������[�,@�,���b+���<x �ZKFN����f~�)~��R���J���ү�H+Ů��W�e�v�xui����1��.Խ��w�׷C�*��K�6�4���`����C�/� �&ef,d���,K��_���LN���;J߽Xx/�d���'�¸��s4�B�)ρI�g���J��g��(>RH�o�./�u.0Ov\�~pA�ζ������HC��/� �޼C+���q���ݥ&&&V�R�}dv�e����Fމ3�ы|�Ʉ�����-C�
�A�$�_D�[��Ha�>���,����IK��K��ɗ> ���8��xK�+���W�Z��p�		ś%��"�Me-��L燤���h��p�|��LA�8nN�ț���}����+���6&]|�8q}@�᱄� �H�~�Z���3 �_?l�G��'���q�VF�r#���fO`�F9+9�
�z��-�Ŭ����S��1J:�jcVvvv��;	���8�N��o�����Z�R�)��Sۛ(ǹ����apЎ-<*j�Y�]�o���Ʌ�+'JM���Ͼ�<g=E0�SQ��cł� �A����众<�k��R+���	����6�o��x���#	d�����s`�S=�Z��&&�{������X��a��	��׿�g����V1 ����O�z��[�����F�و�5섺�Ȃ��"X��m�b�bq�ƹ�P���������13��%Ď�L�-Y�.>Ś���6)��C��9GDD,5�i'D,����s�gga��NE�Z7J>��"����=W��t8�I��U�2���C�[)�Y�j���̆cev�`'Oâ:~�6��j`��MMHK���RPv6�Y��%�J���2j�^\�TN�˗�����o\������ �e�ms�䝕��	a��ƅ��1ܹ���w�ܜ��J3�e�xpԜl�����>�B�X��J��M�MH�37߭ �/������,�Z�%��<��lB7��K%%�Ž}k}�?)�f��FD�8y�O��77��8$�Z��({IC��^�D�H��^��>����˗/%,o��j����4��@ꤚbX�ٕ�ݜ^�Ե��F�O�.r%7�|�9��x��ͪx����ذ0��b�#�w��eHH�84�����~�BCff��/��9E��0%G��6�aa�#CDv�b�P�{Do���p�ss�Yoyv�A	!��\]/��:ҋ�G��ⱥ{HA�̩t�EC|gn>l?Q��� �XFN�^���0��&CI�TNT���E�N�xH������Z[5# 4j��V���w��Fp������q�V$��b�FF�W�pQ�������Re��˺׻���ߑL?� ��0����Ob�R �6;�T��Q���������(:R����Ng����.:Zd%wW �PMOeƣ��3G�_T��"ԸdX#lzt�q_��57{f%_��kÞ��(u�Z������t�P��˥�_wITտ��B^
QQљKǰ���~T��,+�4�H���Z=e�ީ���dsw[FKOO33��VۏT�Th�v(��Z5_��yk�[YIߏg�vjkk[�YV��*��v����+�}_�B?~����Y���[q�=%�0�C�п���IL,4HS�?��WV��v�ڶ9�����,-�٭��=�g��o��}��XL��� �������b��w/ O�$�u�4����6�����G(�I�RQ9{�fg'�8dϭ�/&�\W���>�N��#��5;���8B#`nn������L��Q�m��0ݗe�|@�������|�
���&̞���"�z�m&DA���^u�0О���cF>���V�goP��}����a������҂�@�Z��������F]r����%�;JM��=h5���`���in.a? φ'��M����	F�5o����|��*Z��К�2i\LX���NRh���|��o1))IԽc�>��0K��2�ּ����%�
z�-hA|C�T�1�&&������u qJi/t���_\�\��>�O�:�3�����
�m��[ ��*�?8\��#�q�1��k%=�3�D�"Ki�`�e.;��AXX0LݖTRz�y��E�,�!eOs]�s5 xm����g���h�����Դ��w�XS��2�2i���v�)�ZD��W�ejY�v;P�aȚ��D�������S'����
P	;īr!)1����a*�Y�3�|}���� m}I��vg��0X}m8��bv{�62:�Z���s۳㩾�{=[`�)^���R����l�{_�p}�������ӧv���F��J��#ww�W}�?�(j��'�F�m����k��N�q�왷��nὂ��ͯ��9�j�7oLML�pkEJ71�i�3��񮳜��1߿��i��l5���q}�~��+��0���1��ه���㨜���6��?�5]7�|�p����((A����1!���~��x.�
���\����Lq�����Bzp9a����D�w=�n�L̡��LpSp��o���C�Y����3�966F�7����laa����	�z�j;Hx�a�\]ծ��zZgz�<<<"ݔ
����׍�[�n����\t2�`�T���:�+ڸ��歞C>��W��Yf-�G�e�����&).�{@�ru0�x{HG����zwS����!=�d!P�O��k����ߪ��K�g�7�V �� �G4f!�*,���#)���jYE���!�ñ�5|#a��{ߔwx�IA��&���<Ѐ`I{FGVSW@<���Z�V^�YC_�3��]ǌL�-�9�dL�w�dw��mP����*nn�5OB��8>8��/; s$;��O�o|���6�!ǚy��w����9�������������
{�§7��/�ol8Ay�1�� =�-��u�|s�]|PF��n F�	X��S׶��'\��c&�/�
�9�
�E�M�8�ӷ�����EL����~�aO%�t�������ҧ?��q��'��� �]㦼sԙL�%�g�"��J�(�ư���CX duu�D�fx-0�):��:��y��T��l��#Q<�������j� A~���C!������(("_�rr�99~e�嵂J�����w����!A�V�� �a�	�����Y���B�O���J���2ܜ��P���C<I�b1�{OQ�Sx���F� '&D^N�C�Z��g{+M��%�N0�:::2=�^)aO�o\�̇d�U���į�.Bj�1�v�k����_���U���l�HS��KU������"`�$I߳���2��h����X����v ����b�˯�b�"..�q���&��r-��WWW�ޝ\"j�=��z��lP�[�l���]x�8�;���8~��QD�p���/����@���
pp<�٨�r��F�<�x�l��~��XSSS^�f�Ź "�W��N�>#%!!/y<�$S������ü�H�?�T�cb����@��q��~;�:�=�ӁW��2U\�ķ^��El�ۛ��� #z�-��ls����l����U�K���]1��v{�oE�������E!������0;���j�3sL֧j�7 ����������� ��t�T���q���I����CIq6 �w�:|#��Ͽ��Q��4lie��vŐ�/�i��f,��;�����muuu<||1�fe32YYQ�nOG�hS�JY�S�D�}	���g�WQQ�c�:n������SԁlC)�ǡ}�r ��������by�����t�U��ƃ�?KKx4��	���j��LL��J��������}����!����t(�   � �?iiA:�����n8��y���k���s�>�]{���u��Yw��c�y3'O�K�]+)���&��M�uS-�g�xE�{��n����a<b���2g˗�c07?O�U^Qa�fxǣ�Y�8����F_�A'�}��ְ(e�W�s8�b���׺�4qW'�S����8g�p���h|A	#�폾��CLN���}dt:&�!5�?���E�6'��?H^N���I�(����o�Ů��O��������q	��M������MC0I5��Yd�yb�
���r�vJ-9e�>F�	����pvO|E�!? H����eAr\��[mں,�X���������M���V �1iE(��*ɥgmU� �}��K�W0z������@)��p��B8�����n�Re��[/A9��g(n�);�;��'g��p���Ri�����ڎ���G�Z$��(51Y����^#����&4�H:�"�t&uȨE�����׽5w�Va' ����i�C��F�9��3P.��tt<���RQQ5����hڭZ'����;�wV��a�$M��|�:0���=`�ye���	����%D�oC���1c?5CZ����F����S�X�:�����1iI?~0Y��������;L�Aߩ<=�i��,��	�)V`L"��gn��vw��U44�9�o�Ian� �p�,���/,L�:W�	oUUU�r')5�H�/=c��j�f9�g��Bp0!a��O�*0��*�d0A �-/C{��!�?l澴�8A$"@��ɭ�'##�u�E�����ôؿ��M$-����W��swq���jw'�y���2qnjK33��R4"�T���W�^5��h���S������kq��ݢ�d�+v=T��_X��e��q��G*�+nd��(f5���3���~(77N����obB�D��oo�Ű3�ǌ��(r��a�E�����z�&���r�.�O@�+�48Y�9�S�>�S/.�`�5����������w���h�a��{��P�&:Pmq:�]�PS�Tد�����=���,�=�O�.#u���k麪v�4C�mݯ?�g������),,9+�N�Q�6:6V�2��&��GW�V2���)F�t���l~�"��-P��GFj�H)�牗5)����Bӄ�����^��plx8���c�H����rM��~�s`2�,j�l�w�9���g�@�i���~蛝͢!`lO8��.%F����P�u�^vc�Y�T�ggg�,��*c*�ٌ��"��X.B�
TD���
(SZ�X
m�"I=����%{�:,a���11o�÷�Z���o�4DDP�h�$''�z�(�H<��QqY���8o&��K<@S�N$�����n5j^�TRB������^�U@�F�%c?n�<c��e``���Nܑ�2��]ݔ+B���je;=}����l�����]I��(�bb��hvW7j��A�������`�����D|���)8s^ ��AY�Ԃ�#t��g�>&.F'����ØrC�ߋ��x�����`s���LJ��|����� �ה�ǃ>�;1\]]�JʍZ������P2�����G	er���|�QC*��I��L�F������ٷ�\�طo߆��`-�����v�ٸ����u���e�|[��kc��3�e#��vu0����F��@ws�ji}]tqa!��'e�I�-�
*��@�}��uj!�B�@���S�����@��uv���zt'Vy�Q�o�� ���s4����K�hWW�6�5�CDW�7��Z�]�P��_W�_�gd���C1H{��U~�����;|||]��>aN�����ۃX��DL��eq�f�H{2�i`������z%�X���ۄ�c�c������,��� �׿׵z��f��XH���62*���뛭ܪm���l�V��Ņ\(�z��3L��|���E�%����=�o�y��9͚�< ��H+��R�q�����NU��<��V�i����������Vg6P��1z�oV�Y�ە��;H�]S��p�WOW����>���M�::�#��l<<��U��j^7Ťu�p�	b��I��}n�Ui��>h"�
s���!��Va��IH���R����$;�n.|:>�@�c��.&f��(�ud#@f���dea�����R7Kv�F��RssT�-��7UL�B���v�z�]���9�<���	�B�׽���*�h@_5�����`�y�=*1QT,ՎO�@��/U�c��I'���8����/��sǓ�|�YE����w��5Z�׈�M�դ��ԣ�4s �nxP3�xS7pz<C|W>C�CVK*�/�(�F+��)�9;P�j��Z.h�Ĥ1T��uwY{q���x�]ה"�������������j����!�Ӹ�z��S���=�ؔ!�bRNM�)�{�!��8w�^T��^��]K�ح��e���R��׊���$��Q\�7�8 'Ν�zbk���i�yR#��y�Bg�����Ɔ�.����J3l����r>��r�C���[���M��Re�L�����"���կ��ܱJ?^���D^�����=%b�ؐ���(��k����Y�>�����Q�VJV�	��R[{{�A�*iu�C����["��.�W��>nN=k��j�٘!�C�I�u>�P�L�߳3��{�9�>����(e2�������r2%�'�7��ۭ`�|�oA�������Zß=9��P�st�I�O I0�i��F�.`X���p��Zl$�&a��pOF���>�!Ad���	��~�j,����X��=1;Қo�
FJPY�a�qE�����A����5tt���� �m�)��<6�£��K��$��5T�����u!�\]E?_#s�]���;�Ce��F
��a����/�V��,mlT'�R2��VD~g*�|�����1�;�ɼ3)bb�F���x_�Wo�d|'1,1�fbc�cٸ����-;[�RW<�Ou���ӓ2|��\�Gn/�N���YD0�B�b	�'�������Նģ����r?S�YilqGhVt4�e�'�s 77�T-@�����C��^wT� ˆr��᳀��eee@cW-N36�E��xj����g(z��98���q���$���4ip�Ŕ�<��'Q�X�z���}H����e��3�6�*JrH���ˆ��.��&�Ť�'���y��jcy�	��������-&5��4�; �)}�h7�#r�>I߾�o4�i���V�;;��1g��>��B�/�;�F�Y���3(��UU��h���@Ǣbc�kk ���&)��i ��Iy+46�,rVLMM���ҽ��F��:�">������H_�;��R�V5�[��y�|����C���^�����f���)=K�	�`h(���~�,�n�3?�|��V�n�*��+���q�y�8a�dw�=�k*5n�.BT�2��zǲ�y-���?]����(+����G'S��욂 Vぺ0����l����nnBUǰ�L����s��܏A���EE�+J�xxWO���B�����6s?Ш<�fU����d��K��ǎP�߼�BĢ^��D�m�vj�ZUUՖ�v�m�m�F����
����<���R�o͏��87G��� ����߀Y�z
�߾�64\A��`cg��l\���֭�@?��ȁ35��,���tJdI��+X���:������/��j���]]3�E������y=󸽽��S�~�'�}3�5��I[���單.�'OPb�iRŤ��͛=ߣ�̱����>���K�deg@��g``�,9Tfe����5sß?���n8s���>���éCJ|�1��w��3M�J�*��ܖq��U.]�BBC��,���o��X��:�geA��/5�(#&��[�Mᅕ������c�7�5��ŵ�4-.,<��^�������j�L�qq.G��LLX ��:�4���Ra���@��2y��;�[=���Tn|_w�:�G�ln��"�Y	%00P�֖ ?*:Z5BZ��ʧO�>FD@�g@r�����id��[Κ���^�AhG��Pl��i�J�������	�_��NJZ�:�an�.t�4�rGg�v��i�; ���*��R��荟]Q�ƻ�^Y�}�5�B;���qF�-�QW���SP���P\�v���IĶ��QQQ�--�`R@"Xe��A����2���hA|󙤤�uM�~õLR����%6�ӧwmmR/_���
���u��	����LU�\kGǜ�ӏ
ɏD�N6�'��ٯ�I�6�{�YRsz=��=몄BqQ57w��� �pۣ{�VHѕ�6~� ���37�t����Wn�@�N�����&���}��U�:���ٳ��{�SŃ��E{ y���+������2����{A�����C7�1H�BH!���x�~�(�1�`�5�a �C��w��לh.Ug�����2ʷ[��o�^��PƯ-���+�t�, $��b���1��NB�i�0&M�� Z�]wz*�)SQ)�Z�!���!��VQ�墾Kg�KX8$�L�D�Ǩ�s�W���QY��lh
��j�N��	���x��
�&���N��7�Y7ղ�*ԝ���3k�D���}��JJstf�������&:1��bTA�5��fffu;���\��@����JIU�gO��f$x��Z}X|�q����������EL��˭6wwvB�̴^B�d����9��3倂QQQ��iH�*����b!�ŻQ-7֋}���1���f
�?�C�RRR"

��
:e�z@�����\����aq��fMH�������6z6|���4w�E	�� P(�t]'ss�6?!�Ia�_~�.�}Ν�E�������LUU-�eT���S�w<x��-R~�0�$_���r�A��ו�w���l��Ֆ����Q�j�K3U�y�2�;O������&qps�@�(f�d��Ykt/�'��'�{";������O<%"�P�nh�aR�&�\�"m�xp�E�#nnQ�ʇ�@�nܸ�4c�7;d���Rx��E%6opO�5���U�耂奬?\I��'&��� ��*����Ţ>��,@3��J4�voS�|���p��M���W�\D�i�/��=Y1�e�q��g|��gZZT>|����7�s��$?��Wh�_�Y�Ģ���!���b�����+�YqQ�lҗtI�Ĩ��%[���=���rrs3�W�^7�φ{�QR,o�7��=U|��m����.W����Ҷ�R�ni%HA�A����%�S�=�6߬2��[}MM�{��v[/����v�P�g��X� .�}}�ł�3���@i���H<L��ʯ���]Q��e�0��!�e&H1���4[�����HߖOP�M@��U��rƖ�����f�w~NDj}xav��k^^c�Wbұ��AC�,7�rj��LݥI*Z? � �erJJ=Ո�������bc�G�|�����$��!k�&'@)�x�kX�]�l��'a�|���"r@G-=K����?	���|@�P��SL��n`"�i�����ʩ�LB���EMLLD�7h��3�*Ɉ��#񻌡׻��wBi�K�o��%̉3�n�W�QL�Ŋ&&1�yŪ����"���^�92�ٛ40����m��XM���&'u���_N��}�};�ss=�G@2��`��d���#{r������p0d�a�q�VS�lZR�ˮ����uj\�uӗ����n����̳���o"��!��V��ں����nȸo|�_G(Y�Ggc�RF5� �m�<ruz����5�O5'_�����_��#�3���g�	��EJO��^4m��7��tx�0��%6��=� r�AF��`/�vmrt�L�'X��hZ^�������ׯ�'L��J�a��B{��ٰ��<���h+�?|���5�a��#l*�}�y����bddd��$�
3���3cq����S�xdb�"k&C��]+�I3�A�xY�9���J_�m�cwZs�y0?L��y3��*(�]�@�2����񕓚���]��Q\u���ritx�W���/�PPP�a1(*����?�G�OǏK��ދ?��b�o �uo��C����GtrI��	��rS:������'Т+iG�>>��,�NN���57�P`��l��0'����׷��DI9����
�L�zzC;M���&1�2�}���'*)ٰ|��GBB���\�#�k4b��T.Degg奓��[�͟��$HHIE�ݞH���<��I.���#��VS�T��!��Vf��3���)����\�CV\u!�ݕ8ew�T��_f�Q{��\�$��G.��,�Y�%��E��8�O�~Q757��4g�14���#�轜ݏn�aa�#:�f�s��/~�PcԬֆ���fb��[e@��`y[u�t�'���PP�;;W��@�-��J��f���T�J��-��=}\���M�A`I+��uN�Y�?�r��������2.G]�����Y���4hYJ����X`^��ލ�	-�:�Ց�:�W��f�Z��0�ŘZw _l+Z���������l�\H�j���ɐ�	��Ɏ%<4�O��X��n8k�����'����(w�h�)�eCb�<��1i�f�A�����ēݞ���X�k�4��,�rϞ���Q�����V@�.o��.�镞DRh����M=�\���ٹwp0]�b��(�u�][��^��Z4v�"% ���yC���«�"���菷��ee|���C�*���P��el
T� ���9أ�:��IS�����cR��$qx��|�o߾&��=��:���t]�?�:8�&��������j�ᚗ5>{�#��t����R|�y��%Ar�K|��9u_�:�C!Y���ҧ{�����,�V���R�,YG�_�U�4��1P������ɟ;&mz(O����������J�&^c�xNM�Z�����en��q}mhNpGQ��o�)��U���Z�߸Y���X{VJ
�ĳ�R�;2l둾�3r}k�B�s�m��@G'�B�	ӻ:�H1��B�k&$H�K,�+6�+ŵ�+��-�
?����}s��� ���P�@�9��8x||}x
���R�Wvy6]ݳ��	�I��?:Ip�n�vt�D�k��[�2.�!P&���3��7[}k�.Ql�#Тs� %)	Z�C�p~~��T1�Fv�"�J/���M��?��A�jdi���NA
�C
���7��٢Kx�<i)b 6x��'_�Y+=�����������=ݕ�	oRғa�Gv���[w�\������M���@Gyҗb�v�P�3��>�Ht�,�O�|6w�Ǘr��ꛦ&	B�^b
� �����	�f�L__����t[�aruiC�@�$̤Dw山��w��~Ml��2����l_��߸�\�A>~���qs3n�ۅ+"���\gb�������Z�8]��F�"��ȿ˴���H�P*���{����r �{*T
�ŷ�@��Av��C��s�WX��\��4�����V(�+��G� ��f�_�
l�&(��T�o��zom;;�-b�]�핏��w&z�
��xTY��M��BX�}}i�Ύ���{֖@��KC�ˁ��	�,����k�
�� ��g;x�ڂ)lllx��~�������Î�||;���>�\��P_ߟC"�c�[^��k�
����____Z]U�Vz�H�b���w �?������"0����yC+��MXH�+�̤��!&�`�:99t;��$TIFFF�%*�]0H��`}+�S��PR�*'������]1�W�������28���	.N���FH���?�B}ӿ�w*K�ov$��k�ϫP���h<�ng���	�:(�1܃>�������a���k*�����AC[T4��MYYY�^Aˇ��[�M�:
x�I��*����X�S��2�ז��� X�(`���?$��u8�b��c�nZ��Տ ����wm<d��qSx�o\]]yl��rӉ�Τe;R��.;��v�������!�P�솭�;o)�	�*6�p���k\y���Gl��B���n�=攩�M��)�
���	�BQ���Rx���Z�����`��d�A��g��Sy�V��.�6��$j<���qc��$CC�T�d�脄&p�ܝwO\N��ZHI�/�@	�	.����԰��Mj���9�0u$�s��X(I�u���yI(���/�e��
��ϽֺyMKCs=R��_�4�R��M�����˚��xnvv�o��Y�7��&@�y��UWA�"�a+
怆�DTj��g ����� ÐEυ���y��������踸��z6n�t5|�N$��Q��6��汹$WSv9��e���C�PGm}o��L��%���3E;�hC������E���t K��ɴ���d5tn�`��N[8�u����kѠ���Qۈ��iH������Vl��yz�DW���+0��*I_ڠe��rr�-��x�3�gؙ�N}S@[� �<x�F�gt4 $�-���� �K�|po�x@��ҜC��V��9�˩�g�����x%��,�bQMQ�rgk�O�c���M ���A��__���M	z����@���~����z�b�"�#=��
2�r3������x��=!^����]����x����B^s(��(�]��S��-���fFF�`e�*B�_����n�|?r!tC�_����<:;;�����c��Y/��8D��jgX�h�q1h�O����%�絹���d
.Ǡl|&V����_J�1�O�n!��/�yCԂ���3빧�!�����2h*�'��$�����22�rœ0St	S���]q��!?�y�'�r�xI��Xڃ��R9�ե;���������A�(��v]� �R���N.��5,���Ə��\y��=G��CNN/��m���m�,�?����,,��K����.�M�h�f��;0��.��.zE5��c��V�;��6k���rwT)��+t� i��D���9���C�J�V�^����r�ة�	vO���d]�m^ ߳'NiG�D �??w�;r�#t��򔊌�HB~24�@&G�SQPhl�s6��������v�� E�k���c~.�o+����ZA	��u9��X�2Q��H��QnR^�W0����ѭ�g䲍s�^�~r}�^N��`
QK����+B��4��w�o_&��V�}�
��2��6��e%c���ۛ���������f�����9d�w� =����|������?��l�:_�|��龘KǓ��0�u��r���TZ�X&2\�ӛ���РJHA������:� *�NC�<�q� ����[iiiVK=ԁ[:�cX�"<�ǜPu�L��:��ώN.�#0�ƀ�6���)Eu�0���}�D @
/ꃣ�&4�K(�[𘾏v�����sn�a�����4k�����~�#�tBw�g�[K�cG��7OI�i�o����-pL���\��E�^2�F(���Dϵ�'.�!w�Mڦ�$�S򠢸���NSǽ�
	��O��f�kxק��k<��C�� 9Mi�F(�Y�|z3�TF�vUm�&�V,9Aj�*�;bbe &�{Q��>�aX�#w�J�G����?�QX������>�.�RM��,�#�6:&����=�4ş��I�Y5���ZS�8{X������ܦP�����b��3ܙc�Ȧ��?�9��������Afᕢ=\�P �u��h�s�HM����^u���"���V��l��V3��	��N���¬��n]����_�5�%�R�Z�a���?�f5ю��6���=�q%EXr�o���t{`XII��9G$�F������iǅ�q:�9'vDZ/-�V�9�բ�Y7!..B�2����H�nW;����`�0�l�>����sna����fU��Oo�����]���ezV֐��i����>]�[�����>�y��a�S��'999���������֨�D,�@���'$$g[��gff��km�JSh5]ςJy���BCC�����@i�^s�8�&�j6�$��v�\�vN N������D�ܢw>��x�����\i�Sig�/���Jb��M�_��Q�|�5�U�6�s�<��o��, �ӤLMM�y��,:�
n��Y6�����!�jx�Y4O�W�vK��=��3|'����.9?�}q� �M
�c��kc(Q��N��N�?lͱY���H��d��H��W�#�]z'�X�wd	ܔC[Q{��5��tC�oA۠���y�
j%y�[ Iӥg�\�6A�>r��#Z@���a�s�q�=p�څhy}=�ӧOF���;o���edd��U�K� ����GN��?B�Q� �9�w6[Ӱ�ۋ�up�s$��\�.}�W��s�L#_eMwZ��+X�g��[c'���W�vJ���{��!�*��E����L��U&ݛ����Kc�q�Mh���f���\�=��aee%��!��e��#������;S����]Яx~`4DD�7������������a&��\8Q��2b��[NѤ��~���Ғ��� �lV=E�I����������g�����GKSFF�f�����j�0%ep������&�`Tk�����݄�?l��������G�A�j��Qe�Z�6S��u\H	���:�a^�#�g��=���f���Lak��艉	�nkЂB �����n�:/-�F���:�H����ٍO}C�!z��YQ@֑kCy�22����p[�ͭ��P
�L8b9����=�����:��dk�`k;ֲ)_}�+MrQ�#)i��w�9ׂ����/Η6���C;�"��n��y���<��D�(��;ÙZO4ދ�ٕ�N�Y�^��E�r������o�F<��h�]���M���d��ZeZ���Q�Ҳ���(R�N&!��i�� ��u���l��̢{mng����Z]�8�|||����6���/ZZ�����m�]@������GO,�P?�()!������x�w:g�-,�A�>Th�ȬY�Ӎ���fP���w������,� ^��`����s]�]}7-��?]y���.��8Nۣ���陘���J���t�ct���321�TT�/F;������F��o� N��u5I[VQ�v�9�?ڈn/���Zp�U�&Gӑ���f%��۷{cg��|7���.�9"��[S�6`l*��$@Oj���}��x�������T��<K��[�!��-/����돊�+�W�������B4ߙ�w`�#1�=���]]]*����J�UU���uy�����N��n��<�5S`8[48�6Z"و��$�?9I5??��r�=T��Sw�sJ��8�ܠDY�}c	��N���^ǹ ֔/�B�է�꯭�k��*�de=�2!��d����rS3�����k�7^���w��sr��C�8���3�%'w��'���ޅ���V1PB�����������f�l|[��̉ʟ-�
]�`�e?iŭ*O&��5i��d+��C1�hOO�o߾�È34�gGnrO6h����K�]�蔕�ޮ�ݲ��O�y�,�0�0ҍ
*@���̓��0�^s^�ֻq㆘�>��沎�[�[K������
l�������*ÿ��\�?,t��;;;���5B#�,Zw�OU����+���t%�!a��X٥go��8�� �b�d���*�N����V������3=I����W߾}���Ls|rb����Ǐ�u���¢�n{��j�~#��5�s��ۆruD;H�k����S|����!D�5D��Rb�/)�ޤ4k���n��XX,��h���.�m5�|�_�����Z������r�f*����)�[�Ԋ���mf�2��ϟQ�L_%�݋�Ͳb��8�='��)m���lh�}3Pda5�Seg���U��/_��"����2�|\d�~
J��JJ��~١���}f<s��USR��p�;��3�5���s�<��j��q�eT��%&�������߁۳O��U�ϴ�\ܒ�ŨU2{bi��xP�sz8�\�l�p#����,���X%OW<!���������\�T�z�F�ϥ�8[u�"����r��h����0� z,��A��!g�TJ�t�S/�V��B�H��I��7���X^���2S4y�U�#�It;���e�-,,r�f&e�l�ك� �����Ykkjr<ͩЭ;�q�f��4�w�Tn<�Bŏ��/�j�>III�d(�ٯ�D�;X$���t%
S������N���+�N�R�%�R�m*�EV��⧄�w�H�b8���TASQQ�����|��maP䒂��;4�3���b�W߫�55yA	w��B����i�<�&X	;oӛ��5���T��lsJ^�
��֝��=`�A&fc��5�a�2B���L��L��L���9�c�e6��(�� ���B�W�*x���AN���aTD���###Kqs�Ngg[-DZM+mm2�� ���%K9��X�g�����}���oo��`O ߾� bN�p?9/��"ۚ��id�*j�$���D��3IԹb�@Qť��E����3���;��j����ʟ1��8�T8n������� ��Ī��M��0nְ�n����I���Z�3�3�"��2�n�y���'�U��5N�&|"���k��ђr[Ff��mg�g��2cڰ��	,"����Ї��,��U�g��%@fr^�5��ϸbX6�|��]	�K���-!$@���3�g�ZL�7�j��4HyW�44�K�26�[�o��}�Du�JW�B����ӫvvy�yl�B�*��Ku-������$�5]�;ڞwJ�=^^^��YZ^��][��p�۩i��:ԏ�D�fc��@E�{�Q֞�,))��Y�w��u�W�E���s�aa}�4���Dj�� ]i�E|���m�f�.p��B~\pӒ����(`������oYYA��4�cA۾�\5�_pd�\$�2�ݯ��r)ss�* � ��5i{$+��Q��n���Xj������'���:X%�N�22L�QɟS֨Z��8r�?��pC�/��O���&���o«W��t�D���k�Q� �1H�ٸZB�c)�[��7�M<T�aI	�߃
�f󁁭u,��Ț��V�lgg� E�b`�����u�0��)�<��'W��aB�Hg,��=;;����A��S��z��y�?�&|Hw�:�Z�8j�gc���P�'L���x\�N0���2�J��ap(a�o�l��MfFX�
9+(w@��/X����r|Oulh<ާq;��b��@�7Fk���2$�i�:��+`vTʬ�3�j�:�Ú�����[ff�.4�Dʂ�%��@�)�yp�r�����&�r�����0y�/{�sHV�WJ<y�$�.�D�����Ø�E}nmo��t@�y��A���ZDQq(w���$K,:˨͜`x/v��j�

�5��HM�+3s� ����xX�ME��,|���B�#���+[=zgmjJ;N�����7�쾵�)ȸ��偸�i��A 
9��_��)!�Am'�!σ�����ք������9�Vw�b�3;�W/%�[�a#�À������8�L��G^r�9��������jjtA��k+��k~��ۜ�_�7z^����8�:�;7J�:�_�A=`JIJ��u�����z�<	(:���F\�r����F#+p�8�q)�8�3	���.�;3G��/��AC(�:��T�.����i�o��h��n�1���z�W����A�]8<po�ꄩ���.~�XZBڋ�[7%u�XJ��b����!��jf�w���ɸ*yCNcA-|�1N�Li�O�kȏ�p�ZwH.�Fߖ���6b\ �t�\b���`�^�����P�L��I L�KL�F�r��^V�^ D�u������)����M��N�����C���L߻����ť)��CU��j7ɐD�;�3J6*tĹ���M��������u,��X\r��{���h�ZU��˝�.��9DF�H��x�<)iH]�ԁ�禍�D�[r�S�'c����b����C$/��e�����,v5�9W��Ny�Sz5�Gbk��9�y�OQ����3T�8���hs8d5g4&�)4����|�	ɏ�%2�nTt?6�h������չ���ʈ����x�����9_�Y6X���b�@���qL��=C2zXdP)��]���yv��o�x�o�7���Fx#��o�7���ƿ7�^�_�~B?R�ӓD^a�����a�	&�`�	&�`�	&����>j���WjL0�L��t���a��[R~����~b����0�L0�L0�L0�L0��oK>CEz(�G�'�����Q�ފ��נ�L0���hes�c-��R�`�	&�`�	&�`�	�?�3mF��}�������rs�n��L0�L0�L0�L0�ӿ1�j�B@<g)Dш�����p���ݻ']��� �o�&�`�	&�`�	&�`�	&�`�	&������R2�+�
L0�L0�L0��I
���X��.�`�	&��W��~AY��^&L0�L0�L0�L0�L0�{���R�wW�(���L0�L���xw����WjL0�L0�L0���1��/(c���{W�`�	&�`�	&�`�	&�`�	&�`����k#yЏ�w�W����ި��
��8��L��Z��v�L0�L0�L0�L0��/O��Kɰ����+L0�L0�L0�L�=��$D�?���&�`��ߙ�)� ��]��<����*7�P��&�`�	&�`�	&�`�	&�`�	&���z)Y�)��w�	&�`�	&������A��\�/�.�`�	&�`�	&�`�����e�W��&�`�	&�`�	&�`�	&�`�	&��=�|)YޝR������_P�>��\�/�.�`�	&�`�	&�`�	&�`�	&���z)���:��w�	&�`�	&�`�	&�`��ߔLʮ.��Z��v�L0��ѝ�{Z���Ç�x��^�e�^�Heܪ`d#&���0p�����i!�NCxO�^H�����>	&�?�Z���痡����ol�yW��W�������������������:�p�R�r��m�C�Csss���`L1��Cs�92p�G�F��g�·C�����\�"z��;76G��I��:8<���o�DGU�^�5T��L#U�	d�L;�!SLc�Q�[��#z��^�<���W���泅���c�Jt�!i�UiW�Mu�T�װ�(Ssu����n:��G�=�"�K�bˡ�ܷ��0{voc�m�k[cpe�zk�N]�ET����躹��iZ�F���VtE���՛���H}�����	Q�ȕ!u}���wln�.L�T�����:�Y&��f�\�A�mw�@����v���)��S26����'{���DI6������$��.$g�ܓk"d!ȉM�(=��⒱��pر�����+R�4��/_����7	�|��c��p���J�w?G��� �C�x�k�V��,e�K���`�����F�cZ���[�o�<L<f³���]�ŗhB�;fQA;˅���%9V�@N�eR�#Q�n��y��;S�r���{�u?t�u���H[\�I�׋T�eRH]�����}D�%��*���g`W�H�xe��\S�[��T��\��֌��l��6�=�Y�7��J5z�bi��a��{d�'<(���>σ��e������ǻ���J�E����3Ol��^[��(E,Y���ʙ��؈�L��
~�(�Ր�d�#
"O�J�T�p�YXZXq����9;��ɸ��F�u-�� �2��=�����D��3QQR�1?�B*)�D[�n6�mQ�^�s�����dC�x����jܾb�~�0�T�ˢCè{8��3������:������l@�����I���~?�j�7�p�{Jt��@gg�JX�Mi^۾���p����?�����9�芔�B��8/�Kx0\'�ݏ�mƨV��w�lV��aw,���w�UT�#��dŕ4����0ܱ�>�2?.�z�t�2;��^WSW���:{�h���J�^qT��0�Gٕ��ObZ����p���!��H:�m;�0=.(��eu�t�`H2��n~��}RV�-��X����]�Z������y?%�M����#���5�B�?%��x:��M��r�����5Q�� S�k7-؁����H���w#ׯ�&e	].�i��*��GM�r�m
qZ���o��I��>�D�߯��ש�S}���}%�._�k��\�Bف@8��q2���/&Y�⨳����M{����
s*%m�]<�E��h�z�z>��x����8�T����h����(.�ѭ+�/κ������fpHm+�msj��y-�I
�_��B�K%�d���a�;��d[���?������^��8��(��H��u֫�5�|��텕~��h�v56FZ�?X�V��ȃ~P&�	�&���|5�X��/>ݽ)�`gWd�yl�[h@���\������Yyb��h�p�aƑ?h377��r�>H9�K��@�A�"F������J��E*D[����6D�9w+��H#g~m�8�<��@6��;88����u!�bu�e��m:�D�*��R�֗�1:ܟ�_��~"�aC���$��ё�����N���0T�t��2y0����38f�)���l��#|>�ko�̗���|{Y�a*��s�l�b�e`@���'Q�Bg��A����S�F�҇wf	F�G�*!"XB.���-��_��徶[�/0��9P�#R#Q��$��-��ow:�۳��9 ��dҡ��Ч�ө�̥7�@�1p�S-!R=�������n�����L?�����zQW�*���HV�����hBv��7�$�u�D��kιv�k�NJ�'����X����ל�]�֊e �ܛ�:��Nϝ*�צ������O���hbwQh>�G}N1�m�����F�;�����5���d�z�]�[�QiQCmL�����V���q~��W�{v�2�e����-"�C��2���k~8���_���a4�(���ф��ؑ;/����st->z���<���k�fW�2������kpegg�w�4�HQ
��n�&���8�ܽ�A辬��N����&/ϴ��N=_c!��m�՟���/���x�&���<���i%Y�nn�s<��w�拇mGG�`�bC������X�޻���Y���G�ÑH�v���L�jv�d�f_�y�b�����'❶���Ú�x��Pݰ{�XR��B^���Z���č.���z����M/8=���tp�D��w�V��	�I�A:X����a�'�`��G~���"m��|?	�0˧�mf�^{�k�Η��$�L�xS��,0����^'Am���o]�M\��������g�C큛O?Tq�QJߺVD̥S��/`.�LU>SUSk�i�2��6�{=a��!�=�%����V�����{OP��y�_�����f��37��(�ڎ^>}���K�V���=�,���篤�������j*�@�RT@�4��;( @:!t���{U��K'�I��"��N@z�.��|�}���p���F`@r���k�5ל;gĕ�6�}៯�)�FA=M�|AM�9����(�77��rL��k?�������BB��t�����)���3NJ��^�7��&n}������\ɽS����d_45G�E�I�pss�]�ٹ��i�'����G�x�G�<�W��_�j]�|)�-fzx�K�8�
�{3�}hP��fl����!�/�sI����O5ǌ��=caA��?W����n�^%���f�"�����*��Bic�$����m�1��w��J���J���h�QǦ�y���w/@\�]/�Ŕ+{�v���D������=��X�s�S{����/	~��m����HJ�0���O�)G�·'S��'ml�'���!�g??�p�p�s��h��0�E@��&ja�m^��J*%����k|�� G5A
�����׹���mm{iISa}��{뒜�܅ВZ����W�e�2�Nl���$b�����;�D���J�6m(
G���V��_��kk�Q9V����㦴�����1ы�������Q�Sy���1�٧?hqKQ߄����I�;�1M�H��P�U���c=19���R� �%A=��}���l�Jː�>HK��[u�sɑ�~LR@O�}�g���ya���qީq>���� �C�OWP*�ْT��
�.�K��9�Mz:A���J� �nO��^d~����c��ӧ�A(���o������n�a�枈&��{g%�r�Z�N	۝�2�����Mӏ6�l�"C_����}�	��:q�[�.���C�G�����/����#������VϷ��2'�d��3%Eg�u��R!��Lԑ�$��͟�'�B��MG���1�� /E��_f�4�x
��4�D=L��Ώ,;8 d�[��Lv�*~��J��yyY�"��v�_3؟/al`�����%()���<*���"J�)y,ݒ}Tk��j��ZX"���u]
$���
M�I�<N�w�c�P��u����'��ʉwMEE�i�n�Fߐ�^������j)��["KP�_������GIќiE]-��b`���k���X�,Goai���򧈀@>�L���12�*�WH�T����Xj��@pۚ����gw��,�ȶ_I�34tvh��w���-z/W�FGG'�<��߇W� ��ﴜ^ijj���O$=c@�ȗ��ir	JI��eNn'v]g{x��}r1�z����|��ϯ:��W��g�SO��΍��_o,T�W�-�j�¸ZY���]���ɩP"�� ��6j��в޸���,f������V~���RRR
�bc1������;Y)�S�PH�[[��}�?"��%z�,�@)M�yv26��'��-0R�Eڣ�Ag�s�i��l_v��7)�P�Hʿ�
8��Y��O�}{T�.�5��}o��鋌� �{O�*s��?�W?X>������]�����z[�!�w�>sh.f���3,��q�=��邟)��^��iE����1ޜ�2A�Oe}�**�$�&�^t�aqDt�����^��-�cخ�޾�U��"�oM�~�zz~�#R���$	������!0=��DP�
UUUU�J��Ard���p��e�Ǟ�Յ����<�)A/MO���SQj%��N�G[�y�.�;zh�II��������+�gҔi�Z�Ҥ���<(Z�w���x��iUwww�e��0A��H�vm�������AK���i�3�D�X�޿��#��v���%g�w>J����DH(�"��@�&r(A��Υ�7h��K'�N}߾b��ڒ��H��� u�
�-��"��X����Z^��'u�����{޾�§ÊqW�s.]��\-9992(I��8$�����'xv�������Ǌ�H"d�n�9�����&_��9ބ�����Fr�b+eD�;�ܽ����6��*�q��q�Bq��'R#��*��y�o�\f���P�w_g��bL�!i�to{�)�ĳ�������њh��Cvno�u難?G�HW����2�V�cl,��4!��	�Ǐ5{b#\S��4Jpp�$�o�A�r�'W�R7�D`Y(廮������~L��VPT�Z�K˅  L����
�"������ɉ��<T���mɂu�֦�f�d�+3�1T�W��:qO��f��O�L1�esW�����e����BB�[�_���b��PT��/Sc�=��)��桫��f�~�%"b�`�����R�_Q�ȆZ�d�I[��ޞ��E.���h��u9:̷�Н�W9H���~��/!T���jJz:�����III+G� �*o�)_Kk��H���x'��;��猋>[~/�ˠ�����V��ֻ}�I�R���(=�~�n:
d��Q{�OΌb�i0��"���QV�znn�A����&(m�.F���c	3k룙��V?��io+���D�xb�`N��Td:�}�;#�%�c~{��OWޚ.o��9pN�a�6ri��x&*�Sܾŵ�C"�m������ed��Oc?���������Y,D�&���oף�8������9��.=�F[*����i&�ZU|2_<�!1�������2�x++m�6�f����]�/94��G���|�3�-�"�����r�� u2�ގ�N��������$�͟����:��p3o����ߏ�$p��wt�֓��t���%bҎ��ےP�����*(�C���*�b����8!)T@�ER����gIK���rkS)H�����������������+W�bּZ3G��z+1R���L�G�ͩ�Ϫ/]]�3�ܙ�����^�Wti),N��#F�b�X�̗���~7T�ADDDu� �gl,��?A.�;4\��;��C���������� �_�?�:C_Sϰ�#��2���| C��ڥ�����'��f �{,�BN~Ql�L��q�'�r�K�1zsz����%>ޘ�?���#x�
UdT�ې�j��I+:p+���:4Y�<�dw���(�?D�����o��ʈ��2fa�}
	�Lj�~��-�&[��?�Y�uJ���H�`{w��/�գM^��A�S��7��TLO�>=$�J�prRgg�|���ēxS�<(�`��9��c?�rH�͛��	�נWX�ĄE~\�2��}��]�=��~�|��2�r{�A$��5�JT��+�劃����r���((Vy�^Cq����u�S�Q���m�y���x����=h�	��>t�����[yI�y�/ehE�0���|�%�{��m�3��&�$�����?�J�Θ#ۖx}F/�Q7�e��ߧ�A�e�~��쭬�
���k�η��?�xL���vcs��EPg��ܗFT��¢㋁ ��A�At����PӺ�g��GOAs��Տ3�\ќ���I�5��95_wí$�`�0p�]�WE5����Z��ǯ�ə[=���㋿�Uy�����bR>T�z���۷oR�ºxq7�h�/Nw�@�(,(7���T����>?���	|MP�W���`&�g���o�����K�r�0���]y<c,Ż���^J����`�Tޏ0�>�8�C���mt]����F2��sM�[?�zBDB�%q;ȭ����(�����Q1|�ř�)#*�-s,ՠ���"���VJ�܁�~���ѝ��E��oO=�Y<��+*�#&���ƴ�N�yW��˦�{ �O"x�� ��3j�O)	���X�=�8�7�q��V�`���첀]tKi(2ƞl�Z'�x)�aަđ��s�Eu1I�J7�j�;<����:Z0��,��}%u����i�H�x�3�h.��z\@h�2Uq���r�C���Vzʰ��~�D!�znAAA�M2R�"ά���]E�V��$bY�6���ⲞVs�fIQ�=��?@b(���W`��L �+�����K,������[��v�J�������_��l������N��a(�}���R�4N��}-�݊�T\:v��녬1+a_���nF�q��z����  ��_����(a�/��.k_d����h�k/��QW@2�"ӟm7cr[�˫��Ʀ��r.F���������\!��j�V6/�"�X���Pv��D��,ȳxk{����J�D�&X��/|y��|2�Ȗv���05��o��}�<���󷶶8"8�~/;�7��N�|�^⾽�����:c=�ަ�ʄ䯸��OL���qDr]�������l�0����2�� �PI��K!z7�W2�h�N�j*ԞJ��k?~�h��%e����.T[�P<E�g׽���PN.X?���K�4��ԍ����hO@�6ƺ1���A���e�Q��\D���(����-���{1�N���s\���1��x�"+~$��y�5��Qc�B���pku��[D�����Z{'>�_~-}��ׯ�o��30�ӭX�}b�rM+P�fp�����M'���C���F���Ǟ��Jp���Wn�I5ڥ��\��D� �Nlm�j���\WP�v[�' �f�7L�b�ș�	wՁ�	#U�<9�C[5��S55u%O���l�W����F��l^�������rH�%511���	��5�ڣZ�)�:�y_fxh��f�D����&7���EW�,#0�������������7���ób��1����sJ����4�4�#��X��a�����o��QR96��kXgeM�N�H�J�x�)��xeϹ����o�qa�-� ���@�w.���������dѝ��U��s]�5}Q5ͬ�5�]�!��f�W�M�������Hy��t~������u������q3O�����fj�,F�e5����-���
��Sab"�>����q|����S�i�+;%ϸ�5+� �����l��?<�x�q�;ہf>��p3��mGp�q���6���R�#�����T��@MebT�<������{|�+k)fdם ����x�'6z�%u6��j��` �J%K�\W�k���F �&�k���9��E\?�=ʞ!�=ư��|g�X���^��|�i`T����%g�miɬ`7*�,F5]���ǘ����0�z/  �OShmm�e.��*��y�)5&%��;+��PM!ѿum Cɇ"�����{�6�c�������v҅�\|d|`
k;;�"	u��C��u	
L#�xXޗ���zu.� 6���I91��)qޞ��(#�`�[���l�9�,��"�5d����3oO���-NuqqyI����ʪK��pau�a�ꮧ��A�t�+�Rp�ոs�Kc���i�Vg?��B�&@6������X���`�HM�;?�k���k[b��;iƋ�9�3'�o�7Dr�S:rǫ��/c��~}����P����)0��/,\��j�|Y���j]�#*,^1#=c�8�"��aK,w� ���1����c >F���<�~hn� 9N��P`bJ�}��(�tf��&��1��ƭ��O�9�
�=�����ӁB��ճ�e0|[����C�v�$��vy(9�L�
G����\A�����b^�>t6��c%�&5f�9�;5y|rNNN"2~�-�\�!�\oqc�ݬ���:Cj;VŽ�O���Ĕ����0�C'>d�勼��É����!h���7�B�����X�g��|��r|f&u��5-�@K����퉘���x�u�jd�M��muI�Zl)����L�ߩ�)4��"_��ͷaz�~������p�&\���W3��������%%mK�ޕpO��@�������>W.�x�hm0Csl���]�u�?�o����{/_�lX��hx�����ˢ:��u����ُD9�o^�&��l6O�ˋ�-���%ip�C�3���ߔ2�+~��V65� ���8+���������)f���PE�� �;2���wgg?��+F*�^��gQKK����R�]C2��8� O��4ɥ���H
�s
���]�J�?[H[6hJM�v��_��(��/N|r�P��	�du����(�V�~͟��p(��Û(+��z��\��I�N�[Cl�[`7�� _�{�,�t&Ԅx�'�n~�6�Y) ��w1(��^�׳��[�f�X���E#�CW)|��eD��^�(MTDQ��U��Ѝ�E�˅���r,i���������rO��APP0b_������/��ɩe'7�7����wz��6彐6��i�b�����ꗺ�u��A�}~L�(�lC[F,u��Ս�ί���P�I�H�(�y�B��oG�s.����sM!~X���1h
�_1�<�aI�"�]���E�٘�����Qu�
��.G��F�ΰ;
���C�@5�J�x"& �X��O�8����!Z��L1��ff4�+>;Y��)�%W�4�c��/-��'CC����m���2�� `�/��U�Wn��8"�H�C?6<�t<����|vy}xy��d����r@�,P��Dh��3<̅\�0y���f������X]�|���H��Z?�"���lݪ�h�R�6/U4�$�'�1����i_X�f���	��E�׋pcu�ľ�����b�Y��:ށ� �(��~݉\���\�;��fll,�a��Suee����1i봬ɴ�kEf6�K�G�+}%�x��X��eeh%k�	{`�k�qc C�nH[���$��Dc������-q��z�T1�p!��գ�C����]�m"�^���`��L��"��}/��58׬jZ��8�Q��|�7?:2w�T^V�mq����!�XCu�t� Շ9?ɬ9�������-�B�>_-@ƃ*`I���Ӭ~~3���
MLLD��
�{*��k��s}6. ��s(?�;o"-�����L#h&�dt�/���ȇʾ���CjF�@K(��xUW��V�x+��OZ4G��\:B����Th(?�5u(2�������C����0<L�!�/N$<�&���U�q)2!���t��lq��,_BZ�oOQ��E�E��b����*�HL:� S�������A�4����Y�����4�q ungo䢚�9�xސ� ��̅Ȍ,8�*?E���F(�Λ��	�єNX���W����2���&GFF*Z}��3[�L�7�&�ߌ�����ٛ�'|���� 8��e��ȡ����B�2�����3T!5�7 �6��{{�'��W�˱��b��� ]@�r��|�_�lK]�b��eh��+*[O�� ��ۋD"5���M�������Mu"�Pqs�8��X*�1L�
ɯ��-p.����k�`c�T�j�+�ū6z��Ewc��2�_����l��w��"��I�w{}��^j�~��$�DR�vq�A4a��jv���|��d��L������#�I��9GFD����ro���3A���y�(^֒��kf�f��>~��=3�Q���Gw�ݛK]�[o�=��C��?n��J�o��~��Oo�a������V\?5���o���MU�A��q�-O��9[��*}S�05�U�������� �K��0*h�9g��1����p5��3�+�CuT�g�7Y:E����0gьC�fdq��{i��}Њ�ɽ�|~2m����L�¿ �Olk��� e��K�?V���6l����n�8�hp1��ũ~����Js�p�oB���C�Xe���X���F���钳SOMO?��Q��j��<(p�ݰ����`#�J��`������A�X��x�@���Ƈ�w��v�xݎ���޲M��<BO��{Z^�� �\��p$ZQܠ󆅅�&+�Fw
����3���`]����m(���2R�8૮u|?M��͎��q�4HR`��"{ii)�����|�G���I�Ώ�-��71�8��JV_SS��e? @��*\ �q���I�$V`Qu'��|2$��)��%\ƚ�б�yx�J3���!�]�o��c�{� � �%�DA�E.n��&��O���������9s����e?���	`{��$"��ܵ��A+�'�0��Q`x?}��/ �x04b��+.?Y�"e��a�ga	����kr��JY�f07`歭-gIVV��j���T따�����Ե��F�r"�|���,�ٽ}�T+|��>PSR��)wHG�hA��NS2����S��KJ�n�g�U!#˖׻
�x�Tq(ݻw�&#��A���S��6� $�i��>�qcY�7�;8Xz���|�2��� �P�$��i�]�o�Xı*#+��z�{��6�����ֶ����]�ّ��C	����v�ټ�>=�/�O{��uyՄ���ڎ7NSy���߹,"�!�jWDNN����|�@�,)N�U3	]��X�	iǠl�:'''+]tqKˍ�����w_�e���Q~�Y7'�d0�Ήa����q���-h������O"4]/�7��l�����AGҺg�������I����¼�=���[����Y�2�,			k8\$'v7�syxl,A\���*�xh`�H5������p��\�b�
���A�����Ʀ����"))T`����y=�jR���nt󋁯,�6oz��OQj�im�##�~z���"�W����Y(��$��-��B������s��51��VP����L���F	����(d^���<`-Z=o�k���k-��_\I�jn?cv�o�����㣭���1w8=l����6X1���N��+yR�L��Y�U0���0e`C~e�X���FW}��z|g��ѣG���$!'���j����¢���W!6I99�n����By@[��@y��k�����������h�W�Y����]���9�LS���������e�attt�Y�������6�G�t�]���Z.�����:�붏7GEݶ�������;9�0-�W5�J]�1���,�ߑ�����Q֡��"�b{{;�O(:���)^��ia�z���N8&̢
����f����+��ZZZ
k��J����>=�X�/�X�@X���^lC���I�M�2�����:P�<S��^���5�,ѕ��0�꼍��]}�8_��g�!�ƶM���WKK������uz_iF:Ǐ��ȴ��ȇ�� H$9�A￺�MD 	�m��<%�ͩ�#�vj4Z�W"M���7��fqrz�|������������C�J�\����q!~_�\l��Ӓ�+ԭ�0-��㣣�%�/?�����2ǮXz��E�%}������������/Q���~ͳ�U��\PG@�����k�� �g�$�����#'��e�>���bTT�^֡�/���,���ff����%�o�:��LC�{�R��-�n`�M�N��n�n��[�233�,�U�+:p_�&�3_��&�j�ٹ��2P���c���O���[A���(Qy�"8,	�*; 3j�֦�2�՛��#	m�c.��q��kM,.��u�,-U���E�>�a����������\�RD�4��7�?�P/*�{L�[�`�(����u���E��.+`��9�����s�O6.��V|�<߲A��iw&l��9��{ɭCS��:�	�g��ߤ���4���~Fmcn.�س%�8	�I�g��kBL0a��%ۭץ4�ov�� �NO�k���J�nc32J\�=82.ʼ�C/��{Wؙo}p{-�u��q+����_�T���y����'���Ffo���]�����c#q����z��?`�/*T����,�f�^��b]�2��B�1l񗁖[�����W�����[J�VX�2�*a�Hcn��5X� K��zh����*[s{O)i;UZJ��O��=*:��~��	AE�?&t�pA�5U�L�^Ħ�F�OW~gn�pr$��SU��oo_~6���l�{}��L�%y`��G`��T��Һ�����A
�[���"##���E�
:+E-��b̠��탍qU����MlZ��늰0��9���A��՗���S��Ƨ��::^'�a:���qbr���zw[��|&���I��5![�@�/�F����񱝭#4mL��KD+�i' U	�i�5;��~-rX��<1(���0���:i����i�>���9�,ɜ�>�x���Y&�~�|���i�S�%,+���m8r���(x&�o��v+���5ətc&}㝌�f8��0���D�#�T�H��**R;�NR9���V|&J��|?���+]۟%����K3���tbr2:�***hA�Wz̄�_WS�����J�����'B���V�r}R����L�U[�+��\�{�2bzxǫ��K��-+��ݭm6����-�詟MStUZ��,EJ\F����b�׽�9#vUMP~F?��d��fK���b�pZ���Sq��$�_i *�Я%/Ot
���\��ܒ��g}64��OF[A1�)0�~�������i�=$�3_�J
�+��_�Dn-e���вS�%僮�w����J]���ףǆ-^��8X"����.*FM߷{u�G9eeo �Cz�Cڑ0��w~|�����k����}Q�8`�Fss�7���P8f�&���:�ۦ8ݺi[P�چ��Om�6��C�X��P�ɓ��ڸQ�6��#��ݬ���7n.l��ܔ�䂷��GOe�p�:��Oe~���{@���K~n��g����\�b�����J��B��jBOJ%�&f�<8\��z*}���>�}����G��~���YԘd��r�k✜k��6�Ǜ~�NN�����~N�~�$s	q���s��,T�C�	N����='n�ſL;���D��r���+G �<-�a����?*��k�=�}$-'��#��E>������V�Y���G����lnC����J���ܵ�4�����=���������%��4�;C��&D����_Ƽ=TF�p|�e� q�岹��r�Y�g�r��|��_R7�0GUS|G~�4�A�\1�kīqm����j��^C���A�����>���G��(���İ8�+"��.'so����������j\�UUW��,=h$Cg>��f��Ը����X�r���x��v|���|$�2�qZ%qqXbXR�%���k� �m$�'n�F����}�n����n�>m��QQ���M�[�﹣�"��Kj���l�2Cͳ��Z�Q����*,���r�7��>�?ꛠy�+1�/ F��C����^�aeG�Ѽf��r�ZB���Q�m��i�;f0�ظ��\�+���Lq�OykAp�$<K�@	�1�NU:�qgW<��Zߟnwh�%ŉi���H� '����>4��i�X*�
~������}�/�,G��$�VZ�e1:7]�p9c��V���o�ϩ����m�]�:QR/+ܛG�d�=��Wjnn8���gf�����Ȃ�ֱ��oʜ۪Y|���%>��j��� F�le��)��z11���x��l�!���5��_+���PZn$�|�0	l-M��zlw��b/w��L��xN���~��� ��[��R�H<c/9��X�!���"��??s��g��	a�pj�K�C|�,5u�2�0k�V�ӄ�cGU�9Ut���j��m�� ����;����Q.��ц�7V��W�r7�\� �D�P�8ifTUM�J8�Ԡ�hu3'�|�]dо����34�w���kɖ��\o��b0���]m���p���C˓z
�G�������f<�^"	�]��$���k|��k���A��_g�H�ޗ��b�d�Pd���6̿8rr�M�0�U%�ڐ#���`\���ܢ�]�qVX������*�6y��	I5�����5P�E���<A�q\���R��*���,ۺaB0���q;�}wm� 2#JY���NS?��+���k4 }r�s�*����h�8��Tw�)�Yz�%h�3(i绦nW���Mc+j,o!/�CƤ�K �R��<9������'s�k���1M��DG"L�h]\�QX�_����3G�Z�[�s��=���F'$�� +�:U��EG��m��`���+^����v�KH���|�����  ߔS˰N!�t�1�������u����v�_��xii�w_EM
.3N���U�b� �	>�wl�	99���yz�o��Lz�iT��EM�@�t&�}��a8��Uj��Y#��%
I�\��E�ٿ���,3�;��(0���}t��Eoks�ypi�) �T����⽃�F"�Y�Byaa�c���F�n�>�}r��ip�+k����J%s.�Qɮ��]_8 �<���z��v�$/��7�u��
%ٵ��ʌ��ן!���9����
��TqGcYT=�m�i�k��?d�X�>49��f�����݉qڙ��|k������2����0zn%n�VK�4���i���2B�qI��M�ID�0+M�&�T�X�������X��jv������܅����^�����:���y�����AgU�߇��W4!0<�e��V��K�5Wll��Aϭ��"Vu2:�Χfp �)����yjZ�B��c����T2$b�茕$XkݽxaW��("*& �Qm�u7���[��;>��X3׷��.Tg���,_yzN7���uV��C��H��[��t�I��R!�����ީ?�������>��O��pq�g�#�NSYX�	o,Ui��Q��y7�B�$j�_4lr�~c���9{�~��]�%�+�6����*$�:9�<�Z��3O���ڳ��E�>a�v�����;�xtMV��D�-��$A3u��u�'\�3kc�B�������9s�tTݺ/�f̗���4�X]����le�P
$��ou�;�z����U�W�w?�(�RG"��[��П�QONl�}�򪧙��jzz( `_fx*�I�<y�ԗ����e���b1�q���lj����t�R��Cf��)����aLl>�qV��A�[s�Ĝ�;z@r?��KJf��)��#��%�h?����X	j���b��U�+��W-ς��ɸ9�猐�0��U6�Yt�Yt�֣�"&:�����g�&�@��Y�4sWHl� �A`���d2WL��,Ϫ%v�F0&&��$#!��i�ɕ�==�q
EL^�"u��ۆP��0�-	�t@�u.b3���n�<lv��P��PO�
�ҡ�cyI�\��peeD����|:ҫ� �ˬ����j^�,���4�h�cc�km1zI�R"/e�εxq'p���{�]k< DL��ȱ$�fcw���b��
����o�4�����K!g���ʫ?c�%���DM �J�5c��@�vI�sA�*�?C�O/��v�-��cd@��񿎮;>�/q���?�0��/��CJ�?�[��
������"A��9�7�7���C�ߐ�7���C�ܺ���0�i=�w'��� ���������;�G��?E�7�e�L��?PK   ���XT��"  T$  /   images/53cc934f-9b11-4097-8823-694d19808ece.png�V�W���;i�鎥YBD��n�k��NA���f���e�%�}��W�/oΙs��=sg�|�Q�@U\j\��jJ���

�(6�U����������u�N���7���]�yz[�[�x{{��9;xXZ�Z��dB��QP���+)��d�g�|��=|�͋�PT�f9+`4�P�ЋQ�[(o�>_�T�1��tj:촶�[���)���t�������O�Y���������r*����ן��j��Z��v����	����}a�JJ�,�����|~݉�ػ��qek��#��M$찮�����!�=����:���L���f\I-��i�=(����g��[I���Q'F~��6��;�c66R�M��~G<�2��}F�D%��~���ڴ6h��;�"~�f3�K�M�	����n�i�{�Ź��1�3G�A�m�b�S���L��F@̩`m���ԓhsxC�[�*���ja�b��+�" m"0��Q�M��O�x��_�f�㣹��nU�0���<���@��D���;�l�����3B�JK�P:�\=�>�{���R}<�^\�a�iiݶD�<䲡����WRl�Fյ�t�ɕ���*�7�R�b�<c�iN��L?�L�|=,u�|X���K<���5/�*�}k�S�)rߗv6�펽�E�P�kJ�v�_���h�e0o��%�H�"�ŭ��,�v���˶�z������kB��&{�+.8|6)u.^��~�rv��8p��y.(��7�z�\(�S�-z��?��T-�0Q&N<�/ٙ���i7-q�!�����{���I�Ot�2-�MLKYՈ�Ln�SI��m�ڱODsO\��3eZ$9xzeU��)㚗�,��M�pN�.$:[Z|='���3���)�����fb�ѩ���Ԣ5Wd��1�4P5�b"��Bg�!��D��A��$��'�fS�Wn?���[�+�=�����<��&?���\,���-�%&h`�W���#��9����ڄFd��>�)�ק��ݽ2��+{�a�����w����ӺS2����h��-w�̾zG� �d+���#c=�G�~�Wؾe�P�+n�����f��G=���Q��F�V�0�n>���DP#�Q.����ųN�^5i������Qc��-kA��"�����4J	Ĳ�[���k
d�I'��%W�k�k����@��b�)��H/L��rxg�CFd�S�����uEt�HEx�3D1�pU{��z]*+ޏ�Ցe����*�u%�9��	!_2)����RhY�n?��q��	46��W�Zv��T�+����i	�)5�pc�C��\ѐ8mZ#� r7{�M7������K�7繥8�I�c��n� ��:z�(f��6,tDODw����r���{��%���m����W1\��-�4k��*�"�قg�6��hp���Z0A4c�]�
E�ʩ>�8l�y�nT��S.?	���8חT_z}7
�Zs9������F�|&��焺�~�	��x�\�;���KI;Qj���Z��x�coSTM����m���H��mʂ�U֊�wn�l��]���^�"�Q��p�L��i1�*�{EX�pr�df΋u���erG�Z�k� ���A�ջ���}�pf��`���������=�h��_����	C�W<�ķ\1Nz�K�'3��U~T�0��%������u�ڀ��Oo������*���V�6O��ɂ��k3J�8�'��W	�5O�}'��^������g�$�����}���C���v�8�S	��?6����;"��C�Vn�Ba�����H��1҄�-j��%ö1���2m�D�9zˡ3�"Z1'9���-	
���v/g�J�q��`QK}hִ=�{� ��fTM���*_�0?b)�Ω�wMkO@&�ut�mf*t���늾0��d���|r6>m�AI�s6��'�-��8�����+Y��������0��a1��"�(-�͋��5����S����9 fOb5��� @����w>O?��`�~�2�0S�ؒ��1��`(L�'��K���t��?�*�K�,�ᕪDbF>�Z�F��`�y�;�A��y�tj�XXja�\l�)�b�=/�P�J��2V��56�Vk?����} �Շ�G�X��T���\��W̯k�;����ԌL^�0��ŏʥ��r��/0�Ai��@^�0���{�WM���[U\���h� s��'n<ͻ)�\Ǒ��t�b��i�H���Zf�"�9I�Q"O.�,ɗ�6���f��t�ĩUm	j߱i^���~��ïs;��������u�)�ф�]]�m��͓�4�/Ikf#�b����b��F�wk,U��D|}��>���ĔIX4�w�4���ENQ>��ShJ�MGGڸ���.��|kI� 8��0�r����qH%h�A�h)��[���)�9����F��@Ey^��k�z���^��}�_A؇!�I�i�RI�\d�(�+�#ʏk|7��V����������<P���bfG��Oĥ���L�����{<�k���^�UG|���U�y�9�����O��Ah��k���q��7�K��ܹ^�Yps��m�3x�k����#ʹ���~'���/1�yb���Mfv��9Y�����镰B�3���5�=Y|�X��C*�+�}��A/�|�\͈�%���L��n�K���~�8�A���ƨN�D�V�Ģ>�чv&�ÿ��`mjg0���?k��=,�~[_1����	:U>U�p9s^j��wa:����� �~��1��+)c.pq�Jt|lto��:�m�;�R>�hx�\�1�;��,b�y���(�*_����q�P�ﵕ^�W@��V�E���SM������5L;��ި�Y�=�ò�3�-��AwZ���L�v��A����m�D�ͳ��V�5�LV����2�\�$�{߁$�P��7���l�"��o��a� ��gfA`7L�p��K��� 6-'�7����I���)>u�����`�]��]�U�>��s�`�#02�@�;$OB��>ɩ���:]Q�t?S��<�E��N�a�UŤ��!�Ŏ����=s�I��y2e�?F�� �_�*��L��=,����;�A|C{� ��m��|^u��a�ӹ*sg��Fʼ��08�ہ�Rd<�} ����,�Ԋ�~���A`×=��ˁ闑o��2��Ϧ	�R3~r������1��{�9}�>�P����f���^	�,O��bg�ꎫL�%�X�e�k�Z0�+�xX<����7������͢�c��ĵ� �9�s"R�^BOXpWf� >�I˖����!d����O��Mr ���Н�F�&������F�D��l!�|���*t���;wZ:w��;$�e/Σ�R.D��Fl��:��st��r^M���3�q�i*C�3e��z�w6�v��,��K��g�M�
��'��]����d�j=�do!��\B�oGԴTM�߮��V��F��,�?���q̠4A��z�ƀ]֜x]���gLFFG߷��W�6�;ʪ�&�ãA�`�A7(�s{�9����f�8�uP��t�7�|��,�ĵȃH�<����w�u4�M�������\�_�i���!C�X|uyr��59�"����Q]5~���'�c;��4#�
t���o���"�4�Ee:�/t�S�|�IJ���4�G�gᵕ����1�\�ч��o�5��%�t�ة�3����'�{�
��o�˦��x�0F��|Һ��S@DQ<�^�P&����tih0�T,�����L��s�wbl,�0��Y��Z@��S��M����&I)V+\���#M�/əϮ�ɪ��6���9W��]�Hy��tnC����U�Q		L�o1G�7�,!]�Z.��$T�GO*$BLP� �$��:z��}���c�98���S8T�1,�v
$ �kn�Yh��AF���$4�͘;�;�Z��#�mUznH�^G�}�����ʀ�����[믔�G���Y��P9�|�ڙ_�m���>e:K�r��I�t����`m��a�z���>9U�~��!�W�mv˶KN��q����L� �J��:�����o�!���[���x��\�UCS�5]B^a-�p�B�ԗ���m�h��'�.�h����Q�0L�ƕI�Z��Tr���h0���ϛ�$e���7/VH��8]�
ڻ:����v�Vo}J^��/�B?�	����Y�G������L�st$�P[m�q��
y{�RYR�Njz�������K��L95n`5�sD��&���Ŏф~�ʸ���ߺ9ǻ#�b����q>.d�c�X�("�P-ç	�d�L�~B�8Gz�cή|;�ƅ�����.^��u�)m�̉9�8�k���p�^��X~z�R~z�$�_J5B�}�� bH�O7�$��~�b#�Ӱ�$>w�$�KR�|.w��=8pr�`8rX�D*@B��m�ON ���u�ܞuNb�!|��aHȑ��co@�į�+�_5�0?y��S�M���NLi��?l&k���,"�~S�u��x�2�H�C6702��J)l��]|��qO|��F��Y�@�pZ�N���|�yN�b`��>Waa��/g���0M5��	��^~k�%s�2�znf�T$�_��Tj_'�?�Y�������o5�FQ�b���C�7e��$�����~���08zǘ<'���� ׍�c?Yj�����? �4p~�>�`�>YӶG�w�$aaU�%挀&��uN��f	e�ݱ�E�Ԫ/"�߸w�B�X�̫����TX�)���4�<U`;0��=BX,�Ix�:+�s���p�%��)���Z��$����
��g�k��E�b���5��x��D�^���a�+�v�˩ax��,�&�����{J0��)U��[�R|,��I�F�.}���&�^ ���̀�\C��^�vʀ�5�R�����r��%�hU�{Z�@wpx�4��I����6&�v�p���9�K[���P'�Xm�.#kQǌ��1b������MJ,|U��O60T����F�B�g��	���H���xYPOk�p:rlE�ϕJʸ�����u������v'V�˛���r+O5�ƣ�m;��1}�$���?��Ӯ�����@s�} ̜n+�ǫ�#�]5L�g|v�©5���	E"��n��1�
��ӵ,�_����-ת��������K{g$�fI��K��e��<9�Ksa�ã��=����n�u=��|�߂I;�π�C@y���l��ʊ����N	0�t�F3�����������>d���o1������p)����|��WU�	o�f3��$xoE(�?z;�(y�#���]M�s�M������8�(��Hx���/��� �:��Y޽T���bc�c�_Rі�a��<�bad�f���9����A#5��d2�pd�Q��w�cO�_�iM���F�O�w���)R��07�b�����V�R�~�`�P&eH��r�!����*����2�?��0���l�{l5m7ȭ��V��'�ʪ��-�����s�����M���]�D�T5������V����4���;]%^�P�(��f�l��@l��e��O��ʅ�λs�����!=�Gb�i���_�0�!`.c�^rkHx�V�_��O,�qs�{u,����ጶ'3��~�{�AJ���������.+���v�������v�Z��	xKϡ�O��!@XiV��\���b��]0�BM;$���?]d��"��%�&*��Oa��f8"
#t�_�Et�#rԴ�Pp@} ���/C�㋚��fV@�.�v�':)ZXfU����MTu����2�^lm8R��o�V�ݑ�K@�i��h�5�W����[����Vp��<����䆸[���(�2�	�ר��}b�ƛ¶�cƙZ	���ڹܔ�&'^�p���L�ΖoM��p�`��6K��$�:�0J�cC^�:�6��QѷG�W��!�W�yr|ߛ��ۧE���Z�7^㘲ޝFr��S�S��.��7)�3+`�o��j�p��^�g��5�w���Ex*$�s��4?"��_��	��A���J���������ۊ،�CD����f�F6:>S	���d����#`�p�����J�2�i-ʝ�G�a�Qr����C�f7�Ol�zY+��
�}M'iN�$���P�k�:/�?l��Zq��}n� 81D�a��v��Nr����4sU���=��|�_��1����5��rcsݍ�h�1*�*l +����V�߼f�'��mLƮ��D�и�2���K0���LP5G-`�}��&�����5M'�0Wԫ��+��dm�_�GT�F㬖��OE�	��������Xel�OiDX-��妙�1��b��B!�{j��-�:��]�rƤ�Fǅ�_��/r$xتы3�9��4��'��I�8�[L�	�C��6;�#322 �H�6���������/���A�h�C9�gMI���p�F���KX�����],7R'�I�M�����;��H6��+�L��G��A����(m��+������5�)�����������h�D�˽w�G�7�n�,V�+�ktR��,����OҭD��g������}�H�lA��pf<ʂ-~X��-�^CQ����wsSn��	>����!9��"�&��h���܎���{��^����Bid���R>�EG��Ex�K�E�{��$�O��GZ��"0Wq�p}�����g�Rk!9��7h�Zߠs���ǅт�_(�}�	\��*::;:>�!dm]\TM�Ա�^<����w���<�&�Jv�ȴ��\au�:�6�ⴑ�֘�BJ�9���`��b���x�}��sۊ��A~��ĳT���9���)첊9�9��w��� ���Y#At56�d��VW<9�*�h@�B��NFQ�Zr�C��ܶ �G�`�.V�7�� �뜧���F���R����Cq�~��z~������,�>"�D;k�teW^�q|; 17�)�|��t?���P�M��EbZ��2�n=���K{��c�ƛl�<�,��FXԭ��� ���Z{��&����˲��T�;�vg7�(~�IrǛn|ߨv�|�bDC��yf��c*G�r�]���?����Kc���jcN�eM�[~�����t�pq`�Iv�]�f�����N�U�\��ЀN�.�n���6�9�5�Y�f��<*�H�@�B��T�q7�5]�/󂖏�V B�F�h�2!|d�m��G�O۰'�ޗ��GM*� HInP{Eeg �K��)��µ���XP����{��ʬ��-���/��B�E�ӛ2�F����._��+Zu;�'[ŝT_��=��g�mjQ�%#�f�e5�������Z��ˠ|�^pO������1.�7�]�#�ѿ7��~=y�[e�i�m(�p�ﵧ�w� /P��<s,$Iָ4�!�����rW�u:�P�y�_�G�=R�u�gs���$G�[����)Sn�3��%�"B_�8�� !OzWj��.�ﺞ�����ipxĚ�u��\�;�z��w�,q "7 �������(PCKnP�� �0m�Qɚn#�뭒	�#��V����g&^�Q��C�q���T}y�	��qA�LMK�~}�|�C��Ua�Ύy�jQh��?�{�)�,�ucn�I$������}��i=6p���^���:�����px'�N*"�'�Ic� �J���d�e�ʮ�����be�Y�l̞�E���Ix9�r�/r}sfm�s���3募��|v]��6P&}.au�d���X��s�j]�R����W�"���j���u���.��%�D�`��S5��>��l�D��'s����H�0�'D���;N����IpX�ʳ��1�&'�����S��.��F�pk�O��]m_N�̖.vJF�=�2��f�ga۶�f�=p)�o���W���n=��$�/����UF>�<ސ	���΁��boY!w�D�\L��輽�hqN�m�x�^w���$Mo��ִވ��|�/F[�5�%��Mww���5G��ko�cBp�KP`�|}4S=�jcU�|��"�xn�����Fz����Zh���V��&�n_�DD`��*JQ86�E�u<��0U5�>�}���tMBn�`�����L�����jQi�����P�)ؑ^��Ǯ7�.�|ܝUF��?�=6;}K�<��;�^��F*,�?�c}Kʏq�~SƝ�b/�/0(o7���ز�t4s����5Y�_)�4��'?h�P��e(N �,zp�R�j�@�?=	���$�v��vya5*o�G�M`{%���`(Ԕ��/�#yJd��5������fL��e��8�/���Ӑ�{ys��y5T㜦�#���$����rC��C���Mս� Rl�7���qd��y�O��Dk���q���=��(:-��SE��x��2��\��}����7�F�r��Y��m�4�{�I�W�!���	ggKA���=Ef k���5%5�� q�6㺁f Z@���%w���[TVZ�c$
�Hn��Z��x�T�V4�PK   ���X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   0��X��I� �� /   images/60733dc7-8aae-4c8d-a308-d0d87ce42cc9.pngL�eTTm��'�F@�������F)鐎��$E�A���a��F@�Sz�x}�9�s��g��i�+����'MuE\,
,  ���$�  � �d��O����=�(�*Ǩ��ޠؾP{ ��c�[����tU2�  �y������  O���/t|L��L?�b�}~n`j�����k>�6�}G��Ӿa.�x�дU�e���wEP��C�?��ǝWS���d2�b5_tbMԷ�'N,τ�������OY�ß)kM����e�J0x��[ĉ&G�yE����?�.��zddJq��3�s���8����Ɠ���[�o�~Ғ�i�cG�M�j�ެ�m�=�g]�m�)�iż�U��,�_��s��&bw)G��w�?;�?�|��wK`q#=})����f�?�nY>o�7{q1��Q64��@q�k�T�����~�y��ͫ7�^��K�Fq�sy���Ki�#e���꽽��l���L�M��e�I!��X1ˍ���,���
$r������Un�<�XtK�<�l�K!,�����p�~���k����@a2pt�r��t-t<v	�g8���{��]���jH��/ԟvNOH�g���M:����&��p��H���ڔ~�ω����z����ޫ:V|�d����.&UaE���v��G]Ֆ�}���iL����#?e�[}jD���!��qd���bgC��wmS79+Ӓ�����D���;���e�ȝ��_΁���"���p��ڪ�XՋ. ����'�((�x��9��'��ԚK�=66Ԛ>���v^}� :��2��s)2�-jp��@J�p�2QM���$i�,,,P��D1#����J#�l>�%�"�rŐ���'w�Ѩ1J�Qq����ʰ�2A�qK�b��<�?����W�)4�`�)2�D�8�+v��ҵ��$r����9�6ﱫ=ާb璘�:���u���x?�$�Ǵ�E���jt�
�\础��P�|�ÒE���c��o�����SN�W}r��# w>���֨�O�����ЁK�\��5&\\�o��AV��3��f��SQ$�8�������{�;#�h�����NL/�,��\�D�Y��\��xN��hv6�Ё����H�}9�\�j��R.\�[�}�1Y��
5�0��K�����8�u�W�� �T���j<�U�e��ý)�����Cd��IK򰙗��Po5�_ZZ(4�#��-������s�avU���̇��陟�%|ʢ6t��!m	��h1f��H�܌Zܡ�~鐗 �_��ԏn������f�||챃h�v^�9�a��5���R��������8_�#B.��4�ǃ���ms��m����t��_���va�&��zzz�&U@-�S$-��U�g:��ڎ*�����W}ӹ}.#ti&���~�?�?�u�U�ns��l��+����
c5��k�!�Ҝ˄>�=�����!Ex�byO[��;�[�?�����P.}��`����Z��޽����@�aA]���w��^K��v&"�{N~#^Kk�\��jn�sچ �uP���L�A�>"�`�v�� U�yHH,n�T�n�)sZ�q�m0�{�!��ޙ�����ox��/ԗ�m�*w��E�~��9�T�=Ή޻$�S�a�]i��СKrN#��:ӗ-�����t�p�����8xL?]���pV�$S�$��L�RYz~�1TG�%�X/XL.`�&P�`d$�sL�M}4��r�
%�m��~���������{{'�ݶ���嶩���???*���~i�����@/��2��>�~Y��-�(���Ǣ�k!Hg_5!�0�v!�|xS	�,�I!���Rg��S��0����A�g��PL`=I�QYÝy��O-[gfsճDK�VM�N^S�Q� �_;9q��|}�O"|=�n�����6{��e��v����^�O�7�f���O�G��Ə'z��X��'EAN�Z�{ګ�)WZn���i��ͤ���H��_Qf�!^���k1�ޅ��Aە{��^7��=�g�C壣#������fb�o�����wE ���1�(B>)&,+�A��%7E�S��$$��F���W�Fbcp-1u_y��lߍ W��s�vM��b.GGN�����NT{z�l=���nK�q�'�p���j���2�U��BP�i������͝ы��o�'GJ���-i�����&櫓+[\[p�%|=�uH�T���]�qɅ=~����;��ݦ�f�ⓕ�[�K�ff��oaQA󼑟tj�s�"gt�xK��7�Ы���4� $�n��]|��*�aC���\x"����a��������`Ƈ�2ʋއHi�$�Cr��Y��s��\Qx %5����gq�h� ��;�o0�X$nϤ�k(x�Z����!#ο_��d*�ߜh�j:�K{�����p�p+�=�9&��6����
��3��C�~�i6M�o�ŵU<��s����Ӎ0a�k_͞��:KO�����z=vy�Y�/�����-�xM�f�k��:J�J^��O�&���
���`BW�=K�=4�=]rf��U�R��X.""<pܞ� Nʀ�u��<j�ǧ*�k=9�:Tt����*x9�"�Te�F�f�=���F���/�2��y�=�wF_��hu]��;��^U[^�B+3� � �1] C5F������v	J\> a����|+OF��y�N�:��5maS���l�SÎ���o��m9�\�A��M�v�{�����2����G����(�����{��7�gwM�]�rłh�㾕��S���l�����{5�m�zv*~��q�]&!%[�XT�����3MsD��6�l5���Bp�{�B~9gˏ�6*:�T��X�t��a�)���RE��u�������|�BR�2����}� ���hU]ъ&U������A.��\�on�d�<�"krtD��ë������|�������W;;�+q�M�_[�D,�1��=�[Է��q�c?���_,e��

:Vp��d=�m�$�c�r)����]Z��hx7��R%+�m�$0�H9��@N�mO?F����]Lkk�������xtܲK�)�v�̚a�F�W4��K9-�
u��Y����$�M��!�V�~��>F���Q<Wɇ����/�%[�q(�F��W]�:8G�|�SB��=�� n�:�FF�=�^>	�R��tW!9��W�)����R����b��������i�:�!@�F�>����c��pU{�J����f6���^�+�w�Y��=�d��Ƴ~2�2���2�~�7�a�⸖<Ƣf�o��۴t��?����]V��@�󱜙��h��"qb�u��tVҿ����x`��/���Q8�8<פvQ&<�\�F��A7�5!����lq��Ţ��Ղ�8
F�3�H����u
8J�C���������X��[����@ڼ�&B����>8D�iO�j2���}'+ުm�� w�c�� R��w�?9�k,��\����KK�$�9p��3��,��f�m7hA�H3ָ.��*�S��h)�0V��`QzUף���pHk�,Bx��?00P8W�&�/x{Hw/A����q�Yb���z��ϗ��N"�A��5�㺢�)�W��\VP%��J!
'��Zi���%����PQ�oJ�gy�_㺢a���
5+%W�&xi���{���_�^
���77/TP�t�f�$܎���G��~��"��SW#����/�EYP�ڠQ�]�Y�@��Ѹc*�Ĉ�N��J���I|� �����j�^�7\M]�!r��͉��\�wX.��H"ٖ��A�(����X�Si�u�gPY�\��Gb/�'5���8����j6Ĥ��*�&�j�{
�q�jr��6�Zu#\Q91���/Pn}V��2r�=�1-�b��iE�c��Z��%�:��u��������(D�ʢ��ԯ��Y�`!�xz�4l^6 }O�"����^�=^�,VQ�����+���|qC��=���,\�Џ���W�Sa^�5�b�L�4�,	�(�9�`{�ͨzj�q���k�螧�ߩX^�(�A����e�^��S���b�t��W��a¤�uQo���5�u�N���7"�f���}f�����W�D�K��4�P��%�i1��*�Sn��!��hQ��D����h����������$��<�����O��O���_BSu|�:�y݇��*��Y
v�1Ƃ&�o,����{�RD�kjP�Q!O�ؚo�%#�$�Ƒ�.$v��0i�Q3�}���Ϲ����6�w�� �Ba�(�̤� �;`yAb��LvX�^�3=G���d��NQ�ۜ@u6#�Ȭ���F[�&�
�:����u����4��ODk�A����5w���%&�ؔ��OO�F�j���6�g�"R��1���hE"��r[5����4������vz���?v�=�iV]k��=�?���\�t(���_����G�nŒ�I}�v�M��Ac�^]���,����-����͋pH�ޠ Q'�y�T5��5�����e�"�W�o��m�
�W��b�SR~t<�-͟�m����8�:g.����G!�J��[�V��1'By���dV븹Ϙ��]׻��W�;ҳG/Od>��a�Id�I��ʜEs�T%:��(]8r��N�<�&&M�&��]�����^��]�fշM;���a4͢.�a��0��9ۧ��+��55A�^��d��F���+�V���'�����'�j��I��G�F��)�WzM5�H���QI"��Z҇�����S/,Ģ�@W^�A_�?��y`$�E�ʹ,}���C�O�LS~�u�c����M�����?���+��'	8u���kNi��r�J�xrB_��P��_���/��� z"W�)�����Q�I�����Ϲ!q��X�v������V��(2��s{H�"�-���6�f�D�8'�^�ޭ��vH��A=N��Z��z�c�X�QLl��.F-���D�7TCuV�"�V�� ���t"�-�a�����4��M���׋�M�o�*�W#9R��Pe�w��!!��F�U�OBiޟ��wmph2̆��p�Ԇ�����ekH�a�.�n��X���q-�J�k5��W���F���;1�O۩f����ц�d�A��M��aX%���A?�z���]Ώ�x��p:�밍�_o���[3w��o�MR��P'��?&������0uo�y��:��he<��_��}fhm��8r�����8�
nmG5ߖ%�X6n��酃D��B�>�D���<��U�þ����m��iqR��#k,W愈T��n`R�v�&��NR��*�ȧ��!T��ʥL)�u�ds�8�V���X`�w&� ��	�����棎�? � '��������Xˮ��D);\h����^�`�Z�J�&��0�yE=7�>�I�M/��7l�5* �1��?	6�y�9����xi�7�I{��,da��-x[o+��*[#�����w�=��;+)�oY��Tc9�[��u[	{zg\�ʸ���.���5�������A�#��������3*�ŝ�����0��.F��#����G�}��=�r�'�����>h�B�����#���~���y#��.�w>t��3��]:��s��[�4�l��;'��:>/�-x�ȋ�W�$�����Ē���Mdm�� �ը����n��u��Z��C��Z� h�A#.��W��x�T��~i�ؚG����6�wQj�1�II� v�ݏ��ԫ:o����w
�����b�|Y����?O�'�7���#�a�E*^\���r���8
،!��˿[�b	߱}/���U(�&�����y-��Vu���ۅ��r������r��;RP��4��Ut��H��xnB4��yÜ���Kt �����R)��}9>��5�h�����I7�SL=_�^��|m��X��u2R�C���v}�+�9*U��ai
�Qq��7c�f�A���H�������a�;����D!O6�F]KTۿ3�-�t2_7��C+�����g�{8�f{���S�v���s% �i��:��"�\Cl�C�Ԍ
� ���t8�6`��u����J;��s��^��T�L����W�0��i	�S!`���D����C�	R����wPl$��1���u����L�R�Z�K�����:���H�9��1����Xc�����=�BP�T��XLlg?�%�ǹ�ۻC�`22�<���F3�������C�Zvg-p�[������c�Ԏܥ�#�K�UUǺ�j�m@�jIY���'�����;�P�:����r�Z�&tf��|L.:�Pj6�E��)��ղ�r�n~���'��4iR�Es��ϰ�:7�� ��t�PuU0؝@0�&H����m'��^_o�̡qC|��`'"�%p���\��c
F�S
�����8�V=dP�%��e���2�KzѐQ�(э�%�p{���Q.wp�}`�������6!\ ��'W�`��L�NziuQ��x;�#)��^���+���/a?��1P'ç7��oX�'�i��;~�S&Z�]a֥.������(�h>I�!�_���׮���J��vU]�
5V�I�����J_Y0�w�2s&J�D���@�6�*���^�i|�Fs��B�$�g���ɡro����7�Jr��: Pg^���e_T�!��'�[�Nh�pE]��p/c��9�����}q���9��~j��l��Ƃ� r+dh��cwt���j���aߒ��_/n�d��R�ן��g�0����)�.�9�xX8ms��pt�Jl.,Z��d��?�g�dD�����"$x՟q���S�}���ɘ�4�I(:X#I�\q3�} c�r_��+T��B��\��NH7���U?�����"4rϺ���`%JUy��0��ZKM��(�����`�:��~�2�ڗ��� �&�'��D��J�8���%� ��Yir���H��>9�>���o�@1�:��11���f)���7b�k�%o?D�L�#�İ���+�Q���1�6.!C:m�����l���Vb�7�.���#h�x��6�_2�s��� :g�,���^Uv�H��������p��("`z0�!����~C�:����x��$��ia�Q=�`0��%xlQ5�2�qwiT0l��H���G��k Հ�A�4Tn�J2�y�(|4k�it����a�ïVB�4������j�H�G���T%�p$�K�f#��p�,�|�L*=�֝0EO"L:נr�2JO�vm��zI�f]!$۱'P�	e�� b󠑰���kb>7��4�ͯ]Bs�#o��@�	�3N��F����؄$�:L�xC��`j�%@�����(]�"��qU��NT�^t�C�
�R&��ȭ4|;�%�֖8��[6i/���3� �ۯ2�E���-fR�>G�5�#l���
��
��؂�a�dje0�����0"S�!&����éSgۜ�*[�d��|�@����9k��%S���S����d�q�łC���ֿS-�*���I���y��#��;�Wp��݆
�z��̹g�>BZ�{cz$�q-�^�xnoc���u�s�7Z2�#���sp���P��R��-�?߂y�����'�P���fw=Ȑr5���ǈ�G�����g)�Ӭר{Z�X��A��Lw�y*�dIE5g�_G0',�_~�|�\qkv9Y����?�r��8�OGa�Li��^�Y
3�����ku���>�]g~�������N��ߡ�xa:*�;�,��b�`N�Ѐq��_�&p�?�r*�;�[_t�u�Io22	��'��"���V�M��Y����Ͻ��$��N���?�ݜ:��st|��8�pN�&��|C�_.f��Ew�p��d�qR×k�RO~�Zf`F2�8[���v����-�[��;(��~�r4O���'y[`�����A���H��!�1������}���~K@V��m`��F=ً�h����?�`ۆ�o�D�i��%p4IGrs��L7� ��⋣�C�Թռ9�4k@.t8+O/�c�O��]K�V�v1�p�|���e��o]|s����-�9m٭���'�3�n�ٝ
��ѭ��N0;k(ʽDߔX�>�!�	�R]�K��0t�q;������������w�.��@����+�S��_v/���-���K_�ߨ��`���E�ȉM��9��^¿Z�v_�Ԋ�o��*�+<q��6�"��W���s�.h�Ts_��v�o!�`7��=M�F��9��� z@oC�yg��~�q��(<]�������x����M�0�� �G��$�v�� >��L���%�����t�
[A]蒒�`y������V������>�*[�+�Ԫ�.+���Y�q��A�E��f@�l>���rz|�4� -)��g�.���
��̂ƝiTu,;;�7a��<]g�ZR�y%1��Y���z
�����{�`����o莨��2���|=����קb�rO�W�Q�ߙ�Ե�@Ӆ�G��9ѩ�F��ui8�n�±�\W�E��bM�/�{[X>�y�w�s%vC���cj_b�U�D��)�-oܱIqc
��p%�K�q��.@i�q�#+��~�V�U�ב�*X���e(�eVA�˂q��Ʃ�:`[��hnK�=�M>=U�C�u�kͰ��nE8�ǋ�qs^��.*<���gkB��7�v�`�z�Hd(�;o饊J��=pm8YJ1 ��wzj<G��܇rί��h��T��0�����������+L�D��n����[h����|K���q����/���l�<��#vy��=/��Il�,'��ccfha-L�7ffx��R���j��!a�ء�S��������}���sL�g���{��o��r��$�V��m�]ͻz�#�շ�^z�y@����Y�Eՙ�D��h�ΩQ�B����m�B��go��H�b�l)���.�ٹ��QS�$�kn�8A����gy�V�T��$=2�?��UC���O!Ve��HZEIt�{�#;��*6L����G!���k��^�4�:{UƢ���)~'���I���8f>/ktJ4u��ݾk��u�=���J��3����Qi�q/d�d/	J���f�H�27�.l�]b�V�$I��n��lV-(^Tj��I-{h�~�.>�j �Yͫv0ۧ�~��P�}B���l���E�A�_�Z����6Ϸ!5ye�N- �Vq�A�`����+�Ch�'{�ǭY�a
��w3?r��W�l�Au�x�Ҫ��V�]�¢y�EC��*zc���������;P�*-�ظ�2Yj?���x��Δ<ZQR����٦7M��7NW��s1±5�r�� Ӯx�-��CZb������g�p+J �Ԙ�>`ּ�_���D�QD£dZ<L�p�Q*徇i�ѓ�>���SϺ�s��*��W��@6�'�Vle���{�\"��c�"'S!&�s�q�9�X����N�W3.w0t�,�6+g�"�glk$�ci�@�I�Y���yt��Ȫ�&��������z��cW�E��{��1�(f�t���t�Ɋ%��<�
�V���g!���ơa8���>����6Zc���`��s�J߰�<�Q6��1I�º~~{�G#�zVc��RCRT&��"�P��_���F�F%�G��&�kYEϚ/7GX�=X�d2A�\O�M��/S�Ԙ�a��|bV_TQ��?cD���FV<��n>\�Ҿ2G�S�vj*�.�^��ez�$�zEa����<�Ѥ��*)�_s�_��E�4Qԯ�Y����Xq��C�a V�c�"�\�ޗYkY��=TG{�A`/���b�h��9�:b>��<TI�ݫ�}����
\E	�d�7kunxs�Ŝ�[Q�K%�wꧺ�A{�s������!6�r%��ۻ��37!|?�<�4�F8N�6��hF6��o�5V�������"�| c*b5<���0��60���^0M�\Q�h�{�tPHE��m0T�}wE;M�5����u��w>*ұ@�h,�T��.)�Z�(�D�����m�SA�l&��p�X�N~�q�N���,,�ɨ��W��l�ٝ�>�ϟY��"g[?8LI]-m&������ΐ�{�R_��|���QWP�ĉ��O"�R��#��y�W/� ������qؽ��+<�IO�	�w�]�5?o���ɜ�q|�S�}��7��y�`#�П�Whg�Yu�B7yu������8�w�l;#k�D �l9Ĥy�^��0�ѽۆ���=3��RJ�(�,��h:*)9��E-�S8�+��Y�Y����C�7߆��xS��jO�i��d<�m2�Gbi؛�x�\��;���׉���L���*5`�.���䱭�<|�����a��ɒ?��NOOf\/����;,��V�dZ���EܮB���pn��E�}��.rt��i͎��������a��P�?���WTl������4^-`��hL6��N�K���EC�|�vlև6,��19!����*;�zђ�!4"w�D6���M'��������W6��ptmB����k���La�ʩb5�����Ur�O��h��gP{��d
O�-�N-���&��T&���5�:m�)-K���A%��~0CsN���Y�,>
�M���l�XWcW��I�|{SFB����-���~[{oP�L���J)�-<%4�?[��6k��zSK{*�Uy�Hi��ppJ����n����,�g��0�hf�;c@z�s��솹y]�9S��̷��*���\�ʭs�Ϟg�|��ܔ����4�H&"#<'��_�Cc�3�	�Q��_�W�R�ω�w6�ff�t�T�i+a�V�C��d�I�Tz�m,.�����j�G��?�W�r�=>(��G���FqY����C�;����=�&�be���sg����}g$�y�C��S�Ƿf�V�M�x���R���<] �|��8�.�_]V����7�'���$��@�sg���Z�(�X��>�(9DX]Q��Ֆu<	����0
Oٴ����}����Cu]7\?��ޕ�C*���0��!�!H���0<�~�ǋ_�h�����~Ha�=��|W�q�����Q��)r^nrZ����2N�[�'wo�_�"���'��z��o<r�-qH" ��>���`l���U|��黿���»&��W��e�D�-"p�G��T_���3�s��p�J�WN�׵[0�����o�{�f�|���?[%u�Ʒ������]|>����e��V���+�%�N����[eM�Rn�>Q�ԫ�����x�{�}�iޯ{�I�M�Y3�k�=<"t�]fS;�ə�*:i�r�L���"pO�R�Y2�v)��e
;�v�)W>��V��@0(eNPN���a���h�FKN�X�J���E�K��/�6T�Co�a��S�G�+�A�{[��t���A}���r�PPc��p^�E��:����i�ӱ���0��ќ��{:ٲ����_'�\�Z��-�_�'$��!�ӻc�MJ5I��Mj,_ݚ=�>�Vp�ɈH]��i��72���}�l�y}�~����+�p���q�Q�g�-_�Qe��x����ɍ(�3����E��3䝕��i�m�D�P"��Ȧ����谁b��Y��ݕ���e�h�1%��]i�-�o�4�^ѿ�����?@^�z����ac<��5�K�6urq��D.��-�ۓ������/�L�k�#> ���p�a&��D���p�����~���Aǀ����ue�6 �:_���n�|\&�& �����������^i,�*#�S��� ����������Oh�Z:�I-�HM�B~�O��^�x��^O{�օ;���e����Y�uuL�j�
�)��x�̤�jl(4l����?G���L�۶�c�j|9�5!0��w˩>OC���J�F�i2����v��f�,�DG�xP�x�0:���3�SA�g��@|e�i!��c�6�������\~ �CxV�_?��@s"]�B@8Y=��"B����/���Nu)Q�z�Q��q�����;���N��
IGo����&Z���[�;�䏘=��o��1�~�ng87KJ?Jc�����l�\aI�i����˹�k� t�k0B6��r��æj�/m���tN����?�*�����ʊ�4�ɜ�j�5��؛���Y�T��Ƶ>�J�cu�\��b��8�����K$pb<M���j:��5`��Ks:�<�jpy��x��9�';�u�)t��4�,���Xޝ�����l2���=Qs�iRI��Ʈ�H%/L?�8�Ґ���΢ξq�-�T��D%{��S��t��6-�c{�v��!�>�L��c�~�s��7�)�����/d��?Z�Г1S�N�m1���Z_ ��|�
T��q?��̥	��.�2��bF�K=�0&\�UϾ���t��H�3�LK0;l�0���4�6�6"��ΙWǴȎ}\�����������v%�$�n@.�modo9ɨ��ƚu}2:S��U`e �=^KN��t�y����y�+�����
���V2�������5�3H��{��&_ƀ�)[w�<�xt�/���3g�O�5��Q"&%J:6Q11f�0ς�1�a���j`����1hz鈖f+���bc�ҭ��vh(w�T���i_���9�sP��P����b�8-r#����ͼו��ipۂNW� PRf�$��*��CV~�ؽ@�9�����ҿ���ч�$�D��y����y�z��^�6�u%��ƣ�X����އ����V'ҷ(Ĳ�϶����+��s�ڞ���}�l�Y.���g�6"��Y]�!����Dm����^���э�dL��2��6�Y�@b��*����t5�ٺ����:�N/n,�����
0�Ⱦ�_$�y���d&����ra%��#�:��hD�Գ��_��{�М�H��P��M��n��;�j���!EL�k��=K%�;]�KQ�	�I�[�3�%=v��=vGΞ��	ŃU>�b����&[1w���ޯYSY+AT�Z�!���A�71�`�V����]�:��������b�� !G3���e��ԍ  -��!9m]$�@�+8S�$T Pe���^�$cg����|c��\�e�K����/��GB���@�9�����Ԯ�_���0��N7+�� ��x��f�yf&���3d�t^)��-;%�hq��[����p+����kQ���죽ֳ���<��G�{�uXP|-Q�O۰�h�I�ԇ�R���a�k�^O����]'���)�47v��7s��$r')� *�d��Y��ݽǫLs�T�?2��CcA	�X�Z��hI�@p|��doUܴ�=��}p������~FU�m�����]�W���M�gRl6�ҳO���$�����^��$t�6X�eE�)��A֩͌?՛n�,H��F��Ln;T�[e�oK}C#���Y�+;׊��k�Px����Qu�;f>��C�.+�葜�G��ϔR&	�̮��\p�Rf0� ���"�UG��(t/_���������z�߃������nA��-M�N�&.M���e�x���w��!1���Sݼ��&����SK2���G��亴�8Z�����2Qd�U�c6�.&ހ/� �����F�0n�as����ੇ���:�9t���DC���Na�I�|@/�$B�R�X��v������ٷ02+�|w�5���Oc��dɓ�R���"��S�&
o:��ju���:|�؟�	�0C�L1����
�ul�ȇ砪1?2��w�|9�d��)����P��9�t#�h��g|)��<^������0�e���|����$�)�Wk����	]#��~��A�g��(E�6��cD����R��2���;<��$��x�a+��b�d�f��2��#4���?1�6zZbeg����I�j0�};���?��x+�f�����C��Cc��o��`����74������:^��˿���o�Sv4�D�+��)Ly�I�ӈo�D�-����:a��o�d�2��4g�D�/��ˊp&f���c�E)�nϿ���E7#@�{��>�ڃ��$"���p°�>���j�PH��`u��������2�@eM�����-©� ��ڻ�d{Oޜ���~үM����h%-�s�`v�1Fp��}���*?�����fv��Uoa�[P6�B��?���E1�ęM�]�J�&�Lc�����$['E�-�--���yC��@�	����M{�4e���(=�\u��Wrޟk<j�1�D(��v���H�xO�:�ެ6{��,��������U�q��z/��oU�	�#8�ʢw�p�흏ҋѡtEzH���L��w�2.�iܟ�ɝG�W�*��r+$�)r����l�Q�ߥ1ǿE��U�m���Ku,KlQ��b��hAW�X�iP(7���>lqVf������r.�g�_�G,!?�J:@�{��˾1��f�����b[��D���U��6��тu@��+%��|�^���ixӫ��#EU��s�0�>�:$��y?`��qG�����a��ǈ�����A��%Ѱ7>���Y��GQU����x�f	fp�{��YS��P%��v�G�32�H�X�p8bW���O�9��fj��|��������y�o�>5�2v�ޜ1[Q9�lF�D�${jQ�e��|P;P��M|������y��������f��R�C5g^�3".�9fj� ���v��z�r��8�?ewxh7��^��6l�w�G�����E���sp收�T6��Y�!���H���D�ś�J��L��n__�$W4�㡭e,c�3*A�&7�;+Sd^��JZO��k�X=G��W��]s�pq�-�pt��袰�@��ۄ��x:xM&B./�����1h�H�0�FȪ�T��ϜJ쏿��r�l�o���3� 1��C���g�iь ��1�y����d�S��hd)u���x������L���`Qn�|S>�6��)�"�d�8�����J�p�c�ۤ1�;��#�r��󀳖��"�!��m�w/nݷ9`b�l� �d���a�� �h�J��:�pE���
�_��w�CY͗u�Sć^�㍈���n��Iq�c�7��Qu~J�G<#�di�&���>޻$oT���Lf�x�NP&A �v�zi�
 p&6iv�����~�!s�0��#�����beu56i�C9b3V	��,��Z��_rΧ�3�<g�aZ�E._���_7<�H9?Y�P������S���{K��d�g�7�h�H��o��Bౣ�Sk�_�vS�A�������J_����{�V/q���~��=�=�6��n�p���t�Z�/�$��{B�z>
���h���Fk����\^{sv�hDp�N2y��}��-�'W�pYjRU_�����W��|"�s f-\���Nb�/$��G������	#_��s!�,����h�2;���U=�������x��X�U$���4����D�C{���k�~�I �mD�='6h�e�\6�	��Yh�vYh��}�0��i$�o�ڎ�����8�%�~��k\_V,ɖp�c{Y�ܤ���jAxUk(cyNiT��h���4�<]i����T��Q�M��B����CW#$ �ܳ�kM�ع&u�4�a��X�#X�<v1�1}�b�����5��o�&4��>��%�����l����%��Q��hyyZ��l��.gs �M�P� X� ��&��gӪ#~Bs��Ǐk(Ḡ�q��,|�l�����wо��|F��1���E������z�q�q
Q�����Ѫ��|�ʃ�,^P6,̝F�����Yl\���~c�_c�7t����lv�0;���P1�Nw�0�L�@6�<ȅ>�q�m�B"��%��&�	�E��m�6�\x8ZϾ�Hxo�Fk��� ��&%���W���ҙ�3�Isz��z9@ԿQ�}8�bMn�	��zp@�Y��+���Y4�/�qbBp����/��b 0|�<���]��3��+G�L���=u�_�}r�+1�W9����\��S�pi8�Gc[ (���*�6��f�'/�H�(��#��Ou̍x�C�(Xk <����f��|1iU&Rnc��8~�%+� !\(��pֹS�X��h�o�C���9��H��ևI��z�ۮ�T=�.�����	��ܐ�L:��~Q8�����D�GL�[#Z��+������m\�6����e�Ve��no����yb�� -@ҿn�	e?��X���a�w�ֈ����{7��o�~�9�v�\h4Qo3C ���ȕ��MƑ��e{�t��>���6��g>�h���â��p���_�p��U ,���M��ىf�Cf,�3� `>�¶�0�L� t�5����SO=��h6�w�;{�f�ᙌ�Ge�X6}1�@eN���S�C�"���9|�Hڻo���M�0,]�Dq�o�A�I()�-�`<!��� ���թ�������Ӽ���3WI�>wv_�u7l�,���7���J�[QEUT��b,f��Q\M����r�֎���
,��|h	��W��g���WC�����(c+x���\��(�c�����9��E��
���'����3�d���P��Gz0�a���}Hy%m������ S� ������0EqVs�,6����� E`��!��3�8X�4�b�PS����O����2�` �~l�c�a��;v�p�q�W��Kٍ'ʖ4��7JT��b���\��D{�GoP3�*@��j�pF`��
���B�P*�����5A0q�+lY`����L�*�{��gң�>� �!�-�����ͷ��>g��u�ܓ���#@��K��H�[�Y�0Z��K�f	���w޼���q�F/+ ~9�P��n�
�bia�~;�U%sTȢE�v��2{�r��j�8�߄�����M�4`S�x����0P�Qv� !ʸ�C�`����c� 0�n�����=O��'��M�^~Ah�Ǣ!<�C9WTQE�}"�Q�@����d>��D�g��G��w�<�X\�����;;Ơ|-;��D���O4�*:Ľc\��w �1��P��S㐯����;��k�7ox��0K�Nc��@K�]�|�6�,�ww_L�O ޺�tz��7m��r�q����+ȼG<�c#ʝ\�Q�Q��j���˺��	���P��16�w�5��B�
�`�����Zgx��10[	�XUg5m�%���&8�16�< �S�����:�2����9���c�J�M� g �9&Wx#�9���kV͞33͜1Mة?�4(�P�����mq^�.�c�mv�?��`�oJe[.��(��#|��P�a�+��I6���3gө�gl��  ��(v!�u~�~�x����P}�ް����/����[�̠��'�`?��`�� |��]�beڨL ą�c�A�� �ì���W����L��MeΎ#�u����\<�Ә�vf�����?��'f�߳~��.3��e5lk(|fQT`�8 �\�!~l��W�ؔ��أ�h��ͥX��(�	�����1klmmV����7s�>i��vx�7�����q p ^&����_}\���"��y:w���<\��G�'�=�$W�?�9_����w ^1���~bwwY��,�g����Y���x#�D��+~�O�X~���.�K�>�@�,�� �e�4�Žw��\�+ ӫ��w��� �� 2�>\�a�kv�E $��h�{4��X�`��CW� ,�S{Oj�Y��+�������i[D��(�±IL��� ��R8�l9G ����bˆ-�	���v���t��9�_S����o���o���r	m$�6xϚD(/�����m��s���oi�
W�M�*\�q����֬]g�(�}%_�����?M�'�N��V����p���SNp�8�5�(�X�v+|e���ԃn�f�=
DxGf ���C������<�9"�I�ݨ��+g�3���:�t���Ӧ
�N�*�Ac��`N^N�<a�4+����ZǶb
J~1]���م�O%�����.���W<��E^�`wjg��	��V�w�ݑ������ɴu�t��1wR$Ƌ��iAd��0�,����)W���O?�3l��[�����[�Ը9��tڳg_��K�h�qܕL'��#��t�]_����DL��P�<x�C�]��s�V�^���x����t*�W�S(��L�ww�ޕ~����W^}%-P�jO�:i�r�~��ǔ�|�m�$���Pxp��"��ރ�nܵ��x��������I�<_~����믥���8 S� �[N&��rT!��U%��� �,ɄIG��b���8^�̙�H:�9sf��b>�x��{�a�*�����iLG�&�)��~��DW�x�����qC�w���~����]�w���{�՗�w0�Z7���.<J��}ɶ���)���A�߶;S{�M�" �ע/�+�Bp�=�d~��
?ލ�M���s���~J���y��vE<����= U�����>9�4������m0 [��F�!�����*�7��?�#�J�����G=����"���4).<�E^��pTq�3��x���KLʫb��T��^�P�N#VK�rr���/��D�3���7y���C���������}�I�K�;ք�^�_���O��G���Z&��
.s�a ����|B�6������~�����4���o �o�c/�8@�t�W Nc�E@q� ��4eJ�q�x�>�~�k�u��3��S!�r�E��K�������u������˖�U�>��Od�L	 �(������ ���O34Fck̤��g�~�s��ft���| \������T0���%ą�d��~L��/@�Uo�%���4� ��8��t���ꩣ�#-X�0�߰���3fv���t���Da7|U)������?�d�ma�i�������Y�x1�x�W���?����̎��2QO�k@(
�/����T���������^�^8^zB�������w��n��;�cF��-K�Tv��2�;U����!3g�b+���|%=��>L�B�s4�i�ӰSr��6�y*a��g�q����y�@!Ϟ=˂h�06�������cGmG��f��˗'Ng��ˍ���XV����ڹK ?��Y� ^f���,N��'ݷi�w12`# �DC�_�. �/ �����e�`z�������i��eN�������`7���YnΥ�V�ߔk�j�����`�A�x���p����x�~uh�i,��_Y�r[�l��`���W@4�ӄHY@���3��)g)� ��"8�5�$.�&J{�Ϗ��Y뤷utF~WK��>Pd&̻������x��x/�'{<v(��!�"|qW��~~���{ǩ?B�_N7��Wݏ0ٯ�<�[���[�_��]2��{�ҕ�{⭁�ŭ�Զ��牙9�5��w�7�폟��~�s�����<�/�����{_�uΕ8i�8=�&�����-��WP��w�£���@#L��� ������|qS��@y�sl������dq)��&��d^D?e�hN3�ET�a�٦������s4!�]���PD������G$�~<��OCj|�4=��G��a{GHY#j�]���籨�ße�i؍�|� ���_\y'�z~3���E؆blCcl
<+]Ҥl�,��b�v�E�361O�I<��|��yf���(� i�_����e��.�O�6��'��H�V��O�n���:�]!G3�J�R�����������1-x��ɬ*@���=d����v4֜����������vs����8Y�Lc]�?K� >�w�u��+%N�����
���o�l�t��$LP=��鳟}��@kK}cV�ӟ�4��_|�����UT6q��|��!�;��{�|��e��RƀS���1�Њ��̢������{�θxE>��2���X��G�4��i��ce����킅�vlb�peߌ.��h����p,��Y3����@��Ya���p���ƛo��������I
9&L�u���4�R_��iS�f����o������۶�H[�mx�No���7Z��L[:�hPT(^,Q�X4��`��-Ό��o�F��W�lcmJf��;�}>���W}��}X���ʂ����O<�y��y ���h"o�C��J�!�$�j�����2���q6���Z6��ر�߅>z䨅����h|�mٲ�i��������I�$�ٳ��GC�$kO����o������^�g�:�	��c��H�
��,!]��N3�Sq�G֯��j�\'\��\?uGx4Wwt�����p��Q�6��eϷ��?�FB1Ȅ���!�;\�H�l����~!C996�����.ru��"v�a`e�a�'1��3�*�J|�3�;��xV���p�!���I�9���z�t$��Vh��G\xG�.~@��9�4{��9�ٿy�?����bE��1_'Y<�	��D�A]EI�tU϶r	���{�)�EX8����m��÷˻<Uܒ�2�7�E�䰺�y�m�Q=�b��)/Q^DO�!�q�[��!*�s�i�����z\�g�'��O��-L���^�Gzg����ٟ��~e�	��3�¥(�"/�/�^�c�/IVc��5�QX��<e��.�&˘��b�A��3xˠ	�wQv�	H�� �b�E���z��h���@���0,�B��1��b�����Kʊ�y�|Җ͕���)�6���G��M�+�w�Fc������_R6(	H�u%�y���wIY��,�ؽ��plAQ^܅��s�]�+��= eJ^M�L��N�(����r�jUw�-�q��E�<Y�ܶ��[s�\��]��.�a.jOR^L�ey���Ƃ�z�P�_v�#��u�	��� �T=�iȘ�T����l�)$�&�1���^����p�e"��2��h�*y�rS�-׵��퇥u��/|!���Q�����������/lN��)���nd_�T���YE�92���̤ϠP�`���Vկ��J��(�o�]�^|�'V�ׯ_3pf5,���=����L��'`�	���ɢ����ϝ������Ч<p���}�g���W�)?4���x/����0�a燴���A�2�W��/��sJ1^QF��;�c�.J�'?��nݺ]���jh���m� ��(L��f8��?����ҳ�<k;Y6O�qP	��|?��_�ȧ \P��YѲ��ӓ�y�ZU*�c��G�F�����Z�)d���B�����x��U�Xu\�B<��s�U��ă�`W�f�]� X�6�|��w`��A4l�#Cx���%Nޥ�,��6޷�F���?�gkq��ٿ���:�'afy�# ���#k�Bޥ�1B�]1��Q�Tat u
�zX����޿�ύR��A�/at�Pbc�\�����qLY��E3��Ι�ėA'T����?:]�A�)���< �� >���!�k�S��, ��b��8p�AR� ����nt�r� �=��\�)�,��e��D9���!�Ο��Ӎ:��Y�b�M�y�J٪�-�g�t�AΝ�e�8M�+�AG�2?���C�@=8@�'X�ǿVv�嗩+~Cؙq���=�/�Y��^>:|eE>��b���H;�!���i� ��❬2|PǤ{����������qY^I����2~F\I��y����`�߄4/��{�/��Ua n	�3Qg�cb����(����_N!��5����Qv��k�`R����1�.�F�x�p��{�������,�E�����L��ZR��u�0�y�U8��0��I���m�6�Aa �n�r�/���(|�?�:"��Gz�t̿�Wʣ#�gyBK��8�
;V�Q�!O�_Cch�(O�r������\.#9�Q.[�����!�-�IT��n�t�]C�~]��q,�sbrM���o��q_D-��b�n����mx(�k�JߗٮɎ�l�L8N����㪕��H�[�y��G"�5sPS���l����@�́�I]������R?��k�z�A���
?,o����\?�|�1�ux�S���eA���_��׍��ƞ�����?���@�U�>w=~�g�n��̸K~�\
�>���d�{����E���k�ǂ]����o�X���b�؍�E�E����.��O�� ��e�������+6ɀO��N�*L)�M���ݿ�w�좴�p��]������a���8X��<4��+�1�q�h�4�ah���4�,Z� =�ؖO��v�)��;��VA��Vrg���1�pd�KA������NO<�x���'|�ӕ�Wm"������v"�C���M�h@�p 4v-6}�4�q�������tQ��B�`�7�?�F=Ϭ�ȉsٲ�����r�'0��,�
'�������_D�����J����`[�t:�Άsf?|ɃN���_�K:��sE���͛��`����[ �m��<Q���*ڐqA�!ʂX����|);q�{��G�A��>�h��K~�)0��l�:a�̬-L���@/�7X�h2C���^d#����4<�����(yƄ��yFg�<��9�*��_�C�cn�z�͉�MhBB�I3[�/ޤS�� �yCDZf� ʊL���~84���0~�����j�fB <�Gr}Q�h\xr\���;>���?�p���t��8����W;��r�%���)-E�3��'av{L<@�g�(�%��ފ�k��[�N�np9�AoT�+������T1��Α�E��'�,�E�9W�į��,�t⺈x���`�N��/s�Oa��x�jH󶵎y�c"
 ��.9��O��?<2x;����w�?�ޱ��=��<Fx2��^&竐�ho�����\���6T�VgGq�G�;+C�t��i�e2w����5ƻȏ�(����s�|<9ʚL���j"H���:�H�|��
�+RU ��ќ]�r=&�z�/|z��~�	����/0�%���>.x�儠���6�~&bU��(~�uJ�-�G�QD<�c��T����cޡ��~5�N�F�Q���19 ��w�S+S�	b��F�_\�r��J��}�;.��6�)�����E;����(��9��6�}1&�_�
��+d�q��p�0���2EJA���	m�Ai�9�~��T0_c�<|�Pz饗���$>�0x��*O�:�}0q�y�"S��Ӓ卶ʳ�0���3��,�10�0ޑGlp
���r�<���f��?4��:p�c5_,�+��[�mPb����o��q`Qb�������������R�D~��7Iv����0� �R}K-L��m��c�?��A� �qD$7�J�e`��;���H[�l1�GΨ2��{�K�����~�z���B+�И�<��sF�hA�l~1S�} ,���L�J�]���)
��]�5	x��n��5|�% <ᓼ�Μ�s���g�ap ��}��i�=�UY�U�|�x�fMg|t�Be�������?�?Ӿ}{�q�W��_	�? �i7X��W�~�k�=KS%��D3�7|U4�L����j+"/7h�K]R~L Xf�@f�#p<�3�;'��ҡ0L,�_�p��aiX�i��<�ߔ9W��l�|T�7q����� ����86���3�Ϳ�0$�P,��ܢ�`� ��&�,�&���M:ʋ�Cdܳvuh/.5n/�)�7�Ӭ� ǭ�I�tR�G����q>�{/�	!cC�`LZh��'鄃�_�W�
�?��dzx�s��E�Q��i��0��(���ID|d���?ihPb�i��L��L���:$!RՇ_����i��Ti��y'=B����/>u �\�W������U��D�Q�F4����9�������_�wD��r/�+]�R�Qsų���_
m#�+$�tG��&˺�Ki7n;�����|��ۮ��Ekv��������v=Ѭ��Uq�}9������h�N�p�'^�0Tw�+K�^��G8��B�Хr�M]�h9p�?1�x�*K|���e*��p&Ȁ}@ �>���6꾃>�H����2�O\��2Q���U-Ҏ��� �p2qK��{n7Aĥ�Ԅ�������=���O�.�!�� i#R,ǡ����qqy;�¹����B��;n��#4��RԭCʀ �M�n͉~R�1θ��;�k=D�Ÿ���(���L����u��� �o�-�<�L�D�O���_�p��f��'�H_��W}R��i�<��������O�%��0�����kR��Ki���6Q�?4ȱ�P����-�p��(Ye�.�H�<���y��=�,⧌xx�R�s%,'Y����g��KڴL	���ش֦�������٥��\�u���_��O��j����3�6}�L�Ѿ��_P�s�p��e�w~�wSKScZ�tIz|ˣ�v1aغ��t���`Wb�8`�B!�UJ!�,ظc���0`��Q4Ԟ��;��v��?��tT`2f��A�$�l��[��?a�/@�����}a�0ZU@-ju@�M!\�r)]SA�� �/]��B��Fp�����,�2y/�������w���`��Kl��l�20�G� �T 6�����~;��c�������/iˣ{���B^~������魷���J��:Q�E37�o�
�w��#�vQn$��F��33��f9�s�i(h8[��
��lmHy�]�eF]c�h4�UG��#�DF"���]�\�\�N�04�h߱�6�N��ppͦ�)��eS����"/��(C�C>	�y�eJ]P�A��:V��@�����#�t�q%nb�4 h�ocK\Ԫ���s�'ow�"��۝\�˚��@&��	��y��9�qD��,�ٴCF�� Փ n��"`�o4�a~���sAFj�tH��`� o�y�k��wڱ��A^c0�����p��7�<{�)�����/���M��[�i~f�$G���Q�*gdм�W�l��6!����8��dv��r>��}�!b+��.(;��(l�~4�f[�:�E���탁r���xF�R����is�:d4����UY�A�<���`���(�m��U����ӄH�D�(�.�`���<���$�Y��3�sx�S�ߓ )�a�R�+� ?�"����4G*�b*����_�I��e�U��KݧN�LN��Z���1���r��Y�������~�#fq��~�a����_�%N��O](��	_x�Q�#���~ADYӷ9b�o�^���/���²)�k�*��}5��W�y�Ϥ}�����8uus0L� 4���o��p�#·��+�(c�/��o��?����	�J�����P��q���*>o{E��hi�����L1��&:\�g�$MV�j�'�%}v��O�A���]d���'_[�?>�Ū�|aN�Z#@#V�Q��^x��ݼ�ÿ����Likc� ?`���p����w�cW��L��LR����XUָ$�Ԭڣ�ņw����hv���w������]@N&�M�D�EUH�s��B��VЋm+��# �.��~���p�!Xѱe�c�'�4�rVd>��bfD�-g��5��1gkd����W��dր���0�J"~yϛ�3��|`�i���ix(>� |�/z�-�}f/�3/��7y�84�"8����O��������V��猱���ގ�����'?���@?��4V���W�y����]���7��R����x9ÏFI����Y�"��ԣ����� ��1�y���Š��.ˊ�<8�&�t:Zw^��S�@�{O����x'�P�b��ޝ��eͰ�E��`#��ehu�ꄙ�P���?<;�,+������d��◈�F�&�K���N� L�ŋ�p���z�?�AG\D<��
��"��N�}�˽��y^w�'q�x��Z��0��]�i淈Q7����B�[�јP_��ru\Q�<��C~VP]�̏�qu<ů2O%�g�����W�r�i��Z�
���H�e��љ�t["�.nMgHE���`.��E�XrT#��P�����U�S"˘n���w{�9�_�d��xj��?��7n߄%m�&p�,޵��A�eP�ۦ۩���W�[{�xn_W��������J��b��V��<P3e��߷�o��K���H��g���$�I5���^p$?ʀ��23��"bx�>.4x��'����G�go%c�p�Q/R����#n��y�h�I��rz�9�Z�38Ec9��IK��l��H�p5sxQ޽_~Ń�s�i��1�c����&���Hf�_�ӚP��1-xf��x '��B�2�%�H�e ~�y�����6�#0�@�:췾�>���d���o�����=h������p�&c%r��|��%�KF1�D����J�c�|�7�t�p�&�J=6ճ�i��|~/؀O�$/^�S.���|=p��` �������#9��#���/�Kz�������㨯�3�����1E��ǃ]VIV�n���Z��`�?|��y�sj�����3��K�i��#3\�X�MM��D�Bz�a�Z�%�f�Mgp߾}�=@0�zU�%U���,ew4�$l�z49p !�T�[�u�P�J��+�-|�ih��`�9��;'�Y�Թ�?� p�t8�-'KZ�MqN-GH�T��9����=�-�������z�j:x����F�������Ǻ�ϔC�/UN��P�u<�M�]��<SV䅼s��4I����.� �z�5���j�j\�E\~�4p�=.��&Mk��>i1�� �
_l@�o��3x�{���V� S.�/9ޓ?+�Ù����1�kp麉Xw����O�+<���R�|�GY�<��aO�1x��OnTnX2\������h�i��p<��8���L�u.�I�Z �!��ت��|�}���}�V�����|�7&-��0c�,UWv*_~�.���N�a�A��E�9��C�Ҹ#�{���}vLRp����A��]���;���o��4��|0a`�fZ t�<��"���R|���>���x�?�	���.`�&oPP�ǂwE����/�Ǿ�<�y�_8���z�:�zO�J��\��W�����a�I����	��=�44�t35�vq������^iS� M4e�&�)e�~�k=M��ށg׿�e�ز�\�!�5g��G�C����i��Ѷ�l"S!_�(�kX ��#��b����~�3����.����{֎*$e�ve�����9�
ᣐy�G�JI�CC
�f�0��2�ޡ,��p����{�.�7����{ғ����T��?��8Al���*<�Թ� ����+
�ˈ�O��h�o�D��!�3��&$ꏱ~� �z]L0��C_�x��,��Z�D�֮�٥�O��I�����M�lX��Ο?�����<NA � ���Q<�����`<�I"
 d0�Ы�l���@c��"���)�a�%{�P"�}����`�����~��{���N�c?��{��5 ġ�MD��PL���*0π�0����gL�JK>�j�d>s����^���-$%A��SY��=@��3�Q��$�e���
Ix2�̇L��=�+!l;8���{\Q�c_�Vae� M*�(����F�*@(iXPJ�&��M� ��J�=�,
MB��/�Z�afH������Xx��U�V�qs��hs�3���@{�m~�䟉(^�W.s��-,w�+(�s�!h4� �R�g d���M㣳�>w��N� ��}���i���~�ӈ��-��1՞i� ���,Kp��A5�Av�o6��q�$��T:��^ �p�$�L�/��3Q������:�JƵ�#�"j��H1�c����%g=��-�4At�r^��{9�x��O�7��``P ����&�2��)]0arX��^7ܛ��y��p/�jW�U��iP��Lc��7��Xg�kat�?�3����U91SF9��/r\�'���ePrNn��>M�8(�Y�_����% NhH�B�C���S�oG�0���*Q=\&�[��SΟ��sn�.�U������������)ǣ������Q��$��1��ȿC:>����f�������M{f<��g�M;�3ʿ.b�}�[�ոEX������{�xUZm� �?V� Y�<!�����0d����bmQ����͍���=��@�_����!��֟�A�<����sݑ�u�U�∫��_��E.g�㼝¢�O����G0c
�є� �U&d�}��'�܏#��?��h}��p����[@,�|Yp�h�"ǅ��&�7�^؍O�:ͫ�D4�8xf\��c���~�_H_�җ�:��(G�aj�q���/����<�٠OޭH�\��A�U�|4�m��;�k_e�i_�c� ��4,6�SF��.��/*+��:Q� �N��z#d��S�؝�i��y>+w޳��b�_M�V˲���D��	Y�'�5ͮ�s�"�[�J���ƒ
�.�!� df�X*�����0��US���0=4t��Cee S&������Z��'qa���
�}K����8���Q�T�	a!/5Gqp�ꫯ؟�3�`�5Zh�?���Ok`�/��r��]�����<|M_�K�t��.:�<�ġ�Л]�9-������^L4�^'eG�����*����"��,G_�z��O��n�� 3Xd�3.:Ru�_��4\ǡ��Ƨ ǣ����~٩ʎ6�h��N��~�5<Ĉ\�A��o�����.@ϙ��\a?w<�A~�D�u��s�����L��� Z� ��w�X"H��k�����nMc�o�59-���|���ℋ�+�尵��g������;��s�#dRS���o�� ����t
�i�ӣ	��}��ǹ��k=?��#_�Q~Yc��_�'���unۑ��;��;�-����w<��S~z�ߵ�*��/UpwYLy�]�C}3�~c���O�m���}�9ʀ�r����w7�����m� �CV�TÒ�һ�L"= ��Am0��ÕˋxY��l�S �"~�	����<r���P� ���
f�� �ӻ�d0�|#��s�0�vt�[k���|�!i�����ޖ:�v�]�ˈ�@t�M*'�8oW8x ��S�]������o� w����^V�p����Y�x�d���<�wΞ5۸��1�;1�`����x�`�<�᷀)�d�����G�l�h[�V���Ӿ�<����� V�1Šl(���v�ی����s�1�%�r4��ދ^��C_���yph�	G��Yf5�<܉���L ^���[ݒ�-]fy�<1��S��@kvn�nr?R&~�(T�,2V��QlR?�]x�`�Q�c)';#BB[Lܻn}��e��o<�P�lL� P�,Q�s�֗�"t4fYNE ����x����J �"�#9��Q�<�K�F��`4�}���eʻc�Tv�
��k�ǵ��0j6\��:D��/]-ȸ"���r���t�:�J�N����Qu�
�`���1Lrpf���N��Bf̗�FcG���q��z�����rP84 W�¯�
�r�1a���(�E�0.����8���|/W{��s|���9�����m_��rp��� �ĭ�V���I�w�Tr�>ޕ˷����Nd&��ǢY�!� �r����G���ݡ��ǹ��wqĕ��.��k������N���Y�#4�ug�!7��
D�e�1��*Os�u���N�yT��@Y�/
��f-��8&r��W�����Ƅ�?9����C�E_� �҂�+�$�ቯ���jQ���|�k��.���S��I!SzV��ᏻ�l��?�
9\�['x���Q|Q��5�ė'8�	���I[[J��4BNx6dX^�L(����?e���(� +
��Ԏȧ��| �"���}z����e��o��񶠐��������.(�;>L��GX�ʍF}�Z�={�֎�b܁G ��%���4�5k@� �d��%��0-@#�*6��Ѧc�F�Ue��p�E}�3O�^x>�[�V8j��<� l����U�{7�k�@9ǥ��	�J�����)���RVD�Z�e��I�� nʞt�غc'hgRDYQ��|��(��F>�����cⷯ�?����E���cɠF��2�C�� Q�%!�?�;.���/����Hc<1�D(0�>u���]�b���|���n�d��L�
��P�n ��rn�Z["X�2��!o�� ����W�^m���K%@�F�E��Mx�[W4��/���3�<y*�Ip�<�2���*��_o���	\��P��;_h��&��r�P�\L�����A�N:\G׺��ƒ"��]��h�l�o{���*�l8 ��)ҵ�J�Ҩ�+�H]pO���G����B�K��'Ax^kH~GW3�i)@��8CC�G��3~�U�O����.(\��wE9^����9}?�����%����:����g��3/�������E>�V���e�uzh�����}���<��Ex�M�n�����W@o9yg�k�G�'����c��O�8B	�B��c�&�_���|�|���D�0�#)�~�\��W)�Ov��_-�'�ݠCcV�p7A%�ap@7�}����኿Rx~��̺��Fv9�j�q��w�"��z��E��%	aq�p_�j�Z�Z|h�΃��e�ml�qJ��ײ?u�0��J�|�D��qZ����w�=�U8�����l�����A����^P��a����@���5� Oܫ�C���Tvy_�-�ۨ�p�O��l�H8H��A��hǘ��8>��[���r�x�eQV�>�3 ,Yʧn	O9`��xր����v�p�����������p�@�^lr�	�+l�w}z��l6@Z��~���С�i�������^��؄��cG�ys>�>l�S�?��g�H?t�:!ev������u�5��*6�ӆ�K�Y�Hy�٥|�\��|�����b�/���v�U����R������v��:����2���ۭ�Qi�x���5�?֌��0c8/�'��5lc��k]�� Eo��[���u��%���l��(ǎMG�z.r�������ѕ�l�� ̞5� �� ���݌* 3���&�S�N8N
�Y�O�b3��3Ϥ/~�K��^�IK�❵���hm�>�Оfϙ�.]�/Wl/hu9�� ���}2������>c�O#�(�X�d��.8�-��9p�����3�5;S�=�����\���.�x�e���p���	)�y�3�yNr|��m^˾�0E �����_�W�4��c7ȯU3^&D�/�5h6��J�r=K;�2nh����M�Z�e?5|�5�=rZ�� �#���	Bޑ 
���=�x�V�h�1�X�&g��ߤp��=:�#Ǆ��I	3��H���X�/c�W8�P�ć6�R�:3��ϭ�m�]áe�h$�+�Ba�ON���KH
�3|��;��,(u��-]���L�W e ���;�!��v���TqR8��,ăB�y����FyT 
&+��0P�A<.U�S��?�eL�Q��	ȓJ^|�w��Jz!��&�}��S���� �|���Y��q�J����>:���xl����YqaO���?�;�[��������P ����=��(�M<nkr�K�	��DX��ʊ�<H^q"��W�m��<�E�V����ܰ�6��q229��}K}��"_��q�82E��n���������=�Q0o���z9( �*�L!�7o��FYz����\�9�Y�2���ؐ�,��3��klh�C!,���3�P"�GĤ��5(�qӀM?<p�"�"�7qd��r ^��1��Ou'��Αf�)fd䓌R~޸+>�g��/�<��&����M����؜8����|����oݏ(/�lU��$��f'��͚&T��"8%�`��;^��@n[�UŐ=�#@n�/`��Gٌ�^ 6�c&�<&2�N�.�8Y���E�;r�"�_h�&��P��cO
��'|,Y���	�◾��ݳ6��l�b-e�G*x��e>u�T� *@տ/N�Ҕ�	��1,��W� �(Ym�>M���E�s���s�:4(Nlrl�H?��3�k㫫EY�PZ;��Of9G-�!��Alj�m�2��,�V�r��a���Ï�O��5�x�mv}�y����+PG�	OP��`l\9��
��%
�ʥ���A�A�1���T8˔g�@)�.:,/����cW��������7oN_��5{yг�Ʌ/�t��R��*ȰG���t��O��ND�@��N[��Q~S���,�<��5*��Y3�U+�9,`�� �6�$1�
(qmN@�L�Pc�Ets���N�;�O��2.� ���σyܖ(C��Oj��'?/��e��s��_ܫ�E9�`C�F'L���H�+���At��	𢁌�N�r8���d�>r�{yp�y�R8��=ڗ~�ɜb�� F��+q�]9�q�.�,��A�I��O<���������/q��p�y��>��f�&��L�h#������qVP��;~y֬ve�K�Ry|h�jn�s>0 9�J����64��1Y.�],���+:y���䍍��ֻ�B���X���#]Q>� ��54=m��0���Lv�+�i1t�\1�b�+a�ి���2kj�+u��pe�J��0x��T��G�s�3��rJ٬
I#�J�l 	G��%�[��>Mx·�9b��_\�b�;��N�H33��H��8�ӟB)ǩmm���!�;m�&�B�c�%]�T�C�HKʛ��#y�?^�=gN�.��[|�	�U����#ܔ)툾A& �2�Q\��8�xx�#0�.Y�֮[��Ϫc�6w�қ���������}�8}�c�ꌼd�B�q�C���:�,��r��
Yp�'�\~�/">�!_d�{�u���,d�����Ѽy�\���$�̰)���_��E�<Y�}ґ��$Q�cL&#^���G c�WpDa��(�=��L&�~(�7����*<Ţ�#R�K�[�R�G=?W�;"EY�%~�7�^������v�~%�f",ep�}f(�P����!��РF�$�T�� z���p�
B�t ���a�L0����?/�u��#�������E+�n��}B(��۶����g�����<�\Q�dج�,���b#|���x�ܹ�~6	���!�Ϣ\\�h���|�~�=�w��/���3��ƺ�(ܜf�I�%�*���
{p��Ǟ�Kb�w��ޕ;�;���;F�0�`L!�A�Hj�pJ�f� �޷��/�ſH/��B��
Fp;:������ߕ���o�]침g��q2x�.l��΃N/w��qX�q�pؘP��H�c�K��k_M�����C&�����'�k������o[O�йh1��d�c:H�B���0{/]r���c9�e���B��gy�_���^|���*�AW�7��>k�^ ���S.�Lě�p|U�.q"�G��T�	���)�1�(�x^��V�tt��V�bد˚�l��W�<���}؍�'�>Of�x�2�:t�K[tj���A�hx��G��=�]�q�qU��<:^�sLU��m�����B�4b  BV�#w���ұ�W|X��z�s����@R�:� Dg��P�B�ܙ����I3 uċ"@MK��R�n���D��7�$�+2󈆆A�N��
�~�s������j�:���AW>�wW��@ӹ���EQ��%jׇ�(O�k�A�|XT�@q��#���rR�
hV:P�:y��Yf�����|����A��A�AU����Ι�����W�TQ���=k�<ၥ�#���.4�xP��X��2�@��ISΣ�l�Qǅ������a" ݦe��#ީ��yn�Ϙ4?��k����xz"���F0�G���R��@Y%�.� �Fjƀ+�)�˗.���Ǧ��ts��`�[��d��ʀ��Ry_��_�z挙n�����z���5kV[B���>�ԃ�:x�"H�[�n�3xko�t��̲^�2a`)\�uc�%��E�EV�J��sX��`��&;v��k����I�V7 :��� �t��/�Q�nV���_Y��vm,�?"F;p���%v 7�wۍ����}?�4���۝��@���yp�Q�M��W�Fα�%Z�)��ql+�l����=<��	�"���s�}�`X�b��l�3�9޽kw��?��t����}�G���l���\��x�gO=����g�NӰ�ne#�$����s׮����˭�%&a�lyԟ�]�r�ˊ�q��vS.��h��y�?��X=�_�q����4ZɈ�ST&~�����,G�~�������Ӯ�޷� �ʦ���؎Y �����2@y�t�{�����p'{p�O>��`����s ��+W���_����"���LVۧL������=s�w"t4x4�*�	�E��d�P��g<��㓿����3j����k_��f�+k3��!��O�:�����ڠw���i��Y���]�	�[4߅�`��ϜN솤��_����t�R�e&EGǧ��w7=�_���p����o~3}���NJ�8`7:+w"�y��X�E�-��������x��Z'_�1q�vyVw9l<D��PQh!1;��N�N�Ή�ɠ�d���lh�t�y2���{ 7�腖���E4N[���E���2�]��H,+!O������T���;l�.���E$5�k �(��� `�<�����)z�A �(�g̘�w4{W�M-���<UB�Q6��j�hB�����<�
�I�۔*�[^�z�W F��S��u�7���A�HyƠ�y�_��```��ɼ)�:��`��R�d��'O��^��2!�t�W傭�m�7 /���(�B9��F��'֤����&�e�iv���c�E]3�Pv�'ι��tY��8�l�phuT햋vl��ˁ&�)�c�9(��m�C���[�E��:���;�"���2�?�!���!� ��},�_���K}�ᇼ�\	�LY� x�����W�y��m�~�S�kT�$Gg"���L c\���@1�b�)K�7���.^�8=��g�T�>q3Π�'=��S�˸�˜�@N93�z����/@��/��^�tx��rD��O�C��G���`B|�e4�6@�[1i���5���/4� ?�c����Lyd,���T�V��xij_�DYG3�=�}dLPc��>��W�{"'y��`uLX���@|����OލOI�Jm2�3�����$l�L?e�%�أ�$�p�}���ӓ���,V?�#�4�>Q�&�u��U@>0A��w�_e�(S���#C�/6�/�����
� �`l|w�x�Ǔ2��Oy�n�
0 �棏>�V�Z�z�J�M�@+��}�?�����μ�|���_���iYǎOG�I'5)c��7���)[ҧ����7u�cu��Y��vݦ�������y$G�b��7Ξ>���F9���5��+�z�1�c�s=��y���
�Ov�f0����"Рy�s����F����=�(g���PzS���k�y��N�B�� -:
��Q���0�E�٥]�`ЬЉP�d��|��'�������{y���`�� [��t��������A�Q��������<� �s��b����Ke Xtt�����{֭��66Mw��✹q��2��*_����	v��>&�ɾϯ����s�������$�\) 2�w��v~�Lt�%,g�7��l�w��9D3�'��#�ot�`�{:S䖰�L��	�5i h��)E�E�,�8r�����6�΃A	#�/v�(q�1~��4q���'}���F{7��N��M�x�I�&	���6�rp`g֡�7��`�C�F;`�'Z*��*�/FsM[���I�G��y��FS��$̛�V�\ɦ��t���t���xGKGѶhch�0bp�#&>���j�Vt��I6Y�u�R�{nf�$�~��1�x�A�E�)w������<�>��t��Ix�i��@)��`l;�B��CV�� J��k��
9�䉽wIw�8��i�&�*#��N'ț�p�oʗ$�U�h��3\��xF��em)��3�GLfh��u>+Ϯ�ŋ�u�:ټEet�ƀƔ.��v�2�&� �6{P�`g�ǋ����	<lw�!G���)x_*���Ï��|�k����C����Q�L&�Y˙����rd��򁷰'߹sg��w��~��J��0��)K�c����ʥ�?c�y�W #|r~(	>ۘfϙm�.rT}D���n�Ь'�`vĤ�I��������j�	���R| [�U��]g<�l��r��-����<2�	�@�ߩ>��1�u�`� N�c|�u�����aH�~���-�1q��!�9ay^�c����r����21OQu��w?�hzl˖�~����/Һއ��籣�!�"����`,�۴i�s�u�֢zW�p���������3�)�L)O�1��@��9&���>.�S���z��>��ר�;ʀ1�r̎r��p6с79��/X� m�����$��j�p����sѓ$�!ȂdÕK�/�$��u%?��EL��L(v���˗��<�ħ��g�{��bz���vm�N��sk�DDR�*~�}������.=���.T �D#��55�>{�i��_~?�ڹK�PZ��0 "@�I�+~ԙa/\�ȕ�P���ʳX����o|ß+�hr�����K��t|~�Ǐ~�#ͤ�*HhĲ`��6�W�S� q!��u�va�@����FА��2`>�����Ɠ��W���L�r�	���2M�����F^�g��T��@�����V(�3_�K�g�'>mA��jw&�Ӝ���A�F9���$���*>�ٲ�^�G��E���[�j���)���&,�@�uv�̩�{�'�� �&t����D�؅:L�yX�����&����jh��Y�8w0VB v�ڕ���eQ�p�@gM`�5/9�>H�b`� ��i�Ny$�l*��b���5�fx�B>)���$O2����Q&�38x3u�k�A{��%@��hc� �3��y'�p�ޙ4P�h	O�S��C�ҍ�h�G$����IϚ5�Ue�Re��ʄ�v����_p��U�y��HB�H>(�i�'8�&��Μ�Y�,Y�ٜ�	���;����	4�w��r�j6���^T*��2��UL�x��[�?�f� ]�r�����
�m�K�A�#��TO����$V�6 ���8�G� ?�Hˈ6���.�7�����:��K�-5�`�YBx��S��v����'nꊉ�"������t�ml~郐G 	��斶~k��K�!�v_|�@m�xᑾ�v@b70#8s��z�k�.�a�s�B�>i̙=�fo�<�l���^T;��Un 3��� �*�F��yN[�E���-p��;�`�����7	Q�v�d J�v�{Q@Cya���K*Y�O��	�W�T����]�L�5x�Ͱqـ*Do�Ф+R"kr�E��X�d�~�+�Um��#�>��h+�K�#�'=D���\�m�<Q�19�2���Wx�hA�#~�i���q�ô�&�C�;\w����-H^�A��Ha�D�|˟>�����Ӯɕ���m?/���^h�(�����ѾS��X�9�ɧ|cΜ9����0 .V�黙��&�P/���0C���(_ʼa�m���;v�o}�[^e�$Q@^y�̞���5ˀgʓ�yƹ�hk�'N�"? �L�G���s�dc�&(6:�W��p]3��C�m۶�W^~Ÿ�D^(K�Ϧ!�Q~P�+���y�,�O��2�]�<��������T��m�w�����1-8r���*\�y�vaα}D�t�4h*Z�~}z������?K<J��9
�kT����ؖ��i��5�.�C����2pN�`�� v��_|ς��C�.�
������F��(ʅ~�������J|�ϳx�:_�c�� �8�ʁ4������),�I�6�k������ߧ��]=C��L��M��-*u�r�+�͔���{9*?��Y���NE4��j��>:�"���4�0G:>r�F�GC�X�rݹ
�1�tvk�{��*���~7?׻��_P�f ˋ��ӄej h9��|YC{A�@�����4��
�۸Q�EQ���/�~w��#�irծz�Fp�5�Ұ���5)m~�a�����<u2�?�_3�@8�ж����z͚4�|���ΥSgN����#o�P���:�hGTt���UN,�ѹa��y��v�Zo�D�K1ҡ�0�h����T�N�~��V�\�]֔4m�,G����f��i7lJ��P���?{Y�픗領���W'9szjje���4s���r?r]@{����'��N��w��/�R�H�~ ��;����Í7���g�6����-��K����FH�\�9�}岕^2\�h��9d �f;ȃ����@2��Y�v�������Ӊ�'mgJܜ'�t�+.�L��"f��t���K�;v��v���y�����=�7-�z#M��
Ђ�����T�7�գhG�g�x|����A��|�qG���sE�@}X��iL7mޔ{�q�M���:b�Gv���}�A��ؕG�0�U=���I�̧PF�_���O~����k� 5a+�D�s�>}�����=�v��c��$]*����r�@�� L�<��_�:"���/��a������L��+���N��H��:��iK�S�[��I�2��/�˴��	�N2q#n�x��m��z�d'�m�����	����)���|���y�?�V���&e����|�2&vJ��9�yŃS\���49�gsO�~�_�S�h��?ʡ����=�ʕ|Q��W�����K��Ą?�=���6y {�Scй��_z�!�ڂ��\'��⏸\.�7��8�O�(q�o;�`�x�p>���V ���{��#��u��n��0�ü��_����O�UkV��'3�lT���}�-��Ť?L��Ю�$�*�ۺʒ�Pʜ>}J����d3k֩ȓ�¹�kN�ۏz�~����'ʁ#�8́�X�E����'�x�S=�����w� ���Y�\�8`��f�k��ʥ����[ʹ��p�۴i���"�+B5�� �4h�Q�3h�a�����S#n����Y6�O��Ȅ��`6y��t��u�80`0�Qa�$oif�G�L�,����y��Pe�vGy'���[�6lXo�9�ĉ�ǳ����[�D�Y�dq���f/�1[G�m0�6�Q.|tv���:!��m�q�\����gn�8�!��}tq�pe�������c�{A��1�"����4�:E'������id~"W�����'R_S{Vs":ʋ��Rg�4�B�Ďn�6oL�4x��99|�P���v��;��Iv�F�6)�s�O��M�i���Q���!9�Dh�F0h�&q3g�el͌x��<���$��@+�׮Y�-��	�Tk��9�p߾,C`y֍��#w��Y��=�v��ɇ�3�be�����,3
:4����e�#��8��~�� e�-��`߹K�䃙���f��g��=�ۼʊ����w��/φ�YC�
 "�rDY���v���0�`r���I|чe�3�Hp��������u�I�2��`Lh��	� ^�_�a�`����8�s�fl ��&�e�o&t���F�8y�W����m%D�%0AC�f�����l�B.�+��"lh�X>ž2�,��L��㆟G[F)/4��nؐ^���s�=��ߴ��/)�4�i����p|%�Dr�	L�n��aP�:��K@�GSa.?�6��/yB��E^#�Y�t뼘3߄�q��r����Nb���E[�/���G�(�5��y*ޅx�F7�,��r�{�H����\*��
O���F����O��;��<�&�?�F�]�K�i�w-<2��6\�G�Ǫ�,�EsE�H�u�B��{ҩ��p�d^����l�E�Ws8~�]>z�U��<�����x/S������}}k��,ß��/��9	�vC�>JMe���+J�� aޡ_��S(�O�1�D>�[&-��[�QE^���&}&m�ܶ�ݴ������%��vԍ�B���-r_َ�[}����6���*��ч�y%����+�LL�(?~���4����KJ<�v�3�7E�(�U�;�C�rDx��	��`.ʸ��
S�O�;�Y�hs�P�^�p�驐I47�OK1@��2i܀=������P��>�천�V	S:&fA�~1K�;W����&uXkװӑ�6|��r����Y����� :��v�v:h@ #=�m��k&b6T��y��t�}��j�|�l:g*�΃�F3��&`�A����*a��u�5�r�!����A����l4Ҩܚo���u_�
���G��N�/���x�}��_apc�����;�����%�?�q���;��J���O�3�Zʍ����w�o�O�K�ϠG����K-�,�9s��36N��(���b���`�,�=u�p��pCjēU�w<l�5�7��fj����3�X���c��mq�ya�i��ft>hc,�+y�K\��3ʰbI�2� �y�r���Gޙ�/Y���^g�9���YlA�m�F��s����]��єY�fz����$���i�ϴV��v�mmmo�=6��,��pt�� P_,_3x�џ8q�ZQ�꨷,��v���O�~Iw�Yީ�`�B�rKm�;<t�G r" �z�&�h�9Bj��.��t�lt�V�z%o�g��&�2� O]0F�Sf�!���	h��c`�A��Z�d���=� N?�Ψo���m&�ڕY�D�(;ʉ<�w���[����4�t� &]C~
��{�� Țb-�y��;u ��� ��6�a��s/|�g��w�FM&f�\4H>p͒�H��ĕt�i��>���"��{�(O�odi��~���O�|�3>�	�=K}B����׌�(3'�T��!pm�.�|Pn �Sc<�_�1��
G���̋~L�8O�U��7�����_�EΉ�1/��Π,&ȿ�d�HX�a���z����k�5~�7 ~��09^�� �"��p�+�+����|�����Zc����nh�4��M���Ɛ���]҇���7�#]x�!�ʖ<�	�#O���k ��	�����3�`K� ~;���+�^�Y����^t�1leb��/��']�L[��q5u�\��f�O�N�ԗ�޽+mݶͦ^�`P�16�	��a�l�5e�l���G 0{E�pAx���� ���H�Q�1f{��>�"�I������O����~��+T�E�F��5���(�x��0EP�=YC�� �V]�9�����.�u5*��ȩDdV�i	A��M �{��В1�f��r�� @�� �}��G�g�{.�Q	�t�>BL�A'F<j߳��sS�*�	}�I�f����^2FX��+V�����2L}I���p�)�eY��������A���uk��r�/׍�O=_G�X�~C��`�� \��'��O���QW��/�ע�s�X8�G��9�/E]=�YxT����G+�~ο���s�w�g��J���w'(aG�C�!ZbyΎJ�<�9��?{� eEC�Wb��a�@gHgK�a��԰�N�<����� B5|����ќ���:`��V$�}W.�fi�:�[ꬰC�;�����C�齅���e��QW%_ȯO:Ф�_�����&�����!c�˦1�˦�K����6� �+�.ED�d9�]�v�خRƜ���ޠ�Oy��H!�'��.Z	:�<�|��~���Pۙ���*��f��7|N5����}�Z�5���}a��mna�jP?u^`�����#΂Bf��q '��19�G��Y�f�C�T�W^�$x�W��h��-���E�S�]⃁�U����f:
���OkS6���%��Ѵ�� 3��ХOD�3 9�M�r@�rD}E�
�s�����uw�.HG�F����Z\Gl�je�=���}����IQf�_�m�
�� X�eW'^7��?���y���K_��O�l��������q����[����t�\��(-�&?�R/�0����i�ǆ��9�����Ƥ�u���/u�5
p�g����fbh!�,WӗP�|	���8C����S<(�0]�e+�W9�i�1�X��SZb�52�����ehd{ ~4w�_���*���a�z���Œ�t�	���3�� RӦk�>�#8Q`Q��TV9�T(	h�L���r%=�S�f�-}.D>ᗰ�/���0�ꤎ�+Y%coqcjE��r9`���P=�e��`D6�ȣ|H�I>�&ݔr�ĽF�Ε&�k0��o���]��{��LQ��-�)CV�Y�f5� �������m6�� ��:�;��8���������L���1(鯸��T����DݲZ���޿��k��7�xS��N;�{O�i��f��(=��l}[׷�V���z�G���7�P���7���=d6&�H�2O�5?�]�. �y��\���5��Sd��.t�,�8���30��]E��@���&a�ʥ0c&3`�q#<1���T �.��GѠ���C`�ɳ�s���Ν%>[%LI�@:y����^�,�M���Q�)��)pOg�ѦǓ4��qa;���`� c�;I~�-fM&h�W�Z�8d��QT��������+ =zD�M-v��.��s�,��'9�fG2G˸���W���<�%N�!=�4n�8:0ۅ�V^\��ˍ	�rJ�ACu'���#<�`����`��S�+Ϙ��w�ӣ#��|f4.vt|���CK�cC f.��.�g�J|�C�X����ov�?Ǥ`��ì�:CY�a��l�2o�m$Gw����]Ф�*;K�N:��Y���:m�Q��njmKSZ��N&`��Ϊ �p��#��Dy�/y� �8(�@/j"w@<3�g���3�x�V1`�6��R/���4٣M�� ��=�GI�� F9��l��8�.m�N�i|
G������e�'20a
Dz�M1�.�KR��93������U�Z����r�)I�ɠ�䕶�DG<��ȑ#	��A���Z�?�2�ޙ1H�7�/��� }�Ϲ����l��p�>��IƩOed`M?�F#��H{��e^mX�h��m���0�6h g��%k�!N�ӕX.f"�D�6��rH�i�,.�2�ɨ�$C�E�0i!�8�)�r�&�' v~�~�q���Λ�~ˣ[�c�?�O�R.D(">�?�?�3PAF�kN�	��rx�d���3*^'�OE۠l1硞�i�`c+'Kj_�"��䪈��R�<�z�K�QQQ&q����mҎ�K�\��6�,�P�
� C��V�=Y?�)e_�'uK�Ѐ���/�F�!��⤼����>��з��A�x�q�:*�"��'��fZ�F�m�"=�.� WeMz8�o ��o���$�S~���\�;�����?����(?�G�)b���#K���m�Mė�?�{�D+�E�ߘyӞ�^�\�}ZH��P�Q�S�G�o0��$_���Y�B!v��A�=~���?H������1n�c��ҥ�VH����z@�@�E��1��?��"���U'�͠���&��8�3���/�����Ȼ�#�9eK]@ѷG9��R�r��O�Ͳ��r��8��"�Ov��=#��>���fL
������G�3K���T�`�L�;E2X0O'LФQ�,A7�3  ���wh��7ˊ ���B�v�/��e�fFf ��;�$`��(C���[@-;2�fڴ.Lt�h����Dy��b� Xy@�0 G{sX3/v�T�@��s8J'kM]�*���В��ƻ\�6�f0�k��0D�u���r���Q����Y���Dy�A��.����A�9�'���#�f��#_���,�t�\�6�r9�Z������<��r��?�H�丏N���i���T��(��`@�@Le@ai��C}R�6c��y��{Ҡ:�6^ͤ�E�6��rT���vLM�g�M3�ؘB�Ј;:5hoU'9�N�"�XNe�-�yst�n��8����%wd1�2�)�0v���v)K䎶�j�*kw�#�@:2:5{%��|�h��;�$ߘ��h"���Mz�7��"��EhN��2'.@<�@>|���v�T����j	�X&6h*�eƧT ����M��E9y�(����|F6u�b*��. !#hQC#�~���nx�|k��sh����~�v�Rl.o���%R�#�����_�70(�wd��� � �eK���c�)����Q͚��ҩ�Q>|B�J�ۆ�훲�G�S�ԍ�E&
�o�ŊKh� ��3�S��Fq���-�;�m���}�#�>����<�+q��Ӌ�z�	,75��	,�軦�Lr9�n�f��@:<��5IQ��A��LHq�E8��<E�Y�a�/�wP�(# ��U芗�����]�ʲa��t�²�	�@ r)��pQ,�ٴ����n�1٤!� "�Ϡ��7��oE?�����I@��%�aI F��ym"&��"���3j��S
O�D�hG8�zC�����W���lPlŉ$h�#9�}9� ��/�9M��N�`�X�~q��+��'/n[�4B������lg�O�d�?o�M9pO>Ʒ�|Ev��q�xI�6��y�Q��w�(���N}0F��S��p�].;xB+�&֦�,H��(9�p�_��<&L}E�2/J� ����SeG~��?ڼ.�({�������6������<�PZ�����]O�� [�_�^� 탼R�ŕ� ��)o�����?�u����B��-�ax�HZV���7ُ�`���sD��cY�B�s�NB�G��4h`p`���������k�dc�f),5��>M�;�zƀ���H��!����k�Va0�`�y��͡�l2��l�˒�yϡ�i?j!�`��i�e�A��e�c�������*q�f�䁎������7�H?��=�C�i�� "~ĉ]�		�{��D�������������`
6�!l�ydG�_ $k����Bt'�ƃ�A��(;�<�O\�\	�O#3�88�>q��c�M� j�f!��3�"��3:b��o���p�
�e�I����`��v�ំ؆/t�� 6��E�b23o�@�Fh>�E�)�9z,]U���i�`R�����9/�A�k��m��O�u��������7o��k⓼1 ����8��͛���5I���R�A��#�tz���<:� ]QG�2�#����%�U:Qd�p��<[���_�+ �t:[�����	��sO7UF�
} ��o ��or��M���8C����c���4�(Q�[��ZLv_Œ��6K��ʄ?�"�!Y��,�c��!��yd��>������q�
�̲ &'O����[H���;hx�'��$�w��������6���=�++V,��Ix��#���E���� �}|���&�#s%�<�7��%�
 "�'��h�z������ʃ2y��J;�:ڝ���6�f�;�������}�݌�t�o������ߋ��	`�7�{�ϧ+�=�M�=���9�|_�9F��i4%56��iRo��7��)���e��-�O2(��. /@��)�{L0Q�b�4�Ie� ^C#�J�)�>Yy��10�c(9���h����P϶�, /J�s?���V��'�������GxD_H��1�+�:���Phj��\�Tq澚+<�8�ꗸ1M�\IwP��ΪW���8x�g��Vv�E�k�reBN������`O��
���q������~��x�>: p	
����/�����]��t�o繬I��Ȼ�b�p��;<I"�G��Ox�Qr�ce�IWǭ�ԏ���W�۾V�����	/��u\�-��}��+8lYv=�S��q�o��y���,�$<����M��e��R���<��d/�2�`:���uا�ɼw&�]��z��0���}��eK; �
�K��̟Ǥq��x�������==>*��H9���=͛'H:���`&UynH��DgLDa�d�y,�2�km� y�*��e:p� ��-�@��}����j: �
��`��W��r@�ȍ���ʅe�;�b�*֎ys�*�j �j5�#�̶����ۆ�%҄�CK�A����0�{����E��q������B����O���]Q�<��F� ���S�V���cӀr����e�"�������-�F��F����Z������h�$�#2����g�y6=���-�,��9�����cL<�χ~0m�t�'>��ti��PG����ڝ��=�Z�Q�iMM5:q�NnT���n횞�/[�Vi���a���!M�؄ՑN���:�Μ;�za d2�w��ME�̙�,���|�6���o�(3��&�'�e&�� .Y�Jy_�n������5PO��đwٰ���ٸa�;k��e��m{����<a�� ��T��9���>�d0!�3w��Ym�㷚tL���F��S._����~���'��=�7b�{]�=��<��gf{�1���L��Zm����g��Б4�k׬K+���aބ������Ra��tU���׸b�C�6���ǹI2�/�.�W�GՏ8x(ф�0�ly�!��TP�$sV�������Կ@4��<�Lt1��"^���N��A1��2(anݑ,�궬��!L&8Ŕ�X��	#9�/f�J��h��쟧�}���f�5���]4�=*�k�/�;#�i����CJ��W��?�c��]̜9/��u(-N�P?�d5�� '�jc���;���ƤB��f���>QFh��zP<ܸ��4�i�D��]�ć��TMf;�u�Y��`2!>	)�8q�8݊Yƪ��wX�y�.o��je�0x�-�B�fQ�Q�C��D8��BL���2�Q?�+
��ԇ�8�L�[n��N� p��ߖ%�wx/�����3~s�xH�:�"���c-qd���/��C� B�$,��<����d>\�"��w\3�#&��]��<���:�?0
i�
n��Ōtg^�� �>�T`7ȱ{\����|v��$�����P�Ox�D�r�I�A�� ��\+'�09�o�y���]�.3�ɪJ	�#,rĽ�XGO9���E��I���"Yr}S��l����&��|�.��Oa��1��~SϾWaJ���jM�\�G���7�b��~�Og�{N��A�4�|(}�_L�ˋ������n���1A����%K��KZ���Y�x���a��y�C��`���+W�ŋ�j@��/�9�J�^-:{�a�qa�	��b�roT�37�6̟�༫~�����E+̬���bV�l!�XcF�3�\�1pL����+M�of�hר,4��d��wm��sպ���3��\*�kv8T<T��t�.i><P��\��N��S�/��.��8b+:b�H�P�a�i���ճJ�[S\lx��N�����x���h�}\����������;,:�xǿKqe?��N�c�t׮]W�'&?���'5���%�66���2�nT��P��	�@��V'�1j�]�*�;��[�5UG���4Sr����b�A�Ǧ��W��]���v ���4���^U���G����Z6����D��䓎Ɲ�D� �aa�Ş�y���Ȫ큶�m�(Vj�AM�`�� y�v9!G�	m������Z�;��M�C���MZ�cYW�OV��8��6tQ����	>��6�~���,�/�u�եN�g�� ؉O^�j�t�xG�H�>-T��-����׀:�h���}��Ɔ #@ܿ��'O�C�{�� $����� Zdn���擭�nUy]Q��9���SZj%����� ��h��2G���Sh�$���k���5���U>�[	��'h�0�b��F��4�W��lC�	x��A(s�&X�4)�H2���t�!�~'�R����"5�#�Y�u_�C��� X��:X,\qo?����t��Y��'Q��^��~�X�,M��%���I��%�˪D��Qn�u��q�
����p8L��c�Ɗ(�G�'�� L��.������_p�C���!�`'�#�?�(��`�=��sO�'���x�G8?GY�N����Ω޳�Y���������~��w��,����Q~�%�'m̓P�����lr�t	�U���~�h�T1�\��w1��_fÎ�N����DY��S�(�y��[<��9���s�t�o�0�*�R����ƯK�0� DY)sꞾ�mO�����S�9e�x�y˦4Lx����W1�*��Ǐ82x&=ʋcʸg����$sz�`�N�6�ˇ	qf�����< �Y�c�������c�jg9��T�3vu��e�B��1�R Y;Zv,Wb*0���NB��3� ]�p�A0v���*�%|�>}�\:{>�� ���s7�����b��C� xd���5͚�f���N�@�1�o4	*BB���`��ТÏ�?y���9>��Oh�0Q�;1l�3��h/�������h�dg�g�8�JV��´a�yY��Y������ HD��\n���<��H4ցd�t~z�U~4x���������q�w�;�W���X���-�h�8�C�x/�Ki`;KX�B?�u8������?��E A7t՗�@����eB�tQ����1T6�U~q���sz\&k���B8~3aY
��Z"���w��Y�p�&I6B�I���R��(�H��]��;O:x��$�+��5�jw6/�{����>eB\?�A�f7'~�1$����������cހu�Z�划m�NRy�	qR�0 ��+�KY�y����=�2V�����Kl�#^�l��3^�S��������W}�3@-�&Dh}�0�<}*=~<��C�˲2NfX�g��|h[�b�)�S#n�k,��[���kj���,�zp��叼�2�7D���?}$�����Q�*�:�;ZBD!�$O��/�}@�1�!�#���AF)� ߴg��ǡ��s�LnД��?�-���RTM����:��q;�o��b�j>T���	S�Ub2t�ԩtJc��_�X���	�Ï�q���.��0�b�C?�����$ؤKX����[�Q��a�7��<��;Gc�`h��͕�c�9�`r�-�0�������3L+�䌲�:���`���u�D�zͲ�R��~H�2 �/Zg�;����p4Z��#plRr�*�I��*�ȱ��;]�fv�4�Dr	�k0bYB��^X�Ӯ
�����t��V����wy,��	�|�z���TM�Q>Po3T�����͘�aC��)6]���;o��+"1�ñ"�<S�!�1�5 U�%m�,�]r)��UX�rE�(W䅴�-[���X�Vj"�
��5�Қ5qzfs^�Z���U�r��֭]�I�^n�=k��0N���p��8�OY�Q-"��	,�UE�w�0c��ޮt�z�A�e��䈖�}��������cR��H��x
�� )����R1�o�"�V-;��<�i��Bă:�I�����H�Ô`�Ҧ��Ҡ=�ܝ��J&N��\�Y{���"����&Mj�f;��|�;>"P�p�B�ٱ�;g:�,P\�3W�xb��<2����㢛����&�������mry)O.[�G��?��r�e��ʪx���g���}�Ȼ��%�x%:p�"���E=�x�4�}W�r��X��.���6�y��g�)xC]?���������/vnK�8چYz[SK���+�Ȟ}����i�du�
�nם�J��X28*7E�Ăe����R��Q�H��;����N�=cm6cX�t�;�{�Y��TtSZ��ˑ��xI�刺����{vY���%�Qu\!o�Wlq�/_��{�����7���t:4��Ź��̓���5#VB0�`e��K��-LD�1\� PᔕfL�๹e������+0�����[�xeȓ���iP���ml�G��>L����?����S�n� e9�,�а
�Yל��CKf���\`OϪ�5�o��4c:�*�왳]�t�+V,�$�c��y�+��n*h�cƠJc�
�����2����o�i�6<_h�n�|�7��'L��D�;߶�U��]����~����� �yb׬���n��e��{xY(�OǢQ�>�6����% �J�eZ�|�R ]V��k_����F�����S�IwF��3g�M|�]�I3�v�9_����Sߍ�4S�o������)�$�I!��;�W9�P�~����Ѧ2��;<��W����#��8~4}���ԥ�nkr�2�Ŋ�������%�S��F6��	2�(�_p\4c����l��?�C��0�Þ<1�s�!|^քg`�X�x��2!{�G�Z�u���)74Ixgۻ���|폱Em� ��Cq�����#+u(��b�������c 2���7+b��
���0��=��e��f
��^��
c8�
%O�3@������w�<�8
��y&]�4�o�H��vK��y��Z+D�{W�G��վ�&�z[2�ǫ ��3� 7p��w%���?|�>�Hk ��Yl���G���1�`������˗/IN�#��#?�ڙ�g��]��Q��|ȇ		a�j�7��a�^�Кo���b��^�қ�I_����0O��.����E�	�Q�MD=�����i<��w�k�QRB��� ���XQg1f�E�b����#}:344����r�<�mݺu���,YRwf�r�N⑱��+�k$/ e^�����!w���ovm�t�
m�N�h���p�`Y�����~�����q�m�_���&�� .�x���^�/.�Q����F_�6:|�l\�� r�wk2�k�+�a���JTD��哆Ļ�+������i�s�"�������_�[~�� �j!E�<0ͥx��k��������; �YN$�ƾ�0���>��D�e:(:�5�צ����@�N9B��� ?��pr�_�rSOL�A5��/�;��1�[��g�0p誃����c�� +>�W٣�@N8x�` ��%g\Z��n{F�	�FSwO��9<z�']���8ȫ�Ѧ� x�c#�� ��$��l�ac�~  +��N��  �2`-
��f�̳���(sʺ6X�n���
�?���SB�<ppf0���X��z��ؼ�ҫw�+�lB=��C�+ g �HG���G�P�����|L���m�������V>�AA���R�Ê�yGV9�!Nc��y��xG�KX�b �LїP��F�X���F��L�K�>k��l�T�����>Ɛ�,���8qmD��M���G�#�h��ȏՎ K�C�)�C�##����>� $i��F��v�Ǿ���ȑ�l�#�.���&|������>M:�vpLO\ps�Η<vX6���Jp2��}P��Ȼ@���}��p~^K{��F �W9O[������	I92 �_����$Mz���9��C�34�Kv��mY`5��+}\�p�#�;��S�4���3�A����Eo&�f�cH_���=aǌ���+�_L�<v�����>�y�c#'��*+en3*%D�B��	���c�����
^�Y)�
:/z�*�u�M��[�E~�{��,����z�o%�yB�lz_��6��I.�A8�!`��/Q��'���Y�i .9�ɡ�'��8{e�.�'OhI�yx7/J��q��3d�{��0���3'����g�I��?�����G�/_҆PZ,[��ǝ.��x���VH`��r�*�5L�p����+g�3�c�����凼ǆ���{ԇƒ�(��L�# /&v_��,׮^�� z}��ǡ��w�T~�����/�3	�����q�|����0)3�����/9�n�>1�x���
}���>�igΥ3jp��P1'@H�g��jZ�j�+��#I4�ޱu�'f�F��a��0w��;�",q��E�����YB�c�����%>3iW�`�tu��O9���"/��3	ŗ�$�!Z �"^������N�����\B*Ȝ�ˠ�rfU�����(����K��_v��5G]p%MG��6�S~�0����.�p�3�G���!���s܎7��a$�`"�x�� T�̿k�r���N�x� <,Ҡ�� tq\ry��@ԭ��//w��2�`��޽���K{��M5$s���dw�"f͙m�e�$����R6����A���>�K-�,�(������~�ka�pE�d;8q�~���;d�I!�H�Q&���n�C�� ���ZJ��1�%<�8|�O9�AƠ�"<�D��|��Iʆ|1x�>��<@m: �H6{�>6ql���	���:�ܹ�Z�����O��I-�Gc�<͓R}�.���r�����I6�h�.@���v��.����P�d*�ʯd�X�Ĕ8z��TV��5���=���2�b�K� �����72��D>�g�,"@�5e�w҇�-�nt埜��s��1xQ>�A���~@��H�w��uk��	h���7i[�}�x�\L6��,р�@ͱch�#� x�8����/1�6�2|��N�� 9k��M<7��Фf
����[�KVLH�h�j*gB�r������"+ ,5��� �h���S�~�Zr�{2�D#.׉~�?�@6H��9������0;���ƨg׵����*�)����e�a��͛pz�_�\ �:�FBY�>y��|�3O�{�׀
�G[��F�x0uu��'˨�2r	S�K�9�r9e��<.�D�"|�m�'OB�ܥE:���!ȱ��oF�x��+�/�!Q�~L�3%�7@���ˤ�m!�dSiD:h����p|�r��Y~9�.;�y_�?e�Ο��W���lyL uQ�C�G'������f��|z�.̃8Q���P������͎#?𼄭
(TP�ޒ a�@�6�f�7[�j�ZRK3gg52?�0���/{f���Y�Ϊ�%���Z��7 ����*��p����|���<�@ivϙ����\�73222"222�H�7�Ty��Y+��6�� ��_p�z�'�v\�Uڮ���	x@����O���e���'�Y�Ȯ�pw�:w�5��m��y#������?�dx��,��L/�x��-��`��?X�>�W�g����#^(�`��p�>F��J#�&�����p{5�+��3��T��Y�eS^r/��5��\���VX�9�u��|7�������c�����D�{P�[�C�B��s���##�^04�[�{�c.�^b�uN}�|ge �.a������r�,k�Q��W�ly|{�(�i��<�^ʭ��<��:���w�}�Z�yֵ��B�Ātyj;�@:�����P������%���M�}����G��c%���o��V��V	Gֈ:��_L	��O����o�{ᅶ�̬OV���QGQ{�ǡ�ߪ2�|�Ow���(l�.��*e��Ȍz1E[>��é��,��Cy�A[��PX?�f�/�^ܿ/�p\x�7�j�Ü�P�?D�x�wV�N��mJ>|�<4!���-��r���~�m�=/EqmT�������T��
`���Z�\1��ޘ/\�BS 䩭�c��KXXt�`�M���B�Q�M�?&��c�oU����S�j�����S��׿�	׍׳Y���<��Ӌ���.Ro�@$�b|҄&�n#����E���k5xg(Y��_��^���,�=�;���/�d:��3B��#`˳��q��W�O.���ƙg�^
��>.sr��	'l.��!�L���]|��c�w!�S��P </�����t?�T��Ґ����c ��pι�f�â���\�a��9��"�A'�2�b�_Y�p����F�f]o�bO	�kK%Ju;�k�����Dq"����k��'��߇�iC
�;}N�$�f9�c?v�œЍ~K��نR<�z�繊	Ms�XC��Vtڀ5_ò�4�|+�_ס��p�8�]�{#�/��9�?�I���O�c�kW}i��׮`Jc��9:�]�2k3�-�={H�xN�dp�'��:f�T��6K��(�qz׺����ٙ�d�j�#D��v}�{�i��qc�����{��6�l�:,3Xf��H=�'C(�^h�Be;�\yŕ�5�f���Hִ���g�V�a�z�v]�w������A������-��, #���{�mw�z��d��{3��w��ߝ~�:��>��%��r1���[�ꨌ%�ܣ8�T��6��ʊ)���M���;�	��*#�.,a�s����V�&�gsy��EyB��3��v��E4��i��<=��!x#��j}F�K!���L]_�FyB��S7��b��|��%v�B㩅��׀o5������&�*z0�Xp*OA�~���"�Χ#XG=���-����vqɀ�y��{U_~���h�RӛQbjDY
���tNS;��k_�㼎�S�G�"�k���K�|6�Es>㌞��Fs��g��=WJڣ�(��g�tT�����Q	0��^��БE�U�C��O�y�hn��1��)أtآ�Ǟ|bz~���X������jui\	�|��צ��	��Ӗ������)�������:�]i^x�t���'�;f,P�X:���J6�ҜB�_���H�2�G���?`�`QX�X<�-<s#��XR1WV�)��űvrA��}����oϴ~KU�ղFP�|Ls�ڳ�c�֓�-w.��n�c	�(�|��l�V���[�Q<_�A>�ԙ�g���I���ʓ0,�j�26�1��+�m-(1�τM�X�w�
�~u`��>p�}�>�
R�����1�}V*�8W՞�SJ��!��"t&}�p��F[x��:v�����1��q]Z����}n��W�6}�#�~W��������[o���k��^�ޛo���A��)�ȣ�5Zx���qU�����¿�`�hN���i�S2bw	|�>
/z���\��k�k%��)�/�n�����Z�~(�:m޲���E��n,PJQx_��_R�21��6���@i,:|�h'uy�|@�M��;n�3[��{�"d>{@kO�Z| ���������Cw�~����L��O�,�0J��(���z�)�������~��>�J����?��?�n���гv�A��e��ޅ#4Q�Hra��O�w�w
&x�|�Qz�	^��ROI�/� ���K:yk4��+�����t�G�z�%}C_������<[ﬥg�৔n�|�t�I'�:>�g������ v]`U�W@,�����]�qh�c���9��i�Χ'{���6�����K��<8P�(��R��󼝼*��ˇ�s�x�mx=�1_�3H!{6&�`�e�m��������5���sꩧ�G�m=K�p�J����H|G~��o�G�v�����;���y��de��{��{u}�t�y�L�|�#��
7�t�tKu*����G��w�]��8����o}��'��d6̩Jc�6�}LP��uL�H끀\J��O�����pT��˫�:zL���6�{�Q��U�B�j�����*�p����#*��#�?�����nV�"�0�zF�EJ۹���]Y���]N��w˛H��x'D�O�z��Sv+�[�+�g���jzV�7�Wa�av�= ��&q%4���|�͚a�}o��:�ǲ�,�O����O+���� �����b�,fe�:�m�>��OE��M]��>?��C�Dh���"�{��|�
ئMǅa�ya��J�{�`	�*�*�H���Q�=v�(&p��(!|��=~�|��l[
me��j1��@-:� ���ƍv�����C0Rӥ�j���YDr��?����?�Pv}��R���/��B��W_��_�cM�ZY��;�=�ƳA���T�Դ>�ן�Fy�U��7�r�Ʉŏ�c���(ԔKn#Q|�����Z����\)�OV�{���GQ0����.4��<��b�%4/���L�.���ܳl)+~�U펁�E��L=��F���׫���ʬv��
c@��j ^�P��攫!���V��!V~n¸��}����m���kW�]18ֵW_�AG��ʟৌ��kS��:��#_aY��sm#�z@�z8F0.�A�_��xg>$�{�]��~$;�x�)\pU'*e��������V)����J��&,�o�B�u�E+'�oò�Q�N�X���U�u
^ʮA�����B٭������fg�VrM�*X�3P@l綱��I5 V�R
�!O��n�[Qk��|���}ɧp\2ƌ��c��G?�~��eV<����l�|R��O�Yt��j��?�gӷ���(K�73��_����뮋{����鳟����{��������������w��oO�s���ow��?�������
������z�u5���Mb���77�^�C�8�G{���ݠ�����i�|�����tY�i��%���Ue��.e�x*�'�}&�-w�
���)V��w�0��c�Q���Nh��Z�^t�t���O'Q} �C�i��ȗZ_��Qv��-*dp�_*߂Y��fv�g���v�[�7������Nɿ��~�\V�oX4�>�T�P�{x!z����^�_����Z�6�`��7��G��ս��}udI��#�3+1�h��*�Z�!��
+9�+�����Rv�=+���4��6?ncfm�I��T����=}⚏���{C)�����4�������?�+����/����o|�4�W*ȡ��^:h���I�ܬ���JS����8�@i�������N~"�(ht7aXv�T�5@�j{k����~#�@�!I�d�Eh�1�\�߂Q��"�^�aT4�a�����/�0+W}�0V'a��W�}U�E,�܆�;"e"��P��Q �2t�f�#7��9��=g�a���a�[p8���u.��|\;�K��|UrX���L@�o�H�� ��t D�n]�1���9[�Y�w�5��8�T�M	��c�f-4�yŕW�R�5�I�A�#��`�V�zתdL��YL�X,>��X��QU�#ԣ�L[�_�v�GV��F��V����4�USG���[�}ι�i��>mټ%���0���\؆�GL�z�J��@kƑ����f���|QvY�1.��#�<�e��ݻ{a@3�C�Ymѯ�� ��(�i"�u�_��բ�J��3[m\��wz6�Xu�7+k���BR�l	
�,�yvW�rrFs�p! M���g�!�4��W~��{�� �i ����/3O�;(,
�������(����3���ߕ��:Ú4��ݣdp���A\�B�E�R�
/��bچU��j��5�z�T,@��I%p����W�^}
Z��A?�>vf:���4uR��_jڧ���w�ͺ�ԱAK0��k8�F���~v��W���P���
v��u�"5B�Ղ�h��׬įF�4��E;>��r)�'o��I[�fN�:�(�ʬ�ʦ��4c�]�{��)�
<�,sp�S���.'o�
mE�(�,�x�IU&ECj�B�t�M�9� ��H?���v��GM>!�E�����Q��L��?��(idt����^�Wi�wġ����>��_��t�O6}�ߜ~����������c;�?���{f()j�w����R�.����?������ǒ��1JH�e�B��
%�3a����:�.\���~��<>��OM��{��W��:�=x�(��{<��OPn�N�p�/`�M7�T�M?���/����8ɹO�3�g�n?��O�c8vnM�	Sn�ݺ�wa?���s)�Qv+
�^XUa��:�ɟ�o�C>˹����{��{,����'�Ns+�u��h��
�O�0\���n(p�>�z���iHp�a��^c����OodT��^�o��_Ԓ����D+AA�J��KV�����?���_��;(�u�Y�������,���*��7�:�v����E�}�]z����8����e�V�ܪr��z�@	[���S*	J�ٖ3F��Ҭ߈!�q����O����("+�1�F��rPN�'�:��2+G`f:��L[@�m�c:E�0�b"V��0a6��'��e�B�2������o��~���3-�q򵃇�[�0<9ą��$:�v�/R�ӧ�,⢸�P0t����bЬ�Q"���;@�B��Z��������ұ"��!�([^���]E���j@�WG�f���� ���#RJb�*��'V���=(F��k�~���](�}�_�Iv���C���I��
�����N��J`f�h�(��ш�3�Km���O�)7]�N����8V�A����z�۔̝��Q�K��*��'�z�6N>e��#hEjY`2��of{�z�`Z�����B���
�r�a^\px�^��<��iH��i7V�О�������\��e[�����	}�Ik;V�"�
})�-_��k~0i]3�~��������O�v(7�Ւ�:D���m��f����)+�{<e�LRu�9�s^����[aT�u�p�R��,�/�x ���VW<��cŲ0�%^;�'��
����+e���� ��,*��򁧩��F�pѯ����lկ�ћ��Y�U	տÒ�Q�M��~�+_m7��J 	|�[�?���P(_Ϡ�JP�Q�Y�(�RnM��r�xd��]��cF�MA��A}X����SJ{��j�6Zݗ�k �]���zk���zΗ���S-��9���
+}$H���/��>��3}_��_p�3K�Wy��ӏ�����/�3=�t����R��_li����?/��o���eQ�Ϯ�����x��/����_����t��w�������vh��p���������lo����i�n��cd|==v�q}������{������hܖ�zYLw������(������)H�u�0��/�[I�^�u����Q�E�®g������{�������$�ed��@��Ϗ|�������ʫ�̞���N[ͭ:~G��]���#�kx|�@[x�������w�G}8;1����5 ����W\;�	@G�!<�2�����:V,4TE� ��:���j�[O7��q�.2�+3�6�/�Kou�����ĔM�q��`�~W��Uȯ���<ߜ���S1�n=O�#�?������oO��v{�_��U�T�\�f��cc�9�3���{���}~�ݏ��e�G7�|�t�?�|a�����O��?����od[@7LJ��B#�P� !���@5dŷ���CZ�ù��_�����)���-"���iW�\nF���u6�DTJ�W@)��<Ӂ����B�ELF����Q�2�BT�bQJ44�S�<��|��뮛}��X|+����'���b�XMY#6�Ҭ�\���z�2^-E-���>�i{��},Vd+*�bK(�e���+QD�ۇ;|/��s{ʺ;���v��U��Q�T��M��5 ���C��QLv��h���F��u��L�7���8����GH�*)����?�6r"���W��*HF��茣؟/͍�7u��Ɣ��|�^Z8���?��?�Уm�p��v]�1p�U�X����
�C��z=���J�Z9ke32MFb���v��v�q��Pe�Nε��JJ����6����F�K�bx�m�	�v����2���Ү�:�v}�w������{�k	Iu�=V�Q����dmQ��Q�Io�z��
�IHr��רO�epZm��T^���t{H����Gp����	L��f��Ȁ�~j�_n��s��=3�H���3X���mڲ˕ofu�=�U�R���͹�>�J9�p�:��:V��ޫm��\��h�睆�{Ҭ�~���Xvge������l7�P�mh���:�K �r��l�tb,n���Dթb[w+�R]���(��ēOd�߂�(�����4}�K�6��	x���H	�+�-�}~��N��7�H��3.Ǌ�����W��u�q���@yū��={�O7�t����w�]�0H�+<��K}㘢�?��?ȶc��vF���;z����Pv��[|����ݗ���`f����)�>�5�\�:hg���4��A���v��G�Z婢�����C�"�o}���f;-+���XuL^�s!�܀�o6��,�+I�����OOw����_���/r�b�o��_�җ��0ˡ���o6n��<��.�ϔ�O��_�zF��ڜ+����[o���޵_��e���|@����Q@����y��e���n8�3����c�0���s}EfҮ�?��S�=�2�~Qv7�[��ރ
�d�l�f�)��G��^�����
7�w�V�=b�w��OK�����nLi��9�1"f6lO8,��o���'>��]�,P������Z�F�5��^�Q5��^w�Xm�hj0{WV��hcI�g.����C�H��حC���������j�b2U�r��#t���(V�� �Z��?�B,�Ĺ|c	���睟�l�	���V]ʮN"��T��?�(�C+�	hDz����?�/���8�S�txBNg�C&��!@k@�p��A�Y��Л�;ۛ}U���:_o�G�7N(�=ub��|�35��B5��{D ���UYi���-���*gK��\W��GS�<�P���~���C�Rv+Y���A��B�fKRtoy5��w�of��zU�]�m��ӄ�d��gb,�#�j 7��� �E�y����$���E.�a,���f(Ŏr^@Կs�Cq���,�VL��i���yYN��~# �Q����N�=�4� ��������	|�u����뷅Tb�"�	)!t�T��f�Ա7CsE�K�a1�\���޽{�f5XQ�$�����Q�հl�e�ŭ���b�a���k,��sDں�2XR3C��&��J��U>�����jSl�k��3!�r���f�}L�A�ꍆ���ZuZm���~a�V���:���7��X*���aoi��̬��6d��b��I�ʊ��O%t;��aZ��~������piEb�a۱(��k.�mp��������n<~S"�u7�K�}eWP��W�g�na'eW��.B���B��l�jxk`*<���X?�6(���l��&j{*�B�8�ĵXA{Rv�g�q�=�x�R����H��v#���LXg�������.O}]P�638����W���,z23��F��)��.���c�\{*�µ����b�Qg�r<Ee��(%�������(���
�A��ھ׃7�D��?����O���ק��9;��,�ڵ����[��vy��Ƿ�`T�t)��qY��?���?�a���|�ㅳ�ǅ��(7���G��z���<���<���`�K0sU���"ߓޱ�C_�͏~��io�׫�����Oր���Rш>�]c���(���oۚ�ۤ��s����5����g�%�*�[��[�M��6���g��Ys����SPj�r]�R�|�� .}���J0��T�_}+�����5��_������ ѝj�~�O�d٥s�~)�\��������J�!
3Щ��>���R<J�(�����f�P v�{5��;j��ܳϔ��|�<����'>�����=Z���������R�����u���k��D�y����R���<U#v�?�ЃU惓�������*����n�SO=�b�cA�c9ոj���q��=����ٚ��Ξ~�7���t��	'P4LwQ<��b�v#��H8��α�*C �@�;��Y�-⻧n�
A���aN���N���~���~�
V�JRN��T�(H���^Gp�O�u}1}�T/�Ci����Jg�?f���7���*�a(��I[���PТ��y�k<u�_:v����-��a�\W��!��n�ZE鵠A��F��G)�P��OU��maH�{yL�g�ֺ��-骲�C�,�F_>:!�y�X��	L`�B���H�D٘q:.��/\��������V����д�h���g+S��I*�� ����"l�^so]�3�eף?9�]
ԧ���j����OO}�`"\���A�j��,e��!�U�$��*��h�0	#\�R;���d}�.���PD
��v��O3y�"�?�.���@��x�n�`ޖp)nIP�c�!�gxI�9I�8�[��P�MO�qtO��`�?BW�x4�Z���e�`��E]<��<XC��c��������+����W,�Z�Юv��y�D�3��B���j����`&ʻB^�c�U��������dPPJ������"�u�՘�|	�7#�~��N?��Ϧ{�'�bp�'	h
ݒ7�|S5����� km-
g���_�å��z��5�7}���Bw��'���ȇ'V�C�l?%�oK�=����σ��������X}~X����W�x�4i�B�m0p�j�%h�pKY%?�HR��C<|�>>e�g��o�pCѵ��6�p�7���p��Y@��/ŵ�?�r �n~��
�K� l��-��|�����C��'�mG�b�V}�_�ܼOߒ]�e}�=8�_��\P���Ey�Y8�ѯ�&�t�r\�����F��;��TG�&��_,��ś|��~��=�����CjQpōAP�����sϗ���t�G3m�`�ZΛ�GkW�g����z�W�g��K����C ʮ�&b\:d��X��'�>Y��];wLO?�dQ_d��d��=E ��ȾTʧwi5�2)�;)��zꉊO&�'�|<
���駦g��g+��|��:�˥}��ơ(��a�[�6�΢���:�۳/;(l/�2z�X��R�bfܫA[$�
�UWS�w�uW��D��\sMF�W^ye[���S�)�Axq,�U�^�/����U%CY�U�F3|�}o�b2x��1��Q9�k|�{���F$��g��G��0����m���{�|=7:�}�fK8A�͚iU>�CB���j@/��� ���D�*��y�w�4�w���~�}�jX(����jw������=������v�4]���TW� �a@u��Bg���X��6�H��s�����`,XX��}�-�u�{�>���1v�F�A�~Avb+�Fݮ�qs����[7������SJ|>�ZG��Ut�h�/M���daU�_B�UgueeQw��m��G]j�x���^p�<���2�>+�d��O�Mׄ�YL�1�g�V0���}����ձ�/a׬z�E�2�=t$�
�el(��/����(-�C흅���}���uƓ���b&=��r;?��_���>�������EE�   ��IDAT�L^B8�[eGQ����.Z���e2L>��"�
C���X�ଞ���ڎus䡬�q,�k�_
�QG���:�� �}��5-P:r�O�����������,x��>��c���;w��Ж]
HgŨ����������]\g|6�4���H1Z��Ԗ~vy1{�ӳa�*�V�m��#�fo�r��>3�����5�x�?2���ק>���/
'>���K9��s�{¢�+�؍�(Rt���&�op�RǴc)R�@���A�9���1u@�����'g���v���c1 �����{G[)_�����pb�E���/�_����w�o�q�hփ~a&���XmgW��wԑ�C�2�M�+C�xGz��E'�i+���uNw��_-�{�t��{o�P��=E?��U���5h�U����Rv��oU}_�!�!\m���Ѵ�tdիd���1��4������}�'�����I'm~oeQ���R�|��>���&�ew.�Q�E4�b�5Z��)����t)�*�������J!���!ӹo�J�wιE$/gk�� 0@Ͽ}�:��(�>���s�)̻+��H ӹ2샸����K �}֙E<GU��蠐� 1Ofn����(����Z��t�bV�>L%��I1mi #��_�����q��'�Lʦ�#�W�~��=�g�W��:�TfG�Y锘jw�}�.����t:���:q��O_������S沥T�F��5�A,��sQ���ę����,�)a6}G��3ϴ��x�[o�(�Ub�ɫ��G�\�g��`nWX���y������=
fw���cD:*\`,k#jφQ[�0�B~�86<]F�R�|�?��������PdM��P9�o�-h�(5@*x�b$Y���X�:�6Y�]�O+,�+�!t����k�U)̶���{�'<&�ʣ����k��Z��%��W�{�1���W|&m��R�#��nL�P�����������p���L�գzu~+4�gn���cڤ�l���i`0�6�q�WF9���p���Tx%�+�]}�j����R�� l�Άw��}�y����х���<a��vXM	��-x��	�Lp�Y�vT���o��e�ȼ�r�Qŗ�>;��Rl�Ѱ���P����}�u)�.��7[���O/b��<��(ϊp^P��?էlkG���r�> ��� �W��\����}u빼F�s^'��>_G�vo<�����4q�3�Ͳho�auƿMw����{�/ک�B���x�	����k�������;�Y���7�e�����OL�>�x,������B��F��Jy�oD�݊.���t��~3ޥԡ��wE��d^uՕ�׿��(�۪]��f�1��nLsF��7��n���`�Q���{e v�u{�^P��ʏ�E�/:����z�@��s�̨�煒�ϒ���i�T@V/ ��ƂAlj�D'~
.��5%g��ebQ~=F���QwGw��;��<\�6y�����@�~��s����X
*���Շ�^ܿ7}@=(�>�mq�j��Rl_�?�߼��w[��]��3;wT|�t0�ľ�s��8�7���Yh�|jC�f����3RfeW����ޚ�{~�����d�0��>����y8d\��/�۲{����Z�i��C	��.&uZ)tUNÖ��'a�E\�J�SO>�
���rR���m�N޺��T�c�#Jqy�:ű�h�[�pˉ'eA�#=Xi�*�?:J����غ.�;����q�aX�[]"�Nl)���O����-
��e1���>?W��g�|�Q�x����g>�:"L'��t���bPE�:,\鬬Ǧ�X�.����\���2Ji:}	e�����:L��+B3�_���Fۤm0�e8�9�vG>��(4��7}�F�L�a��������X:,
Nҗ(��K��=���sϧS#��W�)�a�o\�e����pk�R�`�P�#@S�;�gv���",�;�_�Vm%\�$M3I���u��c��W�Ց�S������"�{ZVԶQ�y�B�q?�^�~n7L���G��p����d孜E�k����X��:v}G=]��S�ͽ��]�0��X��y��|{��eTn+�/g�)B�@���O��������/#���Ƈ$��3�-�h� p�K�W����в���{�0�+UW�/���z=w��H6B'�."z�w�����ڰrk(b	�[�V2SW4�m!M�9�9��w�O�@�[�F~3�~��%C�G�M�*����7}�u�U)�G�|,��8��՟��}߾�K)�p3�b��T-�����6;��UZʦc���Y����x��=d���z�
iB+�%T?��K9Tg�̆�|��v���PJ���b��|����p5�o�f��N�,��f? �	y��R^[�M��p�����(��O|"nL��!�6n,�����/u�d�A�����Kl����/|�?�#Pt�����qI۱.���m��p�%x��m�\q�ٸ\������й�y����K_�bE�^rIɢ���f�H�zU>o|k�7岞�ͱ]$ڳE��m���N�r���S��ـ5�Q���+�:���e��#�-z%��K�����s�Qҏ�>�~�t�)ۣ�OY�Qbч�$�*c�Ë��Qr+X20����`6n��>Z>���1�U�ЙM�ч��^v���0�l����G����bW�̐��c���:����!Q�������X������97ҝ�';��~ᛦM5���e4�:���Y��[���k��a�:��Q7v�z6�0�����$���n��w��$���*����Vv�z:���kJe(����k��4_�V� DL߶*ڳ��R�6N\p^�m	q��V��j�A�=;SŬn�t��gĴϞ�>�Q�E'o=i:q�qs<��u������-��@Hݺ�Bri�s�p{x���Bl�Ū@���h�'B�[��s΍U����:����rU焃���ꐦ?X+,HS��:�~�0
�\e��YF@5j��F�x"�c��E(Xt��%HR��`�_���⋦�_��(�HYud�6��K��B'k����d����a�sA�J�(3u��(RHN(��p�LC55�F�����H�����G��C���N/��<_����^�Յ�|5�����y��Ä���b�|oq��|;��(�E��D�P	�t�]̍e�מ���puF���ׇ��J:��'1F�~p���{�v��<��:�ׂsJ9�V�u�·������|�N����F��>�*^;�^K�6��y�a\���~e!I?���A���V���L����}��4[h�1uX����_�F{�!I+��
g+m)�Sf�����Y{�t,W����#���el]zǔ;�K��b�11�ԓ:�>U�ު�`E|�ϩ��}>]�o�6E7<��\��l���69�x���5���)�tqA1���#���p����{���k�͎:Cʟ�Fey�o2+
�M�/�]����o�j{Y�����b�<�0 �@��}�1�ɒ��G�TUU?8�����.����l��a�;��!����ib�/_}��������%��t�܇CeSRo�~��i�6�qO��v}�Q,��f�<%��Y%V���rm���[����j˺DG�Pª-�ϓ�l�찼^}�-�'��m�K��9*2��M��Wh4X�g,zV��Q�w@V-�X�ǭ���ҋ�(�q���8��+Ӿ=/L/<�\)�d=�����p��Q��i_�W��E�˔���,����re���x¦i[�\�K�bI��t��O�>YWd��СWS��ޙg�MJ�8�肝2_5J��,QW�w/�����CO7�|st�Xv�隯X8�]���Gmq�����=(mn��S�o�k�L�}pV�QL'Ǿg��u���t�5]t��������}���������Q^*p�"�Vⷦ��5�PyKu�E,�wk�O)%���N��9����j�3N�^��)y���3��O>>�P��C���q)��m�(g[Ja>��q���Η#�AP��C�*�i!�(ЗN����a�V'��3�6���v5}���ctm�:v^E���U��P 4�-B+�����.���O||���>:����)_=(�`k��NY!��[�I�����0�]4|Gp�\�^vi������g�57��t�a�	!��8��0��\�H�|mڑf�����)�I���h��6h$��	������_),���Y�S��������Z��Q��0�E��E�kI/ҴP!x�i�?-��FYo�}R�������N���η��g�����9,l%���JKcܮ��$��Pɥ�&p�Q�+|��S�O̺���7�/�mD�y0�2t���q�H���hZ9��_+�Ϊ��X�X�(��^���#]�d6J|��oت�v��^\�ޛy{�ll_�K���c&&����0p(�U�\��+$���Jd�0�D�GJ��<�s�}�^vY>�}�i���v��WMg�sNf2Y���c�NP�:SL��43P���g��V�sJ���ڔ"ҋ���a���r��G�1h�4�(G!���e	�ۆU��ܹ#���e�9ōjd����|�z<z�`2�&_��\�
�7J�ǽ�i�7�+]��>W���u]�B�9��k��i�����
,��^�V�|�_}�:_ah�9�,]�P�x�/�4]4���&3��jv��J�@I�]��\MՃ�i|x��V�g�K�dl��9�SegQ�~����k��27�vq�>u��!�>UM�4��ghǚ"<�U^��4�������=��B��IX ��n �fԌ��-��7
o]pl~��������{�-��Ľoz�����7"x��b6?�w��B1�#�07U�:��XBMc���j�"�C�J1�;�t��@�S�'y�ǧ�~(&v���nt�O%f�g��ȅ��X�n�S�(���Kn��u!���Y2|�Y�e��wM�zNX��}�Q;D<��'XZ����o1��Ҩ��0!W�Po�a�QŸ,���\��"�K���y�#��>�-v[n�)���0��etݑ��������ק���35�	$ֳ�1�Eh%u�i6<�O��(��@�C��?rH�
�5�_Š&O ���ݯ��|k��1��w\#���xHl��x��
��ûU|���?0�Jf�#N���R(B��#��6�/k_�%N�KQc�E�n�y
��ֵ���5s�b&w�Q�)0�sȘ]Ŕ�h��C�_7�s%ь�Ƣ�򍵝歷�:�q��=��>E�mV��HCB�_Z�HC&Թ���z�UW�E*�]�Xi�u�����+E�%-꯹-��������Lt�4.��KScۖJ;"<�X�*R?U�j��Q47^bi�����k+�e��.ʙq;_&�g���lغmk#��vjf��E~�F�;0��.;�D�S�2�[��Pʵ���{ֵ`����`�0y���$#Y��j#��V�죏<4���Ow�q���}�e�|���yq�����`;DV~�H�c�^Z9�sJ�8ZsyNqd�f`���<��ч�v<�D|u-�oW�g��л)�^�EQ]���}	��*��Kg^F9Sv\��E���v}�//�����ӽ���t�O<}��ߙn�����{�5[���R�uQL��j���K�a�b}��n�_��aǴc��8:��<F�诹���%�^��~Eh��	: �T���K�g�>��mA�)N�>7�-��t�	���[�ⶆ)^zɥ1�?Q�j�M!#��أ�'��'Sg�ԹE;��R�#f+��/�``�(l��%Y�f���aJ���i(oF��"�bί�j����`�{ҙ�ɶ:������[o������㓭��ר�N��Yg���.�Q�|����\PF��A�,������_�|,�3��x)�|�(�|�v�y!ʕmd�=���vhb�5�W�.���h̰G����	�rv�������!>Q>�c]�P3|��Ϋ��yeQ�"}�I�>�{�j��=�������ú��-�����*��Zi^x��~g0�S�G�>��w������y+:�'���������U�e�w�Y����y�:E�5�����Mwx��ޓ�0��+k-��IV�s3����ޒ������^���K�ӄ���.��e{$��x��|�y��V��ǜ?���P,�4�	x����*��/�,��s�7���6y���rcT��gzVTf,�3o(��e%�k�m�ݖEY6�'���_�A��U>�P�'������."a��8p����/��U��Y���;Y9�j�ŵc�+��K�r��X]�au:e���M�Սܣ��!�.������X�~������N|��� ��	�?pC�x��¨ߨ+�%���ʛw��ݶ:���F�,���cV�ϩ<<�Ϡ$���|� ��h�d)ur�2��šО�M��|�Э�(&A��n��_��:W:E�5��g�Q�������Ed��=E�G�-#��l���W�T�꼪sh��*u�/ǆ�`�p�!�jzo��;�gք+�g�(x�~���.� ����7�t��E�E/��g�Lv.�6�������l͌���X���|��ӓ���S��:}��O�m�Rm諲0�>�8*�ZUhƶ�OW����{�1���Wyh��c�1���˲}�5S�m����ٍa��8��z�:��|��i���j���(f�C���ou5�F�ݸqS!������s����SKɺ`:������b|/M���"�#�`vLvL�XV���O���:g���H�fƷ���\��ig���KJ�>���2�ʹ��^u �������2�>�9�'\�n�d�lK�������4v�@����Q�sv����M��Y`&Ǚ�:	����8���_���)N�,ʿ�����/D�fY�	���&��L�Խ]��abf����2H���齠��
�m�QZ��Y�}%�-�}��Z�p�Ǒ9\�;N�9��;��G�`v=�ּ�=Ũ7a�J�	��sG�F�����	.F0@kp��Q���߸����-���a���=�M!a�A�w�GZ�U�Z�,۪q����k�wl��d�K�s�s��]fϚ؆̮#'����ȉY=�m��	�z�g�|��.[]�U���p�MG}䃞�G}޹�F!�{�A��#��,t��B�� Cy��DS�zz>R��!?�Av�9�s�����흩/�����E�z����|�h���v3?�è�ڰ�?+�z9�B u=��<'D����&S4:�5��}�3<�r������s>5^�X���l|a	p>���XuM[�^�N囯�y����-��\��}�!G��e+%S�xJ�K9�����)s]�[��g��3�q���`�eo���,�������vM��zk��	$�?��ON��vZ�ʰ��b>I/]v9(zϭ<�@�����I�p؟E���k�L
?���N�l�Ԡ�A
��Σ���� �?��릉��g���{��J#/0˃����Rv��~=��ǻ��*�m{^;t0;��ق1
oø��,�Q|�2�Ɣl�P6���+3���\�\/"EW��y�US��?�B�U���J��F	�a��~>�_�F�Qp�U/��N�Pv�T=#�x��sp�;n�.Zz����"�����V��@[O�6m)�k_�3Θ�)<�M��,<i޺��mM��q>_�+^������N,�v��E�ʫzn�~Z��w�ig�􁮓�N�R�Smt����O?��������h���TDp�!*V��E�ȤR�&�<�W�����SmQiѝt��\e��Qv����aD�x�-�-��Q �n����RҌ����5}�[ߚ>��W:̳��9�|�H6��2B�;���7��~x��?��g��6��r�-��!�U�,�M!7�UyAU!���CW^1�U
�U}����������(r���*�6+�a!�
�D̔T#��L�-��4�Ǫ�{~q��ӟ�4+1�V��q�2�w�}�qK5S�2��g0�Y��X��b� {�Rn���,�1�s���M?����[��{�|�L���=�?��/L�Ԁ���)�BLu�W㡙XN�/�����\�#�����|�����ŀ�Q;��[��|��?����H �RF��`T�$H��\��;ު��wG�.Jh��V�y�/*Q0���_+���޾�vL��f�i+�,0MK�Y5�Y]gPRD��3��mP����9�#
V���z�h}m>�0�3p-���0
��u��.B�� ���o+0�{ב�Z�����W�.�i�*_�J?���]�ma�mφ��a�v��<�b�>{�վ�e��$�m�'�{�nࡃ����l����>��/��O�a{&�~t��h`J��h��j[
IQԂ!�������uok	��/�T����+_�.���V�J����f��2����M'�Py����%V֪[����@�W?�Q�R��{��W�Ի�t�UE <�ph������d�Q�)*���+;T-Bs�KzT�,�dG����*Ɠ'�?dW���~���n��|do���2T~�+��&�q��� F���<�h�<�l�qp0p�BW8/�����s�,��G!�ud�j�s��e���F�pD���Xn������ɥ��?ʿ�8���/Bo�Ի�������o��� ����������/S����rТ#��� 9��ݖKw���_�#O��>�}2uΫ�d�q��;�g�R��H�i�ѕ� _m�=���Kg�k�Q�l5���}=;&Yd}���C ��۲Yf�~)��~�զ��_� ��9fc�}I�&����\"G��/8K��9�~���a�6+��*e���瞟v=�+x�j`�rN�A�E�[��+h�\�+�_��� �y��q��,m�9�.���w܁����~k:�������(�mo}��1��Q[ 4��J�^ŉ �� M�W;Pt�"�J9T�1�Jc�B=ڱsg�>�g��>���L�O�^�uC��dYAA��*ЮM��앃oM7�r����տ�n����gu3��=��ǿ�[��-�%]0}��W����"R�x}��]yՕ�e�\�Ɠn0F�(�
�4�&��� j!]����W?ʍk�#��{�O?�`,�O?�3	�`�F~�V�C��C�B���I����5�`RG,�!��X�%�,��w;͂Y%��;Ą�%�Sﬦ�c��Q%Bm,�c�ʂ�bp�wn)G'��Y�)L&��W_����
�	�pǵ!�.���Ƃ�����E�2A�P�#�->�uN�哂���U9�0{�����#��>1��J3�3#��鮯W�C�ؔ��V~I����{�M�@��m%tl�f��י��eD�x%��;jS���8��j�ʱ�MAr�f u\ѱU��"��n86��/~��o��oO_�җ���W\Y�����#D9��y� �-�}m�r�F�%�U���.����_�b����O&�ܪKQ��D�p�ArҖ�b�48��$ݰ��Et�mk"|�R�3ϊr	�6$Y#�(����L���˧O� ��g>;}�s�����s�=w�]���#,Y��~� �y���z¥�)��A�ŕ�h��2�AW=?���>�aKW+�Y_�њ�OY�����Ě9��˔���������`�����>=]Xm�҅�)_��*~����;��*��Z�D�UG�s��e:}�W�7:����+<M��#����-�!_�yE}�Uj��9�E�u��Q�0�ݻ/A;��.9'������¥]Gl�8���7�j
�}�ߟ=f�7�h���y�)�Ei1�%:���.�:�6��'~l��S�f�ШA/��zo���e�+����O����U~���'o?e:�3���@��]Y��ۻ�jV7`�.;2�9\�C�Z��	�'ڟ��0{��b<�0Pе� \��Q��ޗƌɦ�}pEn�s���R�������V�nYkz���&��p}|�G�Q�瞯�,�{���u�^ғ ϵw��[�R��:ח,F��*}��΃�E<:
.#�#y���Uv�ꊅ7��՟r�'c��68P�� �%/)�ţO����[2Π��H+��nb�����Eݏ���뇪�7��^�s<���[�����k@����ߪ�2.x�,ӑu�.U�xN�ǶO�O=��a[[z�u]E#]��ϛou�6�r��3�����k0�L]nZ��ځ�H�n�e��sF���Vvw��T��T�+K [q��7���Af#�~��s��~W�*�}�at��=U�+� =7�r_�џi��t�E�>���{���<c��y�s��m%HJ�n=��A�3���&�U8�8f��@1�y;X@��8+mu��A����vL{v��%�M�"������P�	�#�L�^Ζ�T�0�?�ձ���P�02
%EG$���L�٦���v�o�p.b�c�����B���ݙ����yT�u$8�:�mM�F�ey��^eI��t������4�+A���VS:|��`�}羷}N	��@qm�"L�";������H��f�&P�ul�U�+��R�XZ٩��G>�2�:�촍�:�F�h��,�ձG]��^	#�P��~��9$`���ǖ��X J�gB�r��S<�k�+?�(E���l�5"\�A�j���k�z��ʥ�r��������Vx:'���VJ=���Q~x���ޟ+e��4!�ep�K�K:��%��mQ6�|�^
y�uh�����i>��`u(�,���Y��r��ѿ���K=���OQg�@s�{�t���Ά�ݴ>ayr\�ΫggUn�k��}���VV����_�����TyS�zj���'B�9~�V���i僻�+�n�sT���w �)�Ux�ĕvF>��y(.Ɗ�Bc���\\k�e�g�s�f)x��;ʮ5d|�[eX���Ǧ�������Ν����Z�6,
�����U�\$����a�'�>�.E�4�m��:���;35.��O�ӥ �Q�Z��a����Z�����~���W^yE)�̧��*�?�lUVm'����p�v��c,�s�n沈+�@n�����I;p*���-�v�J�9�����K�.�^�aQ,4,~�y��y1+�V��3�=ٰ��v*�6�����`��,+k\�qG��RH���Zh��y�X�����QK�#��y�J�W>��y�/%��H{H_x�_�C
��F?�)�f	 X*��{�o��cf}�]"��;��F�)�����`9�����/:���UA��q�^ۖ�q��:�q�}��}w��b�j؄&�K��3E�2H/9n�28�O�iE�N5E����T�h�(��剸��K�w��	p�������b~%e�߹��0>���~�WT�,L@�B���U�������A�J�O!�PTy쫆�SȷZ�j<S��8�-P6� �+F	�d�>餭ө��E����G���������F�.������H�1#c<���E�t-�gE�-�G�g�����#b���@��Vi�)�\����掙���K�.�N`��̳:���&��B<:N�0m)�Jo������Mp�P�c5�E���"������Cף�N;��� ƔY?�f�э�N�y�q}�'��g��Ĳ��,!>�B�1�j��X�	�)%�����8�o(o��6C�����_L�r��*�s}��NgŪ�mb�/�`�í��G5�g��wWq-���ʕ'+,��=7	á��a��N	��]
E���>f'�O��7��R��wǊŏM���� ڵ���S5X�#�mV]]�=��ٲ����7�)租�Z�5�.�N�ޕ~e��]M
�d�i<s�X��ɥ��z�S���)Ł��-� �̖GP�����,�W�F���`�̟�kJ���ײ�1 � �A�iL¯�U����(p�W�RWB��XL�l%m
C�P&e�rڀ����jnQ�tO��v�w�r�Ђ��n�ZQ9�뼻�	u��G8�pK��?�� �G�����n�Ϋc]�?����C�x���~��ꓔ��o��Dy�|IVu��?`�N��!��tB]
��q_l��;st~Qy�T�v�����?�n���,��-%�8�c�?H+}����.n%7��»�q~�E_9'���λ ��J��W�P����YX
N�m+�uaԩ0p<"8�/~�ޥ��������㑶-�ݧ�/���������hȊʢ(du�Tv�-�}�ٙ��|ڬ�Yg��ה߬O]�zan��{�:Y	��B[��9���Tt/�n)�qm�� �#�jЂ��\2�9&V~AQ���>��Jk�K%ew���&@���f�@V���Wx�p�NU��[/�~�xݳ�>�)�"n��"ֳ�_���s��'��Q��N{ku|��t�(�U���x��wB�4���7W��Q1��M�^i{qZ_�u���˯L����[��_x�p�F�����V�ݪ;͈��@��;��
|�|2�`��,�����4g�sk����o�Eؐ�y˶,,�`��y�t�<��w�tj��N)�����荹�Ċ��oD�9�Ҧ�O�4g�P�\#;�׷��N��G!���L�er�ҋ4Xx�B׎�<Lc�����*y;��0��y	�x�h�;o�Ru��	�(�E䄉{�M�~����ڐ'}�v�I:_VJWg$��n��q�AlM0jǤ:t���D�{�~ł�Cٵ$�2�e�:uê�7�ҋ�Lt��-�=K�Ez��ʵQ�l)f]Hg�΁E� ',X0+�zL�S��p��jk��	þ��{2Ԗ�М�kb`�6E�G�2��R㳘���)�y�P�`���|G�ȗ�aq �o+�	��A�!���զ�Gb��~Ţ�\���l�g1��_f�D�#�՗R�)���f�W���Q�պX4�!�h�=�ʪs f`T������/�40P�)�z��A�x�i��>)�]5�c�=��J�2�5��2�;�Ҡ}t@y=�x���|�} 8�ϥS��!%��ܣ�<?ax��h�vYXx�ۆ�9:_tܾ�䢏�G�74X<��n�)Z�?u�lq��Ш�����uUl��e�Eu����nB;�w<��m^�:�"�v�G�=�v��*�꫍ǠP8���_���2�h%ܓ�Ս>�s��1���p���$�A�Ȕ
6k�?����@Vz�8�������:LX��"MS��~t�:��Y����=V<�;��v����p��������%���	S�h�U��:�K��^�{ "�����r˴��~X���
�퇞� �|�B�Vp%�W�>`�sy:Pg�ח���m�ˋ5��iH��cJ��Sp�;�x�>�*�cb�c����s\�0&s�����^��� Yo�\���K�.X�a}�C�S6N��YV�{������Ҡe�D�S�P��G��*gӉ�U7��k��Ǜ�Ҿj+�*S=�հ��(��;�C�����Ri��-�ד����`��}v��v�T{&ֹ�&���c�؟�}�^��:���� �	u�ֻ��۵���
_�*#}�a�����-/����G(��N���	ݩ#�gpJw�z�7��S�?�B0�����n�N�9� ��N#)lt,@{ޣ�F�< 9����"V�4�)�h�oT<�:㖓���{�tn)��^p�t��5R���K�?]|��ӥ���}����+��.��t��.�����3ϙN�Rc�Rp��Y�K8qԆ�쎙�:��.�E�����j��%b�J�"��'\k�;V��8�w?���U_��s:�:��r���W:���^�fclp(B�c�����,}��w��\�?i�K�R����(�*��ɓ�q[�	3Df�7ƪn����?���x�˜Ϛ �A+W�˱���ѱ�嵸L��fz1L?���T����YD����u',��i-0�~�E�g���ր�E���C�L���&8i(��C8p�1sʚ��.�������i�ذ��T�ߞb�p�s�����
�K��"���?�aM��\�� ��c�ό�Zޔl��m�R�_[1)�K+��?���e-#�k~G�R��z&4=�a���%��Kf[}
��O95�v�q�_����Mǟ_�SN�Ĭ�7�	�UQ��U�f����V��}�}�)[K��6����|����m��QJ( �����J���b]�(J�(�@C{���q�eE����+�c�tt	���?*i�o���L�M��W4��vfr���P�l�Ŧ0	f���OqO)��'�y�R< ?�u*S�ڪ��e?��o�,�d��05j6k�cm��s����QUw��K��ĵ�NW^}u�f��Z��:Qu~���jopG>}�K��	�K��#��\8]�+b=f)�1	[$�0�k���|f���+#(�q���xD���V��͊j�?H����(��w�ܑ���[�p#/C����V-��,oq,ԥd�}K11;�ēO�*^�o��oN�Y�ݸ��wvo�����/O��;�����Oe�zK���N^_I�#x+I�J��3Vv�����|�P�?O�S���l�_bZ8�Z�.ZV�K*e�"iǏ�Fgf� ���¥~;1Cv������ly/!�ۑg�d���^u3(a��Ӫ����9��?g�>T�����l���!U^�_�RC��ShC�`xi�	��G1����i��Y��Z�%�c�e�}azތ\)�\^|���^��V�n������Q�yT��5��܁}�Tv��.�W�z�_ݗ=����ILn�V9�������}�}Ǡ1�Zf���"�\�B�
��0�.��H��Z�hĎs�s�X{<��z��)���rQྰ�M��'m�6o=e�z���)��5�Ƈ�l�p+��^x�t�yNg�{A�?o�v���'n��<fc�q1���2���]Jo1ʊ�%a3�D��!����Ѥ��=͂���zF�'u�j<ʲ���0�L{����B��h�>�p?��]��sT�2z^��c���"p*?�S1�\
�j��9W���5B-"���V���$�E�2��U@l:.��zuz�;Măi��e�&�M�I^�=�6���a&�ٛI�;#���s��4��D�\|e��R:)���G��(8F^r��(0utM����O��;h����G���֭,vO�Խ`� G�����Ӷ������p��5p���;�Ԯ����{+
�{}�奢��V���:�≛{���X��ā{y����9�H�b��U�+x��������ӦEO�TEe�$3�W�4��Pm����%�Lh��i����q�nҰ�k<�'m�u�q�F�M��GO���i�_�M`�5)7}�x��=S�|ca�2�Mq`ay��P>8P��b��/�S;ryA���wյ
J�2��Gp/h����V��[�k��p�O.4�'i�Γ��[V�s.P�M?�z��X�W�D�l>i����?8}�K_�~-?Pɪ�N�\�Y�s=S�Vp�O�k���S�|�E��;]6��,0Rt��s�ٱ
�/!��HfY���'��~���U����ɷyR�Q8���nXzVf�hݭ��2xϚӬ�ٙ橧��޿���R��0�*K�,։e������/L�=�l\��y��̼P�z����{�����n̔5Z���~u�������R��L1+S��������m������w�w�^|	o�i4�|�y�;��":p�z�%��#��q���w����P��J^�r,:�v�q��I�q'(��Z���Y<E��O*-��=
��+��Vn�X)�:� �������>�m�,.�Նޡ�J�:��]7�·�^��g�y~��|��x)�.�gU͆J+�:��Be4�,������ܶV#K��-�Z2<��o�W}*�m���8�j+��h�U�L����������Q��,�{��Y�Dt���^:���&V;��î]��L���x��t$
��-ȇ>�`T�錦��w!�8�ֆe�g"D0��5
Ica��ъ�������U�f][�Ƃz|u�F�!�"�z��Lbe47����0�ľ��yr�?�CHFք4�%[B��w0��JSpVCگa��ū:���"3��,��s�(�r;�s�W�qZGw�o
%�pԳ�'�e�T7�N(#жZvH�V�0�IT�t:�$V�'���`�:vۮ��w�݇���O�|�N�N���( ��9S��4:̣�`":5<Px	S��O�λ+Q K+����k GI���K&	��{���3���PB�S�*��3�	���zp�]�jX��	+n���eQ߶���ݹ��YPc_O�ٹP�\翾��RH��h��_f;���;�̳3����v�ՆP#�(k������>�>�넏7��v�]�A�]��<)B�Q���_e��#8�ր�%Ħ�����2[�Q2�/}x����BqcQ�������|��΢i=?�^���>�k'���v��sШ�'A���ni���s|+�������%��6X��n���OKQ +��=~=��I��g���(;�g�)�6em�o|��9%Wz�%mV%T%Q�d@p�ֽz�4Xw��P|��dk`�Y |`��臒i�1[���¸�s}H�����4n2�� @��z�H~�b����q�H�p>��q.�#>��}.
��!��[�����������/��?���l[v�O:]���$��Z����/Eנ]�)�,f,g��Z�I2�60�ŭg,��t,�S��+���6w3,fa������Z�X����\nH��˻��X���2RN�ƣ�<V�~(
i�v(e��^.�1�z/J�6��O���h��~m��Ӽ�U�
F�|����]�&Sћ�ff�����iJ�:�>��i�JK�
����8��C�L����^x[�3{,s�3��ʤ-���6vT'���^��Q/2E�,�޶u[f-V��f~�������)�q=X��;�i4Wpi�i-X�ư���������F�=�\2����l�d��SOO���gU��Y���7Z��S��	���au(V�:�XC/b��R������"3کH��Q�l�)Ld�QyYydW�m�ҍJ^;d��3��;��*R��:�Z�V�TD�i��?_Y粵��;Dw�epo���l�"����W��+#�R4-V�Ļ����t�|�[!w�����G�2G�7�m�<|�)AB��/S>�3�M���R�d7���y���CBa��0���sgͽ�]j�^<[�V��=h���v\��	��9KK�E�AQ1[�QXԵNz�7����E|�K>����(,�l�%:e�X�X]6�]�����s"). Q<)�l_�C;`FY#��Z�0�����O�+�mÔmq��Y
7Dxa��h�!��B̽��y�+��Cү��J�~``�U��ψ��r��2���A�O��bP�:xO�oZp?�<�H��y�'B���ֽ}��SU��x�1|�p�H��% ��B��+zx�kS��.��|���,i����Q>�F����;A��ST�ƊsH*���*�@��c��K/���!^��em:���=��S���1�=�a5x����3���!O0������}>�V,����F��՝��1�U�+8�ט������@�`���W����� ��H�u���$�Y�uO���Q��^����ڬG9���Q_���Ҙ]�յ"̦���S�<
\�E�@S�7���\��&�Y�b����2�㘭�䵟�V|�r����}o��曲{��y��኎���r_0(�h���CW\�A
���xz�hǖo��7D�-�(���<��mɃ�X��]��7�����Y˂�9��ц|�#2�
��UG�\>�f��Buo:�1a౯�E'�4}�P�x�_����Jٍ�^=��|�Q[��9�����6�x�{h+�����l=V:�bv,���Eg{�j�����Ա�i�ç�?���6@h��2�k���~��}x���������`?_���e�=���>��H)�f�Nɶa�N��fW�c��Ӫ�N�ίAJ֜d�|�����_���
�z�z�8�M]r�x衇ʮ ~|!'�!:n�!�n[������n^Ĺ�e��Gy4# �1��km�
�Q��a��^]ۑ5�����qd-�H�t�i���U���RDT�ӀD�f&�[h���O�����U�iZ�NՄ_#[��8gW�wt��*j����b4:jJew��S���F촃@Ս�Ca	�	�S��Q')�̮+�tV��,��x*��]�u�|ɳ�t�Vx�)�3S�qw(&�֡��H���C2��X�7�	��.���?�����t��қR~���q5�8?챢�=u{��ե$xg������hב��o���P0�=����]8�a1p` i1���2T0uD�<4�D�蓔+�oد����%�-4e���d��/�7���� ��i�V�;���p4�䴏}N`P�Y�<��bIɗw3��qg0�o�J��ľ�/�p�x��|s�}��d@�����&�|��~�R*���~
.k�s�X���F{����*�|�%O���m��3�*~+�}��F��L�M(�ڄ!֪­��l�ۃ��)G�SP�W`^Y���_��>�m�oh|m��7xM��w���}0�g�,A��v�'?9}�c���v��>N٢�P����e�_<`b���(��M� �)i��;�
vW�B��`��>\����v���kB��ﷂC��JO��S�8f !�l
>r.���Uf� ێړR��Ж��'>�X;2�4��Y�����5�~�hA�s�Bч���C��+����k�����[��}���?�E������}��Ņ�Z�o�>��qشF��6G�L)
H���4G�uz�S��k�<�d}__4�	���QQ��Lr�/3����Xg-j���e�-��ɲ�4�D�����E�[�֞����|��Ymi@��b�(� �<:�c�+ؖʮ/�ni\_�Zߐ�q>�zTw��?i������s_�����U��#ݢe[=�z��Y�b� 풣������}�-��V��Ғf�=����_u���P��.�F��(<�A�s;ǲ�Nٵ�����w���dW��x��Fä"|Swc�.��������ӡb�Q�{�|�N����{vZ������Q_:HIJ#�������q�����2�.[U~����*ܵK��|ۙP��!<)­���eL��"�AC���;�y��3�u��u�!�D�-�&$��'1W2\={ �Zx$/��q�v=��w�,��H�h`�0���uh�^?��w>�
ڪ�f��� �S��Y�L�U�F��2/����1i��[����2�`��{�]��W��%�i	Z0�S�u���Sm�z(�`ӶYh�Svb�(�a�����(�F��mF�E=+�%秃!T�i�:|��{������Eѡd�FY#�>�|����e���Z�'��&����}����a}�#�N�t�_V^0t�wtb���2�@�|�L�)>bбw�O^��xW_�彿L�_(��/����Q8�F����b@0���7�1��',Ka�|9��oe����sLZ��-`��z-�zz�Ȫ�޾h ;_JR��[x���O_�3U`<��V�z�Vi�e(��}�y�A�o7�b�Y�������_��4ͣ�[�wp�R�`�_���r�g��>�R�W��N}����J����S��Ӂ�ͬ�3ʢ�j�7T�_�ȕ��gиz+�(��4����ߨ�C��7;jK� �-��\j2}�J��j|����YI��9��Ϻ'������=F����E�v���χ�R�����/���wN�-e�Q ��3�q٨��#\Zl	�]_aCK7�x���� �0`��5W	�m3���]���>�x����;�XH7��ڼi>���h���ި��#�[����˾�V�:{�_��z�v�r�,Ǻ��Hb��� �t���<��@�(���{���(g�2��L-W��+���x�2�R��6׽Vt��|����?lֳ��{R/X,����R�]�g�7����-O�I�t:J.����̽���AY�]��X�
2?"'��|eq����p)5��9�ٳoi�=4�3���)��e�e��wUv�J�C�Ȑ�P��2}%�#�a�F=_��f�I��KC;�s'�s�JV/�ui7 L[|��������G�l5�A~�8� ��r�"q�(ҩ�|����Q0e6
m��#x�����Z1<�#P�E(�	ZN�Iw�eDx:B���r�:;����B��٠�u���y���3����L����c �>�KRpQ�;�ܛ���Vt	�@T4��[����4��0zkx��D��<*=X�m��"@11��R#U_��Z��X�������y3+s���"��Ϣ��p��/ѽ��q�K�T�6wn��vGF�h���N۾�`�YG8�����id��f:��BtoLc���-���߅k���]>U{C^Z岦
P*v�x��E4;���B6��>&�6��UV�z�m�-�iS1�m[O�>��d�֡���W��Է���V�=�3��o���TN\��Wl#�%�w�e����*0Y��-0�sT�+E��d@�kG��� <ȼ��ʝ�Oų�EgE��) ������B�_���|��lW���� m�t���A�A,&%\�
���۳�@��������ལNʅIy��lQa�����c �i�8+hW�����>�غ��$��/��H�������_i�T̫��j�����<��(��g|�����w}��j�K.���b�t��C����N��ւP���=�Ѱy�b��`ao�IR��n�~��50-b���wzf�*�բ��CՋ<���l>�}�G�����0�ڠ�E�X���g�ǀ��r��|�'��rf�����U��U>���W<E�O��ӟ�����~,reg��xp�������_���r�1K���K���~zo����|F�U�ځ�U���c���|ʹT�kX3��<�|@C�[N��gʀ;�'��}���~�e�v3��/-h��c�����J+�g��ʧ�Pd�yZ����X��X+�E%���1/h�ԕ$y�Е��$tR}ՠI�����[�I�����2^�����TT��s�>u�B�������ك�����?��Bѕ�zW>���#C(�`�*�^��,i�����}��u�N�3���w߁��ǟ�#�����ރ���|��	�� ��Eq��H������⧑�G}�F�e���9Jm!B�ir*Fѝ���~��yǊ\X������>Y�>��K��,�����qE��B&kq�
��q��_i��^U܂S�_��벫<�h_D ��۝E� 1D�ǃ�<�!Y�0�L�W��)+���w�Hq͋��~��J�y3JAm���x'���61�<sg_�I8J�w�읺�"�'�z����������Bԩ�Bh�h!x~�3o��^���k�(<�|5���0_�^�1✆򑁉X�F���O씙�~�cQl(֔��W�۱.j�5,/
.k��PϢXU�w��^3�9���L����`z}��ɧ��i�;_�+����9M�.�W�6�1SPV�����K��1��0��2ȣ���|lnOI�tR�FX��w��Z��N-��e�}_�}
���;��������S���P	��]?�������\��S<�����6�2��t�&��&� ����:���S��w*�fI��~BIb9��
����-��\U�b���l��������Ơ߆K3RíC��Q?u�¦�`t�4�v��Σ����Tu2x��a\��J��������L[pV<�Q��2���|��Rȶ�S�p��v{̕�����eH�gB�i��U|
�Cq��a� x5���ٕ�_����.�-���_)b.kݫ��~[^�*����>�7�L[��RЫ*�$��Yx
�`��u���J�]
K�T]��~�e�>�����W8`��+�k�����/� �	��A>U��n=�7��
is8e8!S��9bɎԣq+O�]'_�)CT����+�}1��y:Ml��+�^��m��Yў�,P���"�(�{ou7��G�+��j@���l|�;G�?��=@���C)���U�u�Xљ:�+f���ao۸��,�*�X���}��b]���J�9�[)iF��ӛ]����pM	���^ J�]�&�� ��i:����dD��I��o�3�D����
��97+b�C$��>�����J�_�z{x��΁<��A��E�ƴ!	���=-�|v-P��Rhc��(��)|7d��&�����N��&�"v��À!���=���B!��e�>�a/bU>VT�=���bb�҄:&F �û���r��ˡ��g�W�ht.q5,��"]���n�0`��/R&��Q��o�B�����YH	:�����0��f���Q��T�����;��M�j�%]��{���'��b�������`�d�꞊}�8��UǼ��l��yE����X�����7��ϻ���z9���,m�hϨ^���c��������(�_"�q�8l�F����bw���?o:�P�H�>h��H?���.�+- V�U\��q��?n)S���y�����mDY�_�!��Ä�pt�}:C-%zX�(�-�i{)8�0n�.���N�;�-ˮv���X@FW��73e:�i}@�hWZ4��\|�E)��O1�C}������_�}wp�M�z0�Z�u�}�D��P2���b�����{��/���'E��H�	+m��� y��܇7e�QXO�Ҩ+�f����׊�ϷgDtL��N�������z��2��y˴}$�6U��n����'k]y���ڵb�v|��3N�Z)u~��ID��j�c�U;��b�g>�r+�5p	hb�����`%
P��{v�?�A��
YUf��`o�{}�ƠY���f�)���\t�7|�s�ѯ�����foŕ����8(���y�_����_;/�����kd0�ys���rʩ�o���q���g������><堙��-�q��6,�`5D06\m��jG���Y���չ�s�UV�*�ٳj�G�ӯ�@Î}/�����xʨ^b�T/F���K>���[�����c��xU�#���fx+-�5���$��Ti���͹��P�>��!��(��DhE��z��q=bߧ��?���^D����<}�`7����AJ=�Ģ��6ʤ#]�@�m��&e�2;֐��.�Go)�uw��Y�G�-���;<�ˠ�g�{3r���[o_|%y��W#,ڤ���1>eg��[�z���+�
+|rT��Wf媼N�~��x���*rę��>�4=R��Y��p�o�aI`u����*�%��y���7���iJ��{��b	��)��8�W�!�z�b��k����9֙"�_t���Bdsc��릇��:7b*�(��;#.x�a0 @Lٳ�f��<�Gt��c�9ʏ��P��R�Dh��G^C�:�5L è3[�qXhQ�2̫�{�8�\h�j�t��jnC{��Lg�k���^��Gyԁ���QGy��Z�G�)[[c�]��86#?\@\9X��B>�m�&�5m5�����RZ	5J�턆p?\�t�5�N���6D��??��!Kj�Hv� (���C����c���n��I[6��8��s\��o��)�����W�i��GW<���Kah�p�}���^�W�61x��-��g�yF>�q�q��%�	0l�rB)ŧM�_xAx��f �j"�����G�����p��:��u�����]=����w��pi�bN"-:�S	�10
��}c��N7�tC��R�g
w/�R���]�*=���	�����B�u��c��k�]V)���
�����v���*D]�ãc���z(�~`��|!���ADv�9��0x��b����%����ց�ry�y�L���ݳ�Ȍ�6���j`y�G��>��OGA�o�{���e*Y�/ͮx��{S�vw�܀|�P4�\O+�"�Ǯgve�L;��i�`lkb�m�Ѣ��d�98v�.u�k�#Cל��h^��6?&�!�N;��w�~����|o��w�?�s�/��������\Nd�|������,\���{ԑ�Q��~�!���(�	��ƣU���⟩��im�e�1ǝwU�t9�v�x�x��Q���/ŗ\����+���~ޑ��w��e�n���Y!���v�b	f�U����GuL|��mT�'|�l#z'��շ,��O���?��|@�#T�4�`u�_[Aw����14I�_��"���(z*���lｉx(]��Sm��&��0���/�r��T#�v�s�y��K����JOc�n���w�%R�����yE�N6"ă�-��^�@�Uɂ�hq��� �l%��O�)�L�产8ҁ�􀙡���K�FW�L�&��(��7S�ɵ�W�6a�0�˱z�Ϙ6�F�~Ϲ���v
,S5Z�EG�T�b����AK#������vk���kBcG�ڱ:� ֎��k�HR�1(9TK�	'�Pfh�:��"ւҙ���2嘢Tցb
c`�-
̢��G
�>F1{��9�#�8#��~v���i<�Q��٧q5��9]<�C=/�2�5��{�#fJ o�����)�ﳩ>�@�e����4��	�|�1H��������^1V6S�,�-�w�w�	�zT}A�`����ܰv���=3Su*����Bs��\���o�l寏M���[���� u��3��F�}���6�)..A�i�YHuy-��C��}�#?<���t,������Y��);��δ�|L=�/:�`��KS]뿔����J''u[S`��r����1�R:�>�ptFx�>��쯛>W�E�U���G�G�d�6�nF�u/�D� � %��;��޼d����i��bb��&�s\�lAc��}���B���f{�����̷�SR~�����Y�)o���w�]�����3k�O�|�󁹡���mL#���qUn-�Y�`��v��.A������O��~��N?�������Rx�Mڦ����FF�����/"O�����2�S2g��34fv�_��쳠���H��H2=n��ǂ��n&����������sf3�Kľ�f�y��CA|}���1�0�8UG��a���OXu@Oq�(���9���2�B܊�K/��˺[��G��#�t�@��̚U٣��k�F_�?�T��t��� �l*���>��Å0nU�t�ea:a�86p��4�� �RO����f -� ���\(����3�)��X��а�B$BZ�!�F�_W~��yi�.m�Cb#����t#0�a*���:��"\_�I	N������r���G���Qؒ�BR�+�`������6_F���F=]#X���N��b�
n"��X?s���,�Y%Vo`���4�^tJ��p�cZδ��	N�
߇�W������/�s~}Lt5+��0���X�&��S�q_y啋Q#�9V�L���ɻ�S���v��PP|�`0��u��0�[ӷX�	~�,^�Xu���	}x�su1�mM0`6M?Tt�S�2t��. Q��O��XX`*��[F��R��x��І��-�x�����s��+:a��Ä��zkӹ��տ��O5��L��#�R<�����oX��K!2��WU}{V�pA^�#�P��pc8��&+�3`��W�_w,�}{W�� &m���~|�QS���郝�h���Om�)�����_سoz�J��Q�"Д�m�*}�E�����	�.��b�j
p4�n��2
]N�5�화ƅ�����3�/�h:���۶V���i�zM������0���<J�W;�qc��2 ��e˶(�������e�9Q�4`���:�����1����+��+&�o��.�4��G�Rj �k��[=���4f���/�xڶ��S~�p�� �7��ͪEw�Ls\�c��O��~FѲ�����oJ0C	Ń���.��}���~EY�?)�m�V�c�aa弭�㼣|)b,��p���?���y6^G��i^�R��^�4[��>,���%�W�x��|�}�v�_7�r˭��΂�'�)�ã���{�@�a���"��u��KE��a����-��ѡ��Xw�sO%�9��s���:�������o;�L�Fl�K���)�Y`V��y�P����;`pO;XK�8b�Oi��|�G8�w���c׮W�?�}vޠ('u���+��c�wn���j38��K����r�i�C*h�1��}���/����3��������[Ͼ��Zٖ�n\�M���~��|���C��d��V��%��\��R���9��Ҋ�	���3����(��u���c�*J�r�l|��Vb�<���l��eaF:��r���V-��Y�?���<���}���q��1q�~��G��~�o���N8��KOHcbR�f��N�N�� h[{ᦕ]� �!D�nu&i��j?ç�~z�뮻2�s�}��(�誋M��n;9#v�i������1e�w,�z��
�!a����0A�a5��m�K~�����"C�\g��a��1�H$�`���]�fF:~F��@au��3Q��?v�E��\,��(��uR��GH��є��Rr%i뾈�o�̅`tp���<K�c��+�����{��W��[���5���k���h��i�2��?+��
�]��F�
�d��^�gÈ~ew��k��oKw���-4&�g+�)��|l����Oc�&���`�;w�J�c��?($;�fE{����dtas����N��Zt�+R�A�r�}.}^�;VR�}�0��ۢp�	�S@��}m��2��F��*<�Y�te�����K���e{~Rl�)�h['�k���m�p�qV�*�c,�T��#l�����5��Zq��3���f��H��g��&��xx�4~�<��\�+�}���颋/��)e���M���^p���7�����)Z����.8?{!��u�tJ�kk6�W��:��m��7�9��A�B{Q.�(D^�a�$/P(�,���a�҈d�bs��}|�{�YgQ��
_L��l�0�Cڿp��Aɽ��K�p�����h�%S��������!%��E;w�-賉%���_�2i������7�E�d�����z��'be4��L�R�~���_~O=�d]?Sti?챭�r���h�4�ϥ]�x��~�:�?��hm��Q��>%	������C�j�4˲9RL�e�\1d�g~���u�]՟�)]gOx��+%;+_oVh�6�Q���L@�P�bX�v\,�������r����#�O��ܺ�&�����Rv��¶����<��Ќl�ۛUϰ����]?�?T�}�[]��R`K/�Z�<���YG�����1���[r�U�h���ܧ[%��6�p�Ϥ��p�`9��[�{�U�s|���|8�x�_�Π�A����.����C(\�,��{�{o=���v��b&F! :#�*0��O�Q(E�,�� 8X�n�uC���ҫ�-�����{�T��rM=P� �B�譖ǜ(eF��!�FH�O|3�1R,	��4p)���P
:%X#��7��iR�y��Ǧg���×Յ�&(��(:���uRx���q%���J3:B��.��{��K�n+��K����O7�)|�x`ᨗ���"-O1#Ҋ����ր�L�;���i�C���<5���C�F�?�����R�HX�0��W	<�O������!)�=p91N��U����3r��dw�b�/��G�v��9hB;�^��|{9|v\�.��hME#�k����+���b��aM�2W0P<)ã�Q���`�wڪ�z�K��B`D��_�eA�]1L+vp��e�n���<���~^J�6��+�-�n��Xh���}p�څp�:���:Xy��H�.���%~��oP*.���~��.����|D�W�_�S8.���d0_W���a=p�J#�7hA��ܫ#��S�'?��/S�-$��` �]�O��d�kH�@�hѹZ�%
�Vq 86�g�v��]y�~C�ky]S��gZ��EF������*_�r���{ι���a�h�_8,�sL�s�F�؂.�Q��'�4�Q��2��|5.�.Z�ݓ�����k��m7���fC(*�ő/4q��$���,�hMOxd򪐺9���eʨ���,rǠ.l�l]̚�o�{|h�x^;,��	/ ��1�6�����_�'x�\��3|�����}��On�;7�ze� ���ވ�욢L���ٜ���Sz���K%pX��ҳ��
t�9�8�~2�1x|�X����$�%�mH�x�<c��P�nI[��fڀ΀��b= +J#?�+�s��g��vh�0F�z�|�l?士i_6k�����.4��Wh3��>?hʽ:��}��/kڨ۬ڥ΃���ۢ��T=R����Y士Q����D��2�ԢM��<��pxI��o����J��t/�K��&s���W�|fP�>?t�ޥ���ݓ�x�=�����r����nW����z��9a�O�qnؘQo��*��k� BE�z8X��A�ҍ�^u��������M[����~�_>~�B��^Ai�ض�T�*'�)�uTf�ǻ�G`�|���M��<��c��1�!���?�/1F�)�b��
:PU�4zF5c��u�C[�
[E�oԈ��m+�|���\v0j�0d�1�C�[��f�w��vT|���|��"Җ�}!6���S��!��Q�k�W��}a�����7���6�i���)L�a�V"�OiY����Bh��Ճ 4�o��x��*�a�-o� �_,]����R�O�6���3QZ7x�˧kPc���E
PQ%>D3lS�2��>��霊ހoD�L�1�����/p���J� ����ua,�P�|��H�@��2b��%��*l+���G��xc�"����wSg�j��w��^�n#�^�K����]��ː�)7ޗn����ÄV;���u���]��3Ό	OhT5��=L���mŵ��v� [_���C�h;B-���^<z6�X����'�ϵr�j���:k��s\-N���i%T��Jz;H�;���"A�
h�6j�<)ZgW?c�nWp�J\�8��>�Ag��=���X���:�f���xk��0��֫���'eտ\�%�pN���Ǫ������S>�����<(��R��J�q>����Q=Юٿ��4��3��P��'_p�������,|K /�t�#9yj?�:������G><}�[�ʗ�>��+�+��Pvk/���)X|���W�|��g�����T��a¸+�">7��V�>���ƫW�w�YO"��Ջ�T���_���X�)��f�E.��,����	fY}x����������W���S�1�@��~�?�+�$�+)?[�d����j=��=��9~������g�B"�Z��~�5xښYF(L_*vc_��8<���g�=/��令ߨ�K�׳eo�����h��R,��~y>�:�hp��I�,t��Pt�O,�]�~�G�=����{Qv�Ϝw~oIi�B<��f�.%����3UXT(Uԙ)�Q�P1oB��c����5rӐUN���yg��Ns����b7p�Vo"���͌:���F:���-�J�q�>u+8m�m���ެc�}�~�7�K4r�}����`Y}�yvWu����W^��b��f��,F��[�(�q:�J�
n�ܪP���J\+��O,���/V-8��t��Ǉ1M*�b%�t�ʨ��RXO�T�U�p,c+� �̋פ������;��b�T9�zPto���O:W���"�e�����w�kq��GG�͛�Z�ch�>[������mj(�� �����G+��dRX*���aY+W)m�0	)�}�ꫳ���x���
�wߞ(ڬ6����!�#P��Nᭂ!0V;�����p,����W"X�i��ݩ��6
�P$��s8|������j��E:�E7������ܶ��c;�{��p�p��m  ��np���n�g���c�f{01�@T�c��ҷX�Ya��(S�3�T����A9Qvgz�/��c+(mB��w�`B`#4ќ���K`�J���u�HO��w|�';�o�FqT�Q����2�T���x�UWM��k�6}�ߘ����������������|��vU`3-J�kƄ��CӦ��$�]��Y���'?�f�س:,���ק��p��E7���s��8����u�Pz��kz�l
/H��J�[�|�Q����,�m��O�W�Nś��#��^��3yW�_�\v�:�%}�zU��s�3*��O>5�~�����,}��W���Z����{)��?|U���7-d�M\���:<s^���j�K�U���+%e���a-$s�j�	]wx@oMs">)0���¬%�穧�j7��{r���5�|��������0w�ڙ�V�ҧ�(�?��#?.��_+��T�vm;��h�'�{���/�r�x�x#�r�ߺ��SO�L� �B/�jG�B�x�PF^��j��Ͽ ���1&}&�q�5��}��i໛�q��,�|����1(���v�;l���M�Իh4�U4Kz��b0/�z�|�W��ն][��;u}l�g%�6�m�]I�)�:�vnB��y�u.@w�tE����V���n{oˮ���d��c�G�A�
Q����)�"%@,M��yJFV��h*S��j�U��@��}��H����trO=�6G�V��Qʀr(\/f�T>Tg��(�Rj5�����>2s+O�#[eTG3�S6��	���iV�K�ۤa�hx`�/�y�G9�����>�My����>���uO+?����Nc�.8 `<����^���S:�w�smK���V'5% ���W��wY~�h��+���Ƨ}�g�O�����[JЙ�F:C�_%H�N!��8����xN���{M�m�5m���ca@)0_|�gE��Q�|?�/�c����iL/���J}����u�'K�r���L�G���V��mV�-<�nK��}�:
��
��yFK�'��|���}�_�.�ؔ�/��^d>��`ҦMY��*W]߭m����I�7l}���-C[@\�(D��5����4�͢w��ʋ�t{(���۽}%��i����7c�B`��x4��)��fm���]��`&C�����o�q=h!�PQ��;�|)�[=Q�����S��J��2�8mO����X�w9?�i��z��9��:Q����� ��K.�����F���+�&�G���Zh���{,�艵ߦ��򖆲{vѾ�zz�-�m� [�H�3e��¿|�cEU����R�7���ovL�=��8��(��ö잒v5���
�HJpS8A7ڛ�N�/��
Ko���ge��[�'z���5΅�eX����/�����ۃ̺馛�������@֭��j������}�)�ˀ�/��&����(}����_�r�c��g���O~��@w��.=��|�p�w�\��yf~W"�B���:rW������ұ������w�i�$� ��P��cJ1֗��}�5n�ݥeW�����2�kl��W�鸸3e�|B�ۢ}ib����U���Ln�%c"?g���q�`����~��A㾽{bpЗ���s��3����s,����Un�q�e�WpZ�Hm�������8�/���WG���8H�������7�W^���|���,�uW���i#p��Ms�ÕS�����ge�+e�~$���6D�z۝��w�<��F�>L��!��iD����a4z��g�y�t���M�w~�����W�ì>F ��Q<���(�s:8ss�4B5���%5
v={�E�Xof�/dl�i6_���7�h&U�q(>�9u#�@`Ź3+۽�k�7_ʡ(*"��yfg	��F�0�g�袋� e�?���Vn�TB�ʢ\��0��PxG�p�c#x�ZG�L[����F�φ�3*���?�L�X�~u�j֪��zl�K�)T��/�G�ӱ��Gł=Ӊ!��g՗�˔�k�,�2��:?X{d"�(!�.�	�
r�C]���}����V�\�6�l~0��ڀ9v�Ú.R"�ř���+�xJΉ�I��Y�z�Q�t>VX����/F�I$�юz���#R�|1�K_�R6��*�j����S��KY(b!	!d�ѧ����3M��h#�l��U^���L��4eҔ��W_5�����*S�ڮ�郺������A�ϋ��)WT�z�߫0�:_�q}��H;�nEwcV�_�᫃g�/�Ɨ���X��rѣ��Y,tϽ�N?���Ӎ7���>��jVP�����{��6�� ���h��K��;�w�]�XE�X�;��_�w)�d*Y^�1�0��D_��:�+��xK�����e�=Ix8�,x�1�da{���6�������BYze�+�0�Q��_�L��s��@��W����7� @�%D�(��J,TY�]y�ۻ��-��/���|�Q�X�� |�����������t~ɇi4�Pp� �ߗ f�_��~�p�Z���u%��[�n;���Ԃ�}�?�3�g�s��u�e�r��j��)O���N�)nxU?�G���N	�����v_(x�o:���E�-@r|<������y��4��ږ�B!�W;����g?��t��7nx�wJ�6�n5�z��Y��O��t��7��|�4|��°��&�u_�.4I�XI������y�;[��B�u�4?�9��w�-g�d0���9d����^��c� �8�V��#_�,~*H���CvW�E��1�.�A>7��v�:fں������ˠ�}ݫ���``��� ��j�2,�g��5���_f�C��/��r0\V��,�/�Ŏ%�)��М�f���'O�0����y��2���W�>���m\Uy��\����s�};�룵����}�m]�?�C!u��\5o�F�e0h˷�1�.C_�}��h1�Dot*���&�{,�G��h�rk��c��t�e�L�}ֻ+�4�[n�c���3M`�1�>�P�#t�N�*���V�
�w�ھ����X\	|��(O�P�Պ)ar�[������dT�����b��l�u�3=�ѳ�Bft�S8�G�<��3����R���TP�3�R�ü�_����«s�ZD�k1�=�Yv���´'SJŠR��x��v��P����h8�N��ć��+�bWY�l��MYN������3m�p���)�r,�z��ś�r��۪�'T�M�Ø�sUٕ'殼1#Ltf�G�5��9�)�8�����أ��������~���>&��8��Yٛ���Pu\�Ի���B7M�C7��\�^�)K�����b���c���Ώ�㙖5=�>�qx~�bw�;v�Sz����;}��ߏ�U��u�T"g2]\�|�-b��� �_���[���%���Z\��>��W�EQ���.KK�}�22Rǁ�5���p׈�R+�?��R�}���oM�K��֨�K�o�����c����۲������o����`��|�&(o}��.?Kl@q�#�����E���,�A3IfW$4����[�
g�Ϳ���|��!�Y�5��&4�= ��y�;}�3����ͯV�: �,�2�+N�N�?�H�]}����>�6k�`����D�������˿��oT<��s��4-d!V�{��|�u�싯p�wdq�w���(H��X�fZ ����Ι����Rq���XQ*������^��0
�m�ݾ�7��>A&�^qk`���N����M�����3������ߚ>V}�0�o�A�X}�c	��{(e��{/�/&B�d��^~��/U��48`�������ģ�<|��]�i�?J?�ȧ���Q�W�x�++f�Z�p�0`�T<������R�m�̽:d U�K�e�G?�Q�%�O�&[��2<�N�:�p��J���׿1���A��F�a!��w��]^����5N{q��K�]�P(��湌5A��0 �[�간U����=�7�]�8'{�/�5�G�@QK^� �z���w��?(�}ǝw?~���k߷է(ЌN<�!��b�c":vo��S4س��m%��4�5>*&��S��`Rna�3{�p��gq��h��Կb�����l�<�gx�s�}a����WGA_9i�Iq��p��|{���CӠOz{�����_��3�2�X���p��>u�(�Qv7���p���k?1}��^����Ӷ�%�i�
nC>E���o�l%uۭ�f�r�8�m�p�. !U���m9ik�E]ES��vg-�ߍ�B��y�2�@�R)V����߬FM�0� m���q����F�Q�w�is5#�)g:��ڼ۔����`S�ԫ��Ff�)�5[��w߽�Qz*_���K�/�rJ�,���ٜ����}���l��^��,�1��I�E,�=�p�:�z�N{���_E��G}$D�^`�i�t�:�G�+�E_������#��V!ՠ�mM����c���m��Rƺ|�/9��'?.XH�(�@�!ȍ��V��3g�*��s�Ъ���V�ap�Y�'��kB���p�0vX��N�_���K��bnD9���u}���6���?����Q�|��S��^Y#L{���#a�_��m'��#������Z�����$1�vpPe���M���c�](��k����oL_�ʗC�I��.1IBX�b�������?�a��Wt�f�ߞ=��(�{���:@��&��^���_�]T�F`��>�zƦ�y<K�P ����*���or`n�tyx�,�sc\	��e�G����/~.��8%8-����/��ڝ�Bn-��R �G�`|�E��N{Ṯ�l�49��3��P�;؟��+���b���(<��[n�����f+:|d��W������ݾH�W�z����Y
����7Q4L��ٟ��tK�W���	?R_�2�~�_�>��d�;������OC7�f������0�/�'X�� �@,�(��t������_��|a���ڸ�~��)�7'���Lj�C~,���x���#H�
Aݷ���_p���h���Վ��:��i�tt	�Ֆp_���r���=��E���?�����Fhv�Y��ml��h��!��p�=��7�롹�K��z����ѿ� �@�Q�3�����#D�:,��Q�:�1��I䋰�۱�s6�ϱ����c�Ime�V����s9{{�+����q�W�y�bh����j/(U�������c�,~5Wg�;�8�À���ޤ|ƹ�]<���j�O]�?�YyW��<��f ܜ�����dZʂς�N�B�����=�-��6�� �@���8H��7��%��(��� �T�����rӽR+8o����</"�x�qE��X��5�_~����O=�=�	B*֖�sQ��)$]�U�ߞ����,5�xߛ���J���B[�{�`�Q1Ԩ����7�L�9>�/����FH�^(�ʂ�����u�[������|d��B�o_�̕�)��S�M�J���%�=���rӦX,0~�A,����z���4��1-,ԍ3�0h0f���`-;��!:{�n�F9����]�)u�8q��P��V�������m��i�3;�WY݌�XvC<���H��"�l����i��ߐ:��
숹d�N��"�(���R6��?�o�����K��ˋq�̂� �5�H��f�\�c�d��b�&֠(��#|?��2"?�E��{M&�8,"`A��Փ�Uu�z~{����J���F4�k�̰-��}~c��H�)"���ǈ��ѹ;�Kϱ�����Xt{Ԃ����\�Cŀ(R�=��F����J�׮���+4��i�\S~�J�H��RW۰���*V�]Rt|�W��i��Y�s�KAY��ئ�����R4�	��k��P���Š�2\�+|e�_qQ71��"�+��}$���׹`��,R��/��)��R�P��n���
JY�����8L���.�� �h�[G��&�eÂ�O�S����.������-�䞾7�a5�q��HW��+Ӎ����n,���_]Uy��S]�O}d�R��r�j��G�zʮ=u�^�s<Ҵ��0m����\���VN��.F�C*?���}j��������PdZAqy]�:���S�yM�{NQ3����i�1�͛������.�h���-���crNqK��捱�/P=�2���U�a='K�������M7�4����e���n�q����+�l��J�@ڳ��짉?�hf��-`���UD��27LǐC�Y0���zuڽ�ُ>T���?������#\�>��f\���®�	������yYjBt��&���3R��O]�V���qܿ7mN�x�9ک�`��;�T����k�|�%1�U�m>�P��O0��z)��W^�h���4����.W�������x{����eP�(�+q����1�8���nOg��a\F��'#���1�D#C� ��}kLGf���|�R����Q��=Zu|j)p�jPEJ���7Fɤ��H\���X���;��=����` �Pz	8�(FV�*��!$�;�hq��{���r}���{�!{�����3�bI}��Ґ�F��:�Q�3��Ye����۶��o�IV^̇Ŕ/�%�V���.t��X����_��|�/�x��X���xPH�Av'�AȫT�ۓOٞ�}V����l>�|��*�/r���ۚƴ�tL��~2�q����c��Ci�6
W���{8�q�ki��(j�����RY�F�y������>��hV����\	!�6��w�{!����,<AA�����m�c$*���%�kO�C�����4�s�dX�9V�(�{���k^��A��׊stl�'��)o��'T�>)-���r�ǯ�r�
[]枀&�ƀ�ꫯN9���B�����c�m�J'��mglb�Ѓ�{hڳ{O�v��3	��9���<VY�}aӦj��y碇-��7{p/�W_姺?n����3�C� t���W�QgA���H�ߵ�oa�F�eն�5[��P�ع+��{��r�][Q(��aC��Le5�ﴹ��$[�����L�iS��o�����g�	����� ����'\�Ѣ�{j0�*��]qE>ޢ]��ઠJ�3��h�,�s/
S�Z�<�E�-�q?��xg]���n���`�zwF�jz�C��k�V���XE�P�Q.WQ|��u���_q�y$Kt�=�Ԏ�x�ɧ"���|���Q��{�Rp���O������+��[�+_�,��Q�؋V{W��`�����9�5=33^���j�E������1�0�
�h�cw�l7V�_�^�ma�O���E�'��1�\�]O0�wZ>�	
���ܮ�j���}���F�F��*R(g�)o��e�}5���t����5b�;����Ǒ�ƌ�{������yV�~�Yt�._l�ɯX�cH M����*5+���<+����-��x�S0��#v�s��}�B�U|�>�c(�O���)��K����K�����x:�-�W�-(��:�gfQH&��Ȍ,����@�Y(EV���e��%�?���rM����Fޭ��F�(C���R��
@8b��:O�Vdqe��vN%���Њw>6�Q�Y m�C��YJ�)ӱE>��!G��F"�C 3a
�FAΨ����JK�ӈ���OM;�~:Q����]��}��r����L��r�t˭7� yp�[̺F�܆N�%&t2�&�a�A�c�f�|�X
.���2��1��/"�:h�c�9������^���2=���%�K���s�b�v
�f�m����
�~�;g㮅\����W⢓̸^��7X�y�#_�{ڐ�%���Y�
�X�~�颁ބ��8
Yաi�w���/6:�U��Q7J�loCwӯ�W�9\@�7\�t�ݿ��(��rGĨ��VZ��N�#��z���`�7*�m���pT1D4�j��M�R��9��W������0�{	���ي��������O�*Vʈ6櫌��>������o�!�ʵ��إeޕa����̅��`lW�UE9�h�ڇ#�?��X�*?�57JW*V�A[��vVq����{��.�L���ʢ��ѣ�*�������ȷ��0��`�W��Rv��"]�Y��8��?�D��x�L�~�*���	l��M��*�k>~M��8�����z衇C�ʦdq��n�x�[p3�5`Y���`IP�pV����bɭa���k�W� ״�v�~�E�8LH~Rt�,1~���:�[��ƀ81p̰��f������U�rF��K�WD罺�?�!�O��=�?f
��A?�ݺe�t��m��qw�+�v�O}*>���ԧ�X�ӟ�t\Ն�ba��M4*�q��Jxq��I�����l����˘�-�����B��y�[����y+s-g���"6�=�����kQ<�~+���N��v���N;�[G��v��c�\أ�`O	�u�i�%���2�\�9�gy]�[�p��5S��;N���X���1q.ۻ�������6N�񑎬�{�K��J/�ɘ���k��^`��$ޑ��.���&�/]1��'�\}'eW!*�s׳%`�����! \��j0@��]$��i�3�3gS)x��{�=�k�}�b�ϖ������M��B"�2�I�u	~B��>p�`���Fk`㼏 r��}�:�^��Ixa6|wY0����M��I��TD)����Se�Q��q�nVaS6{���@@��=�r�h�x���h����R��z����`:���Pއ5��6�>J��|3{�?S���;K�v�a��S�p2�,�<�`�<�Ӯ��xt���\u^��Ӡ$h�&�������NQ�5a�(vf�0.Y�1�N÷�b1���DyN�u����/�@�6G��,y,kF�����c�Mi��ʺ���a�E�СP�Z҅\��1��#�S�2 �]�o���(��?�|�����I4�ﺂc�^��`U��e�^�YV��������w`��Vy�#4�e�:�Z�nKP�K{-�f�>��<����Ђ�/��������/� ����Ek�9�h�}��=�"qE�BʮD�<ʉE�B����鋃��u<�*�<E��M��i���ˮ�D�T�]0F�j�
i�9X�c�,��15�����ǶRď^���(���}5�}x���K�|<�(K�©�ZY^�ĵu.�p���מθ�̌���Z��������n���d��"a`xw���*��cƪ-/�M������S-�z Lo�L�����@��<�\�ha!T��=_E�Ņ�D�dx�G9��-�\w��?K�����D��Gk����ɌC֍PT�y�࿷�~{]�1v	�����ۈ�������zj
再�Wn��� �g1��9�yG��	��`�s���QՃ����9_ױc�J�%��Yp����L龷�+�S��e��Rn� ��ڿ�R;�L�W�\�y_ʯ3�{M]^N�\ڑN.�[�	�c�<��E���9t������+��������!��]\�/Y�ΏזZa���Ñ�(g���r��bHK�T�1�CG��1{pL�gZH��.t�+���:yk��D�qϹ��x��˻Zvenc�g��/'q��Xf ����B�д��'������Ҿ����;�K���O�V�_{`��(��-��X5�ߗ��ۍ�@�Cl*o�/8c�5��;����Hg���i~GV�]�J���t)���}n���EN霋�0}X�폀�Y��L:��(R6���m�Χ�;��߽��i��b8��7�F)��)���	�06�����R��ө��p�z�'*>�����k+��~����<��zϠ�`A=B�U\��88	c�p4��A��3��|>
�1u[�#���ˆ�ň�]w��J���(��Ԗ`�� `]��g?;����ݺ��Lpns�a�$)B+�o�.z+��F̀�k*QxY5.���*�V~��]�Q�H9���ҏŝ���aVu �Ji8�,���+|�R�����-Ş8�c=_?d1ߡ|���<X<`w�'�T΍�-����k���
mW�el��?)�=F�8Y���>�Ĵk�(���Ǣ�`�އ��)��W�����0�����͹0��zV;�6�����L�SL�(�Ӷ���t�Mᑕ ��cu��z-��ڧ�4?e���w\)�V�s�1�U��F(e- ތ�#�<k�7XcE��`��Ry|���#��}�qE���*Z�����V��#�	�O�!r��[��N�z�s�3q��ĵ�F������v}�������x�;�`�yf-�����+����5܂g�7�D�S,��������i��-2���<�"�*tQ�~g�o�uo��,w���Ce'��g-�CS�*�BS\�(�h��J���QD���/����|�~��ŏ,��ߟ�~B�mנV>��\��sG��`P�(/4� W�9��}�C��yc�j��ը?1�0ڸ����%�-�M�]�z'M��"8���_�O^��U�����*}��l���Y��W�|$��H�E�4�πYȳ���#9w>��1�ԽQ�E�_�gO�Q���c��o�{P���R.����[�Kݩg�xή7��\|	]�M|C}A߮<F�]��.۩���ʗ��7ˁƼw�9gM����������ƀq�D�6��96���Q��:�:�ޙ��ԇ	+�*�V|T�����=����X�)��!a�[���E��xu>^sX��ӌ�5,�{#Q^苵e���w��x�=�Y���j�Ր��NG������O���a>[m�U\R��`8�Ŕ�8F�#�$���u#8��=MRt���.�3e���������JaM	�U�-x�7�U#�kKP�x���|�3�)u6�s~�/��V=,���a)���-<ZțjS���a�q��P:��R�X�R��HH=����ӗ+�zY�J�q�z���Q���Ğ�� YX�\:{#%��1#!�Xv	���
���jzp��!D1=8 ��ù� ��^zY�ùT�y�Y�T��SOπ�m�~�WMg�uF�>��Q�����G�����v�*>u�T7V�S���]\�6�9��-�v��|�)H��) �`>Z���ʹ�����<��+�i��]�2�G�/�K����,��z᳣j`��Z���X�Iq�.,��������ǯ�&��A��8�A�́����/«�m.h��j��U�PȽ'/y��EA
�u�]W���(�I������_����!o������졒����J�/��	|o��9�{��y�K>a�{�����}��8g�n�GO�o����<�S�x�*}\������������x�<���J��3}�K�6�ZX��U���(��W��?�n�ۓ��P@�;ۏٶ��3������2���x�w�������NWRy��2���;��GPW���F�kY*�S�" o�g�>��N���(Z�6��z��+I��r��r62j���>8*,N�,�/a�s�-�곎�W�j�F>���)���ã_{/4[�Eѵp5y�}��g�s�qQqQ����.�dc�1�Y�J�b�o6l=;!�/7��G_c�����Jpr��t���2�q�H�x(�©�~�O�.e�B�X��N��+��䴙��˵�g�^����%��t�B�7b���{�z%�0:̧	��Yr{D����W�q��拄��Aϧ�<@FI��W�B�t-\�[ܟ�sXI�r:�^ss%�t����t~�`�wl߅fc(V�a��f�Ga�M����^��Y�;
%!�Vi0ʜŇ�L�
��u
� ;2�,!��/ε{��(����>�������X�N'�(����Ǿ�|{U���0�.�Y�(w�qg|��љ���SϊO���٘
b���w��)�r{�e�?ʊM�!��9��E�����i�c�|i/eP���2�6�v[��g>��,@�6�lhj���N�|R�kC�;_"d�a�R�n�.Q0L�U>�q� ��z���L�0nDi��U��;�c����)�` ;�W�^$��3"Z������#�z����>��ӥ�<�6��/��A���|�	�f�ò��R[�9ĺ ��GEw�y7tTiG��^fcƳ��N���vB7p@i4c�3H2��F�����e��(�D�d�I���k �=�E���]
�Lˁ#�)y�q�Nx�eW%�'j/t���bFk1���-JQSfD{p�Z�0+q�c3y���Qf�W�U�؂R�(����Y�Wp����n~��w�-�p�����%iCtuo)�ܕ���}&ܬ^,��Ό�P�Q�<��-���G��n���1h��^an6a��Mǽe���t�y�>1I*�6�d䵚~��ww�ƞ�'H��wg���u��",ʚ�s}4a��X��(�����M�ߊ�W����nf&s�9���=D�c`��2�����[Fy)�;���x�1��B3oO��fN;-�Oݾ=Lx��[rY��:&�y��s��iE�-^M���z�b�y�}v�v�ϧ[n�3�꺟\�_P��"c�_S �}1s^(�i�Td����ɻ��-����%��O�U�(��8�2,	j�_�"�:9\��{�=�5�WӮUNfae�XI�8�w�c^��+���;_�U���V�s���ُ7*M�Ҝ.r����j�w>��B���enr��c�j�F�V��O��W��vx]��PpGyPd1b��R`�}^v���i�G֦0�:�>�r���xWk2�����Q�����jcb�2�=b�/!afSn�X)�F�e�1%�'5E�pXh��	ڳɲ�w3Z�9ÇA$�ʻ��t���O	��%��y5�tﵟ������?Ȼ�@����D	�l)����+�%�pb�����q�?y��O<�T�(�1�	o�|�˗�0���F�U��ǥ-	fZ��|��`��t�P�p�YHx��vˠ��S�H��is�����x���2�հ��n���\
�����@�U%S���}�X���j�������}�HwO�����c�[�t����sAY��Uu.]���`Uw���+�����j�x�e 8�zWfĞ��v�9�ʫ)Kp���bGxі�O99�[6�e3p�;�6T�n��y��:.շ�p-߫�~x(��I�8pi;<b�[�g�qffYx�C9�p�w��<�rA�Wp�9E�s1}p>?*ź��ڃ	?�q~y�}�F�����@����k����'�t�z.�	>�fTͪ4m�O�3�ĺ6�m��$8j'��my��5_���zY��M��P��o>]� ���E�3��7��1mh��{m�`�?׮�����0�,�~f:��9_j�#��C�[G�}��
+�o�U�sߠ�l%�D��]��fm�y�	X[�z-�Мv��a8}'�
Rv�wF��Y%}�;�B����π���}�� �ݣ��.���0�E�W�,٦̀����੃�	�r�e�}�hP��0�f����5�o�ַ�+>t����㕡� ���~^
��ӥ�����\���Wቩ�[�P|����Y-�i�UҬ����
�U�������FB�>�+a(��ǆ-!�9/�|�"������
�3�j����Sf%G۔��D�<�w�Y�G���`5l�B�e�֭5����ٻ3���BHx'7�z�3���58�:t�k���K��.�1�X��
��a0���v]x{;θ��|����>:�r��.a���J�������ڧ�e��m�Y	�0�J�/)UZ-K��t�K�����������eup)��b�G��,��t��c'�j��M�k�!�F�>5���П{���W���n&��s���aS���c�,���O�1��.�|������RV/&�?���c,��hO�Ѿ~a����:*�P�@�_��Y�Ujۻ|(�m�m����󬁶ݓwxQ�sX��LrI'��!�*�58�g��g�����ICp$�J�=pI�nV��p����F�<y�M�@�������7:J�F�-�۞������+_�j�u�������w��� Y���+O��p+u3����k�)cʩ�u��S���O�!������|e�nl�TTgu�Z���N��;��:�y���5��:���'
�U<��1Ϋ.�O���M+��k�c���G�rފP|zv����
~�C�g��!/�^y��#e���e�7o��`�!�>�=�����f`g!����,Be%ד��ګj��a��
��`�T����63��Q�?�@�9��w�}���6�y�]���j����2����L�����z�w��vA�f�,ĥ���Y3
�AݸS��~>�S�qd�]�p��j��qD�X]S�����V�=@�x�|:��3�|^q�U�����,VƏɪ�>pi>3n0:���{�����W�j>�6���@�&W�w����/�Z����/��o����[4e���\4}�k_Ϻ�3�:3�Ѡ:Bx����(�SΦ3]	�2��C+�?eW=����o��te��-��c�1��,-���J ��4��"h�Î4Yx�X�#��2q�Ό���e�ޯgo8�O�[�	���˱���LOf��{ԳT\��G�p����>{w��������HЀ޵Q�Zn�QK����P�O�و�7�Vڈ��}1ҪcB�i�����M6=H $���{��6?�<���{��< {Z��߭{ΩS&+++++˜(ҍ��̮�A�:�����F�R�t|�GEa����*Xʚra�U����i����3B�}�hY���.��E��|��j()ESYU��>�7^mU��(i�������&#�n��������,J|9��@s�P��s����C�'�rAPȺ�Vs�P"4r������Nc3�����Q�˵:�����+���c�M�t�yl�AF�pWp��LG��|�^�uF�hQ|&����y�A��9��X;��S,w��u���k'��<u|,L���^W���5q�\�q>�8�����*��_�IWZUV#qi��LQ�玌�'��-:����I)���R��������/��tv+ɚ�������/�R����J'�S�Ч�\[]�E�+#�����8��<Wiq�ͼ��4'\>�Ўߨ��E��1H>Iϯ��U����W�(()��g��Yɀ�
�4�w*�;����*���T�ȃU|W���i�S^'Xh��_JZu,63�Ի%����uN�/~I�Ӈ��w��N� w���/������N)d܇B�Rx�ͷdF6��E��j��@{�_����ם(��W>9a�R�E�rA�P�%+�o�%�"U.�{�*+���lb���)��*?0�rء�e�iR<A.���L!��Ց�n���5��v��a�6�W��x�����(=O>�T�h_?����©n�	�]����N]P4F�����o9?�)J�qB���u�����8���ޟg-�o�&�W4J�_J'<�K��Գ��Ӡ�h��쓯>^}�'��?y�tY)K�ty��M�wn֩W��C�Ny��E�+�y�7}�ӟ�>��/L�W_`�i�ʱ���'�|J�U]��k�^�3�>g:�3�T�rRه������������c�~ک�dm�Ǯ�X��;?ۀT��&�G#�9�}D�N̑p��������.+Yz�t�%O����,s�:gpj���!x=�֪��'��Q���\J�k���{W�zRfB�*�9���$8��Fouh��`�׿�ԙ�%`�A�Y!t3�u�%c�O6[d�Y��7?���+���[2O:��W0�9��f��'��}2kvmPӑ���@�#��x�~�Rף�Y�+�[5��u�❊��HE!���c�=��+����e���m�1p���qj�-��!��� 3J�w��I����uZ�g�$��M�
]�Tï�qMX��^g�p���y�R�o7g�@�it�y��ʭ����z���6��u������mE�����H�U��l���44�$�*i9��Ϙ˪|�0��v�� t���F=WôL�@8����[o�%�ݞ%�5um
�(.����^sV�T	d
hJ�hu���K��\��x^9
M[�(�p�<'��5���<St�W	+�!�'���
_+�2i��W8��R�~,p��3�^8�T��	3,:P�yKD|*�g?�i��0��VUL�������2�?~7�8x:S�����r�R�2���+�\N�
�܈<�H#������;(�c�@�ĳ����w�⊶�G��<��<�/l��9N���o+��� 42��B5_ɐ�yϿ�Wz�� ��g��1�M7�\�}d;���qǽ?(���E���#��xi�<��H[[j9O>�]!�;�&��{�XaM)�~�����09J��J�Q��ͧz3h�:w,%�á������)06��4d�|�.Zxv�*W���[�{���3��)�����������p2\l�,\(��WӲ]׋<�~7�{�j<�����Ja����/u���+���,�}����A�{��γ�u8�%K5�K/r� ����������F.�5��J{���a��ıSMo�S��N�E�Y//遌�9r��x��*�lc)��I���/F�����#Gg�]:㌜�W}h�g8�WF��#K�|>�ӥ�^q���q���zgz���}l:����.�|���؟�vdUս����������ˆѪ7�斦�B��[A��
 ��|�O����#�e�+�w� ��Stu�H��|zY��>�b_�g>��|����ɱGYk��c�jg-w��'�����h������L�a�Y���Q�/8���?m��Dal�u�����7~#_�5@����ey՝w������KY&#�I&ׂ`�$o��AL88��/fH�X��9���c�}���e�錈wPv�q+J����U�zwȽ	@�(�A�_��ћ�Ah8�� r7����`,�,qW�4b���G�& �4��7��at����5��Q�~��(5�M	���ȵ�9�	Eb�it<S�bj��hA�T���8(;�sO�#��x>$/�~��B:��P��e}�4d����p�o��S��S^�E�ԟ����Y�z�k��D.h:>y��q���3�M��AyLg�(��g�(�q�ٓG�l�@���u���F��hV]D�V�>�(���:����Ĥ�J'���4+���ϱ$���:��]uf���:�ݕK�Di+�,O����SǮ��:���6��}��\���
#M�aG>D�#�8|���]�Qvo����N^c���!o�H�Й]���F�hEq?�������5����{����J��^�L�u�;�ĕ��%lB�b<f����/~ɳ�N#=u���E��[J��/<?�R;kᶨ�U��|�*�\>'>{�d˨��Ѿ����J�����ԙ�ԙQ�����,����_{�<����L)�.܇���/|�Ӊ��u�x)E��p���%���6��N ^�<)*N: Ї�2�n��b�v:���\><hY;������@8�K��VONָ��[r���Z3���1�9 �Vy�x25�g��:�{2��Pɏ�Q�����~Cn�7�N���͢/��?�[�Z������w3C.`�k�׾��銏]����fA�#�H��'I�y�/��괽�He�y�[��[Y�fO�ڱ���x�՟������Rx��6���7`S��|���[�8vs@�5à��VN���j�Ś��+>�e� �ś�p���%y�+�Xi���+��23lx�����.h�6Ӆƞ�����_�����M���<.���͇qd�ժ��}}��^�N���M7eC-z[�� �}l�X���٦k�sm�~5�v�-�]�г��3_5���>���a�8׵���`����{�tn��<�-��q;O<��1�1lTv9w'��dð!W�`�i)ŭ8e�T�wĐQ�!�b�CK�����
kd0�BVi���a�;V�hE�޻�}U��鐃�kT��1�qy���Jx��Q�ӆ��tsm�5���~ʭS3JV�>'�q��Cڐ��^�)�΂�*�wKȕ�)�Q�'����5	�I)+'�x����?U����p8��kP�`	
E'���S�dg�9e{V���?p�������T��1�<���r,�F�QY7��:W�h�F�_��W��|�!�S�N]8B��!T^{�w��{��f6b�i5�����V~A���R����?��Q�%���k])'L,$U?�Y�e/ׅ��=ȯ���?�4�p_wI���Z���v7�)������E�+���Y.���\��>���b�.xU��/��5�	#�'av��G� t��f!ӑ�қ˳�m��2��r�	��.�+�=��1w��� W����nU7�ÝiA�ɀ~����\:|����*�*4.�F��3 *y�gο� -@ҿ�>��0y�V��^��,#�ay���+��g��a�]�5`�=��ߜ���X����q��g�Lj30�bY�s�m6d�y��'g����A%�nO��C�P�?w�禫?���M�]�KP��\2�wn@����߽�9<�!��>��A�V�>|}Y�W\~Ef.�Hq�	�e��{���[�[;��^�OZ?��C� <���C1-Ϋx���"��D�k��,�,I��Pt7�h@��{����g3U,��礏�3?�9Q��������#��z/-�"�1_��bA6SaM�u�\9���r�J����G���N�(]-�e�m�ǯd�����A��5��������(VG�Im�R��"Ͻ��]�*P� �,MY��]�{��7�w�~Si�6�"o�ݙ�NQ>dd�T��b_$<���/;=k�m�vr��_�|)���ַ��n���f�э���}��WX)��]h��������ݢ��1�|���K//y������pn���|mWx��J��}OF�7��o�����,�a�֟ё��=��tk�|[a�Ԡo_�ƹ˷�[��/,K!;�?���|��E�C)�OOO�fM�ڬ�̅S��4�к1��QN�=��(���<���Zs�i�M��"������EZ��0��tL/ >Ʀ�Q�u�%�f�������hUh#v�9�j��0�Z��,\+o�<���:|#�51*��
7�^�dfʦ2U��t�gKa,��h	��^}�������Z3d����Az\�5EzLek��@C2�5,b�,L��)ԫ�O�U�֙�v�G3uCq=�z��:�*
L#?"����׿Z弲:���!X[c��#�L����BRY# g��fq3������y��C�_��Qe� 8������7��j�]�U�>}]�No�;�׊W���︭��n�q�ڍ��S�+9u� �K��z�,7��U���P�ʳ_�hm�s�K�w��t��0f. �4��������\ʮ�a�8���%����Nu�6N�(�v���Y��"�u���ޥ��`�:����k�Ta�u�h~��Hk`>»��r����4�(���ov���ď;��9݅��(׌�<V�~�r���Uv+J�ݡ^�\���lvTSX�>����E>�ʔ�㼜�jjއU5;�lZ5���:�C2��4_u�U%�N��� A(w��4]:�����'���6d(�m��X�Y�.�����Wg=�g����X�'�rs݌0��-v2X�k�Ĕ4��7 ��a�Y(8ߏ�~i��? ��x?�Zt�^���vӓ[�|(������A�4���|���,,��o;餓K��,�9��Զ�~�e9�O�S��뮟x����2��C�3,=���9V�gş���Yl}���/uc�Nˢ�q���#��R���E��k��!�z�;���c��S����$��Jw����1�KAgե�}���/���Un��|��Nb}1ަ���tė�j����H�e��ѧx��&,��e%_��C3'��E>l2v���$�/�ݙgV;�#k��=��ӧ����z�]w����@��#��Qd>�-��0�h� �����P�{tA}���-0�>�Z���`e�9��ƚ]��p�x̰j@u����Y��#�Ț��^��LS�&^T�UIve�[�/͟��M{IT#Eʊ����\����k�`��7F�jF:��C9��Bi_ Cd
�^�)��j����x�,vԲRix�R,U�
أFD{T��W)��C��O|����{�oz�� y���@�ϒ �*��T�2a��{v^k�����m%�_���R/����g��׈��c��Ŋa���(����3f�CB�@a���iVSx��ދ��K@��y����ܯ��+���C�\7��ơsU���h�6��4�X���;�-7�t����}�և�ʷrՉ�R2��]�wg�j�v�����:�vC�J³�#_o��
�U>�ky������8+o°乢	eƽ�����Wo��1%�Ȥ�^,e�:r"9WV���n���i�h8�U�/��5�3��,sa\+�Y����kj��7�w�v+�$͹��U�� į{����^A��jKფ��6�������2�4�ͅO޳E�&�VB��JmΧʪ�{�RAy�m��.9�ʮvL����[n�1�_�Q�#\�TyQ�� K�Y�k>wM�Aa�<]�)�=�*�P�c,���v������쯩>��QN=(���𕨔�d���$8��}��tnh�ShF�#�|�X��W��&6�}��gS��}��*��Z�1�_���8?��(8�m�J�>�zF�I>}�X^�vh�Q\B���Rn�w�.�s��e���3�s�Qt;,�/�f�|F��Ȍ�9��T�w���΋N��aI<�1�x�t���\�В1b�7G��1�,�bj�i{2�ɏĊK�����3��]T:�Q�l	�{�`e��Z��@Ɗl	�e m9�=5������m�ˉ6��t�EO�ܼ��S>:��'k����
���f�/�=������G��%��;%�-!���M�_}=�Ժ�(���?�e�yu3��S0�y�w�B�ׇU�O���(�f��m��.��X㏧�9�?�o�˺��%�Y����j��3�Z��ei��Ja�B��U��N�u�!�e�`���)^���+��D�}��W�v�!��a+�p��zvmR5������2-o�!���M��|K�pt��UY
�����ޓx#IY��[�����q�N�����Gqf�����s6��.�H���H�im�땇O�y�(�bFW/��Y�!S��3�=#8�5j2=E�Ր5
.S=�6�9��GV㽽��ݬsqH��G9�����-��2�����:�jTHi�85t��=[���lb�B?���P�a�ư c~vjZ�d	��N�tv�)'d9�A�&�M��\�p��&����ݿ�����5px �@WJ�5|��O�mF���A��$���"פ�7��yi���~��zJ�Ƃ�K�^�x5<�?� ��c9�qU?fx���n'sũk������;B���Ўl.kҝ��tH��C5���R"s1�v�<V�w��UG�l2�K�%��9գB*��ŋ�V���o�s�uo�@����.��=�A��ϒ�X[=6?J2�D����7���%O:�t�c�6���c�mz訕?���~fR����*�撟�'i�����-w��I��p��7^�;��C��H#i׏�p/	
-��|�qxv��Ҟ����p�ܔ�i���g|z	��w�l�X=����qt	H���|�L�c���ݯ�kQL��K��!���,�ȟ|2�d}b������R�"�|��~�����w�|��Qƚ��x��l��/���@��ʣ�+eg6ӥ~�a���wڅ�{/�]|t��+35{QѮ7�����=���J�L�L$�V�Ze�t��Y��4^���{ ]>�2>dBIh:>���o�p���u�DW?��u܆�Wq�]u�8�]�w@��)��L4��������4M�P��p5���Q>|A)�5��إ���@zҦ<2�(o�j�P��48Β���,�>�-�p���^�H�?<��_7e�pu�Y��=i��L�[�����h#KZ{G��N�Xkv�1����ۓ�/Ɠ���d�����i��+:ɟ���k���P��Hk;�q�wn���J�a���
ydM��s�6�}�߈��,,K7~���+�����:5K�\�����G9�i����O<p)�>u�p��Y>��Ȧ�g�\�o>[呧��9��!�?���Wx8���f3��`�8.���|T��O}*3��}V��),�VmI�Xf4x<����r_u`�i��mۜ��g)�ǆ�N��{�=�уl	���J]0I�2ڝ�wֵ�9I�2�u�Ϯ���?����;ӟ��VG��	�QqF��V&v�X{�p����ᡑ��c�=&D���O?��ϦU%��~0}����o�?��3i,ٝZ� `����|ݯ0�;�
ʊ���d섗��5:µ�۝�N�Ph�P¨޽�N3?�����?���W5}���|��rcM#��y��Y�N ���V4�~��Z ��58PC5����(G��s�5p��Y�Nd�9@^���8��z)����U��?kp|���G���.�5��KwhMs�.�`����M��0�@.�;�6�����G�x�u�U���^xyv,'�J���3��-���0?��#����ƲT��\s�ĝ3I�pQ�\��\�^)s����z�m�-�8.x[�݉v�Ȼr�I6��k"��ډ�=�8�`���5�ɭi��kz�\���3�E:~n��"ͤ���b��k~��u�x������7`��ke�R��_�i�µ\/����ʒOKNz�<�[~:r M�G�����r�䞼�������38?�2�E����>��(iڒ�)f���җ�4}��_�c���պ�}K�~�r���j8���^�%�,V�,^qT��x=����Q���/�y6��
lӘ�.x��v�x{��PrX�,y���K���R��,4ǧ��\p������Qt���sh�z=�r��W�����)8�S��t�x�Ӗ'cH+��v������;
�x�Hk�?@X�����i���q�!<����k��*q���Q�_����R�r+=��>?2���o70���Y���1#L�30�s��Vŗ�p�k���+�z�����(V���$��fE�ZY��h5q��,��wy�]��MS��r�Fx�s�M_hVϡ]�o�]�?��"���6�&�~���B��&j��~m�ފ�<��TY��ƛp��8�����eN�䎙��W\��$t크�'�����[.��9}Te�?!׼����B��mI 7�/�D��YmU�%�Q�,FfU3�f����^{��}�Q�|&��m+0�2�a���/��.VO�4:TѦ�Lm<��#� 3�S����<���0_�	1?43�ȫ~*��ǜ�S�p0��#����cY���X�"
�
]Ú���2���q�m�]wܞ#:��D#k#�t�&��Ҁ�����=ˬwO�lO=X/�t�Ǯ�?���L�����?��_N����U�ۧ��=g���>7�R�/yQ�u8����
�����7������ݼ'`�MF\U/ct���p2:����b/��� zr:�U�<��6U�Q\�<�d��r4���R_�% tv�����]�[��_�6��@
����͂nc���'�Z|�«�H'Wi��\'�¦#w�
IN��,๑��'(m�S���h6��P�f�v��8�ִ�Q<r�\:�L��{۲~��o%��E��fn�t��2Jo�0'/�;�\X��`���GS39�V����P%;<�C�3�A�s�@�S>ӻ�޾�l�, ��²�X:Fٵ�������t�'>9]p���ѥ@h,a�Ӊ�#Ԣ)��&� h�_<��5����x)G�V|��}}z�]Kg��i��[[���$*�937�,�%�A���kX��f7��Dߛ|��Eי�{UGlɖ�e�̭#����SU/��K,C��v4�9Î~����o	�|�C}��}����s�S��@?rQ�S��A|<��+����Y�V��m�~�����#M����O<|,��Qª��g��F�{��'�tQ�]�b�nn�G�^?ʸe��t�j1X�X�h+�R�F�nY�Lc�@�M�_�TgZr8�W�(�]C�h�{�ωq��1h����ۺJ�����N��绫�/���?���x�)����Q�������Ece��K�A�Q�'q#M�c�/���nj'����
���Ӎ��`���n^KO���}E<�k�����ɱ��\os��CJ�[���D�V�,m7����@*=���kg��Qe������RP�u�w�j��*�P�X���p�����m�����=_�1m������.� v��������N�f������y�ţ�8N��:���BzR*6D��Аr�X���}%PU�������;���O�	͆� �}��MkB�z����b4K/@qҥxhx�j��U��	�b�t*%� �n���g)�|���M5��%^�y�G�#�.��V�M�����Yu��=��8�+�N�M�,fĿ)l�jz��k���h���G
n(`��ݪ��sB�[yv]-F���P�s���Bc3�8�
o�L�ÿү��I�#��;�n#�A{3`�O��qdi#�[9]	��+�}B�a9վ��^���
7«|���Cp�"��hv�L'�O�?�$a�և q��;�2����
�4m\�n�d����>��W�䯍=�]w�t�7F;F�`�Hk��q��c�8��9L�Q_:6����=l��w�e�]��O���ed	�%6q��J��D�(��_��@�����E�\:���;�B��(tO�{�駦�J���zo����^N�s�X�5��e|��r�t��gfƍOμ����a<����+?�Vot�c�o(�K��pUW4a�d��`��{�{R���{��Sީ2�Z����%}�˒	˜J�/EX_��k6�GjB�
MQD�}�c�(���,����7
��W�r�۔��j pr��,��
�㪾}�o}�[�������W�^\Z���h�� |���%���pʩ�ۺ^�k��7�h�����Q�I���-|��cG�V��Q]��S�څ/	J��馞i�{[�Kɮ�m�RG�=�Hp��?��ӿ���~���?��~��r/ox��G�ޕ����_����sR�f-�oߺ��m���iLh��;oMO?�t��w��v��o�I�߭�������������l��;�<�Ү��Aߺ�� �q�7|�_y� �o�ޘ���Jܪ2w��r�VϢ�IN9��3���?�~�7~3��Ё�/��P��R��Q���i�k�H��C��bޯ��ӗ������ϋҦQ8�㙊Бd�S��urs>FI��$mSy�����{��{���<����XƳ�4�3����MiGAf��P	��G��lZ(���Hwu��Ƅ6�C��
%�\�<���/�g]M�8[4e�rEC�1��מ{W\G��a�zxțv�@�ԃu�>�;����W����f��*%��U\����D��nϛ�6Bӵ-���3�,?iz�F������%E��gd?h�+��6C�_��x�s}��ͥܨ��m%l<�>�n��9z�{+�|f>��*�~���f@��p�a���7�"��ʒr�3�r����Ov@�����e|�2�oy�?8.O/�rw;D���Ź_�/7���c
>�	m�S���u�.�	�c��o����(�6�(��/����7���:�p:A����[���y\�_�t��1�oU�z��W23�;��+�=w����/y�t��w哞9���cub%$��ܬ��i�F9�i���ep�tFsy({!�z���;���]r�#�guyu��^��6�W�����`��'���ĵ��<�M���\#�Ce��<���� }�����*i��#U��Ja�Q��G}���h�pXT���۹�]:�3|�A�֥�^\����Fv��;�KaL=ID��m��F�%�m����^5�t��w�P��H`u��X�g��~4m�� x2��r�x��$��'?�+a({�Q�̬I�Èr�	�g�*9��Z���w2[k�V�v�9>���S������o�\q
ôF1yD!,��M^�1����V�<�~�"���E��m��=}g�]}�~���W�)���.d_�k���GmT�����/���|����6 �"	F���Ɨ�X��vs��M\x�t'T�NFj\��ԖK�;�gy�x���y̦f@T�ʧϖ�{�}�Ԡ�@�����KЫ��j��츲:����+p�e�s�TvE��$`nf;�H(��x��(�,*��b�\��������Ha��F �1s��G�T�t��s���6J���:���gW��K1����)d-����4Cк�Np�v����9���9�	St\������ʝ��3mp�a�f)��h:�R����Z=#�W�5���Р	c���u���Ό�]���a�
O@�W�Xڒ�f�Y�M#�������O3��22�ơC9���M_��W�/�KYl��PP�]�U��+?����(pkA7����i�0f�h��_�o3BE��@��ǔ�j��jx@y�kH����J�Ė�u>͋\�@��x7���q�!��7����������4��g������9��K_��wr�:��$��t��0�\#��]�'�6�?�9i��q)^�B�-`(�xZ:\�Lg:�������Z��u��T����ޠ"�U�^��[�m��`�)�R��Oy�"��rF@��< ���|��7�(�(Pߎv�GA�w���0�LZ��o`o�A��0d�Hwf�W�T::����!�c��^����xY�$?��'��0+���k��Wv����*>��g��[o�L���@���d�ۅ���j�o�:V���+/O�Y
��oWgV�)H:��4M ��'���p�`�R���%7�wpX;�u�h�2J�O<V���ڧ��=;�������*�*��̗N��"=��s��.����ӊ����̞d��
��68������ôK��\���:]v���n�k^Ն�?Z�7�4�x(�R��s�^u@qIy�^*@�pI���9v�I��Pv��ӡ�g8r�ȥ�^��B� �̰��C.u�����k*e[�J��jf`)�֢�Lem��#�~���Oi���b[:h6����RB�_�	��}7�V�n6)�+6E�q���z��OJ�)��<ֺlhi�MK��k�<��'?���/~%Vkie�S�)��3}���@qXtu�v���v����Kn����e߫p�u�/8�g�ǖ�o��^ӁE�[��AYG���i��<�W����
��� J|���i󩧟��zf7 �0�#10
9����`rD����s��JƸ�/M�h���na0��0A3&�S�hBv1��w��G��1'5����`������G"E9��Yl�ά�Ύ@�Q�4�54#�y�V��֤d�n�ݎMS2�rX�3��͌ۦgJ0>��c���7=��#��}��F��F��`m����;��}�{�L���t����{S~�8�>/�-CШe��9�r���z@sӍ��"@��֚�Q�?��3�:�C�ig��l�1]x���GO;m:��j����<n���LϨc�*��ӌ���:����-Y�9�[C�!`.�o�jX�)��V���SkЃ>�P��h�;�^�����`z�qZ~Dφ(�����ٝg��x�8iؔ�qT�x��X:*�љy:��F|�)S�g�������ߺN�IL'�j�<���*�d�5���ukќ�06f��s;�nӑG5��)�s�>�5�xM��g�|]ܜ8Í�R��&��:
9��4J�H�[�Kx�掺�BT�k男Xr�nK��QЋ�"�f�ν3^��@����:��I��k�7xe= ��~�f\��+/�gM���:d]�<�˝�I�~Q�_���%�t`��ťL�����v�җ�<]u�y���Kr=��s�SN:93>������e�B;��N������Ev����wI�"$�ޙ~������G�%�Rr_|����o��B�g+W���\���lH���h���2��c��z��j�Q����瞙����^���`�9���n������g/�*�$�0� �g(?u�N��1[����28Ŀ�z{>�.��z�zMrx�\�yn������Դ��O�^����ΣB�9�O�!�#��~=��ʴ%��;߮��a�!O�#PVjXQ����\}fe�8�J�XY���>Gh^~�BNJ��>)L������RV)�f�.����䐒;`��0�����_�������?���>�r�-х�e���n����-X��ǝ��z��O�\v��s�򤜪���+�/�a��� �V3����t>�i'�S���E������̚�޹ѫ(̬�]|a6�^X:��Gz䑇���GYlк�J�
YەG��E^�>��.d΃�?��?��d���9���}>��]�J��n���/R6���t��?���s�s�;'�z��Q��{K�k/�[���f\�x|���I����0�UJ��{T�|e7G����\p�4�^����Rz�!�|�FE��I>�ē��oJ즛n�n���{\K����t��{4�C9����Bb�W���E3��r��t��d����sO��!�E��<�`�Nw=Z�{�x:^��,��}4Sw65m9*ɑgPk��J8��2K�7�����_�R���B�30�c)vX�so����l�8`��:�0]Ca����z�m4�.ϲn�,�QO!bs��fpe��;"�$�n	��~������L�4ͥ�lU���&��Y����W�Wc�1p�4z
��7���#p7Z���i�c]gk��X�%�xd���L�O�O�%̥)��t(ʔay~�}�����n���Z�o��Y�׻�<g�%���JQ�^�	��װN��3Z�3Nxc@����H[��H/@Ս���O�C�eM�ߔ]|L *O�Wn#Y������/�l��;h?�o-���qyC�,��6��{i7=@ߏ��:m;l���sғ>�SFt�d"���P:��S�.�l@#iwyJ�U���r��$�Q��w�����8	����ϫ�J�̶��R�x���f����,+����X�o]���?�¿�Y����^\aԋ����I6���۬v�ŗր���K����U�X��P�ԇ�oz��盎z��WK�8>��r��%?Y�7�,�rƭr >Л��<� ��i���i�����۽��W_����5Md��z��E{{��S.�O������:��d,;���q�9�k�i_�3{YHb1��~m%t���`]�Uؕ��; a���uu�\���߾3�ֿ����<p�\��pue�]�5+�	k�������Ւ;�-O<��<�(�䎾L���	g��z��lh�LP�c�p{Z��L��dkG_tqև�(���@�;E��>�_,�য়���_���������K"X�Y|�U��L�[+m�W���,�.�z��A�o�j�):��,]@$���xnx��kv����_���������nxlW|;��{�EO�����{|�t�M���͓s5@*Q]���::ġ���"���}:�;��	��ǆ>�M��,�@Dv�o���a�Ȋ~�9g��9!�o��V�k�0@'e:r}�5��|���������h0�_�@x�pT	�Ű�2:?��oH�)��3�ʴ��洅����O�ӌb��H�y��Q�OFB�˱V �����T���0�M��Aq�Kو�9��j�K�8:��R�!딳n�F���t*�
��˚����w:�n��]vEF�/eM����뤭~��i]�f��eWN����iZw]����k�ft���Dʫ�Fϔ�&��]�Ų�KZ�=��h��}wTv�<<V��4 0��)��\�d�+�Pbr���g�|ݩ��¡K������m�<�4��5~<�9P^��ke7�f|�d;��c(c9?8���i��ʚ�szs:s�����8h�Z?	�) ڨ0K�5]�������(��7�5`㋎���OXJ�=�Ϭf����O�v"���,qQ�����W�/]n��=�OY�=7��M�oR��olBCs2	?K��V�1赀����S��R����i��n�f��b3xe���
=�Q�����Rv�/�mTv)���h`p���MP�L�~�S����3S����L+����hx���,ya-�+������.����*�xk܊ϫc~�g��_xaz���grX}�l�p���>������<�R.�ܵ˵���e��j�<��7x6�m�pyT�wf%��([��ߣ��m.��9�N����5X�}̦Z͘���b7ڃ𖝡!��W���1�?b]^*��Qh=S���P�(�����J�F��Qa���>a</��iw�,h�W�y7����U����e�|�����w�t��)��	��>PJ߭��P�O�Yy�]���aџ�M�EKg��#K���}��R�|Ђ5���9N���?���g�����ͣYC�S�"�W�C6�;�H}��}[�A�zǀ��=��#�m(����E҉�`���e'�JN7͊��H�E���Vwm�dP��q��w��!���%�m���5سx��� �,��C�_+TO����x��3����=���]r�n�^ؖ��*L ܺ/��e���ɥ�ҥ,�أd�.�]���(��R6¹7�}�9�1���=�ޓ����m�ڷ����̧sn�F�jI*l����F�Q�ѝ�c��}���rpv`�I52��������0�Fћ��J� ��I~�)ZDo��n$UN����K(���o��о��b_#�s�4 τ�/�]p~ũ�DP�~�mYϬ�����|K U>��Y�\A�4S�äS*��ܭ�ÊVc����b��zcB��Su��[f����5 !�5(���(vR�o������Fٵ3��K_Jͺ� keW�%́p�>� ,�N������VT�N�X+D�X��l������Q*�C2��M���5�!ߔGF.u��������h[��?+.�f���ӂ�:���ɚù}�k���gW�i���˥n*9i����t);��Ӭ!�T審��]�ՖݏD�0��!B��zC'�N�u�;�Nؽ6��J;4�멧gZ(�{<W
m��U��F����9�[	�^k*��[Ҩ�6C�ۊ.a�������%/�k���vy�x.�Y���ܹ��x��i���{d@����O&��ձYB��f�|����xYbXp�^4!��(�x,W"[ٽ$ʮz�>�C,N�	���c�Rn��t�~Y�w�	�=k׾��u���Y<P��B��(KJY8����ب�2Pں�n�S�)�Pv}`�wY���,��Z�GM;:�s*�C�[,��7'Vиu]�	��Y�l�_���v�����k�����V����s���KC�\�Ekmq_<'�(�����GO{͸�S�ߕW]�<scj\��'|┵ ᅫ8�wq��ޥU���}����������R��r,��޺��"��ϫ������w�����rx��93���Ȧ�x�����zۭ9^�?�At���}��~X���]�-oˤ鸸| ���7���������dN���/�r<^����;��Ս�0�����"|l��ң(��,�l~��������/~~�t}��7�xC�����j�� ���-�o�z�_�7��Q���������KYW?���6�!z�e�����c�?���;�n����O��S)~u�M������l����C�םA�e0^�uXv��,�Qv�8�x��TĴ���[��t��D	�"���AT�O 
���E�3A�G	Z�`�t!��~��_�B�O>)S3�|�'[�����ɧ�4�y�!0���I���qp�F���]XJ�?���x:��S�h�c8J��4�?�
��cO����C\`l:Y��nAI��1�<3BPZ�i-�C���eJ������_k�ugғ?Ǭ�W�Q�Yޭ�ѹ��,�y ������)Z�����J�"j��	iP����?fC���)m���햀F����,Xw��c?��"D��������M����Q�)&�(=b�����g�QV	�G}��������Ϧ���uM�Vx��0�%�L<x G�T��B��Fi���,�Vώ�/~�%��ͺ�����>c��2�FÆ����h��<�N��Z>�9�ݶ�߀R6��ｎG����9�UbI?n��o�l�iIS[\�$ɤ�!�%�����@�@e��	_��V���K��˪�w��߭z~k�����W���#�R�5��s�gN�����3�;��t�v>P|����]ɈU%ϠL�i�����9�����78�P�Ƕ֦���뺮�1P'���7W<֯��g�p���'�(��YJ񖰕]Y�`����p&<X�Z�	7���
ci��r��׾���{��ݿ�w9_<����wق�
�7�K�ճ������#VT���T���Az�*��>�����|f���>�n�ĵ�~{������1�łw�I'N�����/_���{%��א���������k�L�J��Nɺ���
@{�:�R���?xڳ�ܳ���OQx����S���݅�E����=�� �hei�Y3`�ܳO?5=Vtx��W��oU?�Vӿxĩ5���5Yʰ��O�ãr�K��Zؘ��;~E;tQ�>Y{O)U�>�|�W.맯ж���[nK?ú�'ނ7<S�]=���܂@�����i����x@bῙ�:X�h7���$�q�:��GE��&\]GRs��U��=(�>��+l�ċ��ʊ�AY5`y�h��K��<GY�i����Z��"{�1=�"� #�F	��i�«/�>�7�$���i�M73�W��RgC��ɒ�I��m�+rfȫ�͢ߜ���Ͻ6B���K	�%m����>f¨C�2?l ��֛�^{���{1L������@�A$xTy����\����8像uD�a�P�fc�@V��6��|)�A냫����4l$��������,�R�|�2���)eꩬ3���5���8_����5
1&D�#x=�=�����N;e:�F�F�,F>>!�ff��Y5��鱪",�J�98D��� �JKl���;3z�T@Μ�0�G��yo�R�Bb���mm=-\��R+>�s�M����~&��8��,��Ga�jTFX��XDlj#�ЦG߽��T�Y����j�z���|�B����!�F�,����h�4��2�G�����Y��
����mz��[odc�/�(�u1����P0�qC�DZ(.��6Ӧ�f�zk���u���r�
�5%�tb���.�
�a;ߴ�)Ug�i�4H�&��+�г����c��?0_	��xՕ��Ӯ�#�0��Z�G��1�.�+�4��S�9�͖��^���Í4�f!�Svn���ͨ^gd`��i� �P�N��嵢;�@��~��#3��\�}�u[�Ս)1r��o�t፞�3�^��5�ʗK�G�uڣ3��!��F>��iϾx�N����]9�n��s��h�$��:��P�n����Q���d�8��yj{f��:����jۦv�M�� �k�eY�@9t�:1
�c���^���Y%Ӣ:ikjYm�wʶ�J2��qr��*��VW@)5{P��L�L����҃b���  ��IDAT�uqJUu�X���d?����X�B��Vp��ζ:p47@JBU�*_�&�����:�{,PG}T�)S�ｿ��RE/��e���>�R�@�j�=?���{���R��\b�y��Ϡ����lN�x�a�W��RO�ו�J_f� %ml�r����+b��q� ��8�׽4:�c���޲"ٷ}<�s�[�����Ц�gP t��#�k�羟��rl�F9��+�p�Wt0�ˠ�}CZpK?���6%��VW�]K����2��U�I�_H���u���|+q^~����i/�?����/�m�+�����y�����-�-/���y�a�]��i��/K���ǵn��wyR���>ǒ���>���)������/Ʀ��!Ǎm�jʘfY�"�2SY�\��r�ʥ�*�؉���򗗙�����Yg�5Yz�G�E�BL�Q�H�%v.(%,kW�����vf ����>��O~��|wg�Bj�.˧�����W�\)��u��J�°����j����zQ
����j#֡�Zex3��������G�n%�Џ\,'���Pu���4ni� ��!�h0p��f����O8.B�2x��rC�"ܽ��We��py��C��`mu���������܀5�/��/��~�/��
��_{�(�&��FoEi]K�/e����������nӓ�O� #@ܿB���9�Ȣ�u@6X7e��^%x_~���*�/�=��9��g]��s�{��sף{
M�g�Tď��(���OC�.���/�֎��OV>�ʹ_=�����y�=�a�w�o�3�6�b����i����K�ӈ�,���Zi� �S�*� ~��+�L�V�I(W �ԀS������J�ӔG��k�4�y��^%\��ZVy�O�a���]���Z�&6�Ј�A�ʳ�c�*bǗy9���$�
�#��r��f���-�28
��cW��q����_8Ϯ@��S2@h��S8�"������7�_��D�#��i
����x��f�{faЛQ���y�K����Y�ޘ�,%˷������~��~�L��=X�p�����^śE�9-�C���߯�dGu���qUn��j�D�2��*���k%c
7u ��N�ݐ~�����u+�V�����^���|Ԡ���d먣���\K﮸���/�.����B���Jn�����|/�\dC)(；)Y��Ok���|�g$�/�K�׾����&�J���{�����<\o��ק���躈rPn�ݪN>�d�{��Y��W�m._�Sm����7�몍�Ksо���W
n{ڳʄ��Xsu�������#��!��'�Π�T��'�nO�h�>Jt)��m������Q��Z�̼��s��^U��T[d���.���R���c8�F��󛗥�*-c��Փz�0괈g6�9�ְZ
�x;)�8Ǫ�7��׾����h��L\����� �/���;��>��랕�2�B�$|���/�B~q\�Я�}�y~Q0��].cP�7�|[)>�L������#GX���Tg%2:�A�P$n#dJ�**ӓ���>�.C[���a�$�2`��R0+(an��I'�T��Wߣ�����b�_|>�ð���pI�q�L���ҵL��ݴ���&�N�bskW���QLyι��:2�cu���Ո����iP���bd�q�dxe�~Z<�{�����fM�qm����aU7j�D�#k��� 	Z�6����R�'�7Mb�!m�7 x��N鷄D烮�6��6�B�=�n\��p_��~����%M���av^V�*�o��3����/}��w��'��[_��q5Hۧ�Zyk� P�~�;������O�(+����,�@7VQ��<�ߜoҮ�Gu���9���
�A*�tōe`��/ϸQ�
�����I�w�Ԍi���<+�,�����?d�)����DW`J���0�������})H:�,�h�_�X%�mTy��ݹ�E�@���ޤ��6�_��0�����a��5�������P,��䠧��M �:N�'H}�u�{���?C�������~)B��k��*����VJј�-
Dy�9K��u�pr����ʫ��������,��^�~���;� �@ɠ���SN9%�u�g�)��4X*��?���>��i�ʣ��R�cъ��d�{�2���vuO�R�w*�{��{O�Tr� �28�|/�"j�]_���%sܫm��ے��}�� ��ӱ]�T�+'K���
V4��{~����=r�;o�l�{�������gߪ3�e@"�,i�B����Z9Cǜ0xί��S��R����w�3������iN��A���|(��Pn�3"��m����T����Dԋ�ݔ���F��5T�3ޝe�~ ���ƿ��R�<�i��"����@����2f�.�p����i�:�JZ�r��o�g�x�? a�Q�͡;�Q7��F��}A�z�>���:��y����݈3�k���EI�/^xǕ��
��E[�\9�ЬK�2�O_=��o��t�Yg֠�D���1XO=�l���Hd}��r%���Ͱig�p�L�XدaJ׮A
(E�y?֚���PFӑ�@}?��(�޳��0��t���?J4e�(�4�RQ'�q�k�F%h��e��ɏiS��'�Z�fW��(4v���k��N�>��y���ɇ�׋����f��y��r�Fp��mr�1��L	 G[�j&i����~����4-��Y�7Jlݳ`����E��P�z��`}��)u9��w|� )�6���l�k�!�V������k@J4��W�����X�8x�!늭���G��=Jf�U�:�A��F}�0�fм���z�ͭ�s�6��zT|S��o��*!�y���0� �t3�.�ळ!\9�e��*���(
I@IW�F��V��;��#�������L������6B��9�6(��u�B ;���}�a�]#8��x�|��e�\E���%��=X�����_��Q>\�ſAu�rd@╿�?K�{�\GZ�52�6�< n+H�r�p:F���k�j�`Po����Lg�.ZnS��y3��o����,������>˰v|b��3άN���k�˽l:cqd!3;e��OԿ����B���I��30I}���*>��k=��0��'�߭��/�8vl�R��w+�Ś�_�)�t�{x89�,�#�`�Ƿ q�y�����
����Իwp�j�32x&H'�gR͝x�E����k���m�,X�����d�w�5=�أ�Go�L�p_i���x@9�j�}�<a ���>��0��۔f���#n�q�ez���x�����y�[���mx��@��yح�Y���kCy����V;:<f\x�gx�LZ���G1W�ͥ���%^���ܾ�=����q뚭gF�w�:�y�Z�j�}�K���ؠ�x˕�y�P	J4nn@Ι���;��i[�C}��!��OD�����No�9�I#��ܹ�wL��R�9!�)�(��<��m�x����V���fEou��<5�m��Q��'0�᳘O�"Z
:GQ��b�e0}�V�ްd�2�3|^�G_)��_J�RE��ܱU�	����p��;�S�*j�\��t�pa*}�2�7ʈFp��8:ay�Z�u	r�s��{y��Y���QS�թ�Â.������_�࿺���kvs�ȕ�:l���8�<Z�"��u��ʉ�ch4�ǁN��-�^E�(�w�	:^7�ư�Ƶ���6<��;��V�y���GY�%p�-;ǥK��w�R�(f�S.�S'�Ca�ͽ�"n�������O�h+�>X��+�zS>F��[�#��;�]�F������e�XW#_3Y�U�䇁Qӹ|���|�+eT�A+u��%-�Yq)ڨMm�]���� Z��n%_�,ˊȽȍR0)S֊��H�ճ�5����D	���v���,�����?��[>~��s �u�6�R�{J��c,�:�����<��6ʒ_]���bSp�f��φDhW0s��z���%ȷ��ۣ\�\R����Ͳ�||�W�WJ�٠�����B!�8�qMڕ�\�.d��K�֨ 0zdv2|b I�i�-�ԇ:��K�<�\��|��d�;o�U���]���Kׅ�>�2���q^�M�0�<0�y/Q�/�:��v�k7���W���n�з��p�A�P|g�%��^n�Ύ��g�Ȱ�G�Ϛ6���v�0h�q��dMdg�Wo�}�X;a�u;X�/�gܐ�%#�#a�bK�h|�U�YcX��#8���a���,qt�D�L��A�F�L[A#�o4�T�\��T歷�݌�60Y������꒎i�����>aj���_�u�Ң��L(�Yd�ҋӶR��;\+=�߻�׌�J��n�t	BPg�
p/�7��7`�3"4)��誌p65���5�cG���x6�4��g9|t��VWS��r���N��CnXu��}X@+�٫p�F�9m|eZ�3��8����3���ih���t*�����|u3�=���I�n�Ͱ���,��$��Q�]:P��o��ĪX8�M��qJ�~���]��If���3
3�ȣa �)����z��FXן��N��a+'N�ߨ���wí���F@Cy+����A������Y+�=Awmi?@|>3n��h�i��!W�nwL�ۥtU;��]�@�_�5N�K��.�-uWE�k�����)ŵ������1�7ke�ς;��᝭ɢ�Ba�k�`�-_e���-!�v/��m��9Gw�������r��_��{g�:7����W$(�B��5y~=�t���fP��K�3S�>F=�e���_�>,h�QtK�d�v���X���o+�9̂�kk��U!O�q�4�4����!��v�>�#{ό�}��`V1��m5pq<�����w��ve�X�W��4��Za�u]C���5�?';/gd�V����Yd���~�Q�����]-'ڑUѹ�]�~�!�q�g�"mC�Y����k�� B�Y��ݗJP�rg�|w���:ɭI0��v�WOAD�R&��`:#�1�7::�V�#p�����ci��y����g�Z���H�b�C�����8��U�K��읣�R�J�}R!�+<�$�Ĭ�LU8�!_�2�%ӈQi�>�v6��S߷n2C�i'�t@_��n��C_C�2���|�gi�͈�;�#,%s���d��P�@�\��p`������7�/�P( K���S��~�|����p���p]�u���G���?m�����f�4?���Q�.<F���� ���>�O�E�5E�ـ�nu�9�'���C%�%Jd:�0i%^�ڤ�����������f�����]�S��3��vǶح�S|��߮��_yeV�9��t;^�/���Ǡ��V��pu�{����14�ki��� ����;�u��UD��>�@7�h($K��AB�v%��K^�o���w�i�,���٧p�R�\m�fOysC��at������C�708���g)������XG�nyQC��o�_h�k��Ä���m)����cݲ3�8u.�S�z�t뭷L��vK��]�-m2#f6��AyU���gC�)�����f<��}|�k���{Ma��k�iO�c�t��Ӣ��0�6i���@��6,��0?��ó^��&#lӪ�P��A���ź_�>��=���MUE����I'�t܅����+�N����n���#?ܴ�G8�p���CFΖ/쒎rKZ]�4 s֩����˧O|�u�4���cI�s�?��O�S���'�}����#�<�ʺ{)�/���*�k���&�γf�:��Z��]9^}�����P�D��P�������.����������K��`�zܬ�ڜ�V�AﷂF�9�]�Υ��M��|״	�:��_�
X����ל:���K]������1�өK��� iE~������Wϫ�/���)g�v�
*~�u�!��_T���V_~�I'�3���w=H&Q����z=lxSAv�Pa����P�%�e��K�$Nɐ&p7�q�E28l@��bÍ��CBD
>Ү�y/�\u,�xÁ2���2k��ٝN+��I'V��S">Ry�Vy٨ò7y�\
��{���0������
�8����֘0L�1�(���x��*+�8�P���x�{ĲTb(C�m׊��ך2�9��_e�nN��I�����5ݱ�Bܔ�_� ��3���b�p�CWP� �p�*iZ���2W88ܔU;XA��k�P��%���X :.f���]��Q��u?�"R�%1\{��S#��	�wA��.����bE��h���Wޫ��E���\E�y-�᪼EW��("��LwM��G��Q"ݕ��<Ǐ@Y�ۘ�����U%D�|��k����&���3�B&j��T���kK�v�'+�]�dD:�
ksV+Ý��$l,x��[�fnK�J�I}TY��+�3��ߔ��YOm�,�T�QOx`n3�ƻ�� ��&b���ɟ��t�5}�[<����?�k��v���u����	��|-c�����<���ݬ�(Ŝ/H��^�޾�>��{�3m�s�i�}������X{���y�db"t�4]哼F���� �f�Q��g�H�uؤQqu��q��%�u����U��U��%*��o�����K�,E��._�|%u(LN)D�:ɀ��і,5���:����ɩ@�_�A�����˧i}�֩ܯ}������N�g�җ�Z�_������`��~��We��5��t��Z�jP�\�/$�b*^s]��Q�7:i�9'�8�_Q����d_�U��Oio�y8���l׼�a�2�2��l~��8�r�#�0|�#r�s���/�V�cV�c�����:�g���o�90dA��޷i����W�~{%Y_��M[^��n�jd�W��nu����{g�Sx;���ky/R	��tGǞ��g�����P� n-���ac�Q7���AU���L����.L3Cݦ�%���\�!�S���;��_�uX�wC�:�V-iAY���(:��ր�$��II�dGb���,e�����A8���f���������(�K���X�(��S�Y�a��]<=�v�z��~S��;��N.!��O$��We[�*�K�VT��|-��4~��E�����o���
/���ˍ���t�ᇅ>o�I��yF���-:���q�sM���c�J���Pu@H��B6���4��GA켚��d��6��kձ�XHۓ��C97��N&���	Afo����C:,�pywh-�ݜ�{m,�!�q�,	����3=��å��	:�*�Z�;�eQ:!�4�,�;��f5
�V &�/�-�݋�r�B9g�R�XsW2���>��N�r Ǜ|�TExa&^�E�$�K1+Y����-\�/��$v�3`i�/r��_h�N���u���n����S��D��a�i���>z�Y�?���h��>7�u�����ؑ����p9��Urʬ�>����Ο.��|�I��+���e'�X�wP���;p�o__�~c���pN���O�c���ս<p�o���砃�gl�t��{e �Rgh�>!��5�����u�u�mz(�m��4P�p�kqQ�>�&aw������V����e$��_���gP_�����2R��_�QN��@�0�ng�It��M�4:0�5�Nb�D�3�)�(P33.�p醵rX)��7�C���z#G�x���P�Y���M�1g���?_Ul��8��H�.iN~0�#FG~tb�ǻ��x7I�Nh�:Y���}����y���_%��$��:���%��������we�AIO�F��и��N�C�"X��3��ɳ�*_�	��0����7���wQ�C�����V��d�'�P���N�k��d];~t������ۏ�Z��+�ӴR�V���uaN2���2��y���MB]/QdG�UB�{�N�%��ŷ�Z�w^�?'�}��9,|rF�QG��:������ǯdG���\�^N�84rC}Q�ky��~%(��x`�u]�[��s�F� ����ʷ�$x��=���Я���������K���҄#���gxR��*k# W��R��,��p��[1:m�V�q���W���E����!Gq�fK%�cM�:\��5p�x\mp����N�;�ē���z��N<��i�}�^{���/���jիu�6Ľ�*����պ>������\�V�sP��<��S���>v:��cr�'���SN�ݩө���SO����U.���oOi�xYjvܱ��{\]���Nȇ�8�O8q~.<^��c3���
�;5�;�>.4GfF�w�߃�u��v�7�E��;�v��)3��/�W��o�4�!��9��6�v�o�x�>Tԝ��N�����K������Ș�z����V�<T���kWҐ�0Pi�R�s�A�o?<�Z�Yy�93��;q_AW�jVKH�fb���~��c6$��P!̗@�������U�Q��D��X��Ɍ��?:���o�^�i:4�1�mc�A,k�4���*�����)�#�˸�e�~��ӈ�RNg@��w]�x���I��s���$���u�W]F�G�w��u8����u�K��M`�i�����:{̰,Gp,���z�����(����D	���hK���m�f�c]�Q����h�:�A�V��:�5 ���:hÁ�u��u��r��ʿ)�ޒR�F]���U���ڱ^�y�����J!��������2�ʭ�ї��W .�W΢�Pdǉ0d�)|�L��8�X�-x���N���3�N4��w�/@r���S���*=��n<v�a�!�@mY�n<�.y�-�*L�>�]�.%�PJ/<�{��x�Ĩa~Y��c���X�)���%~��U��W)�u�cFm(fqU�={���)�~D�_�R���)K$�I�ur�M�,�������s���p���N{�B_h����^��n(���N�V.G�7�i�Y.u�$_ѻ�%}]���Q/#�����]��n�xj���4�h�l�20?y����,�`���t�����l>
vE���������\�P���Aq�'�5�	��Ϯ��"Wf��5HxT~�b�2���@6�)ր4��\]��V�;�0��S
��p��ow�.��&HqYY�	G��p;��P	�->���G�G'y�Yk2��\�:��&d�7�,N�FĺNZ@
#���=�ψn�����5��[�i�b?����t����tzD+	�����3�[��2L9QF�Rwu��Bz�x�tw�����u~#�u����}���nS��1��0�cz�%X�\4.��ߖPI��v�QӷyE��a(��=/�N�xYg�V�g�1�3趹1���ܠ��x�۸��Т^�!�A���n��Np��tA[��7`�L������2�J[XB���W�e���]FN�Ѧ���~��n
�lY:~K�O�F�r,����A-�V۫}�|0�z����F�\�^��.@z6^�J��^6�Q~7���V��~#��V��E��biVn�<�
b�f廀�Ag����>����K/)�hO�Y�<����;E�Y�>��s���O�ĵ�}�}��|��ǅ�-E׉��v��3�6�ZF�T��~���^#r����_���{�7GSZc,���?���w���[���+\�m|�����?x?��s�=�`�ぼ���@(�q��������ѣ9c��T4��)�c<]9Ǒ.�A�x�
S}�?A�1k��`�]��Ѯv�?���b�7(ڈ��4@4�q��Ah:'�Da)s��Ʋ[����Z�1R�C��+��uq�D�s�A��0|���W�`�M����޽Flt���$�g�����9���q�����i��%x� ז�C�:���$ᕧ��
7U�#���4�5��y�_�oB�
�r�BmN��I6��Sb�+�h�]�_��X��ߢt�z��� )�0+/���'']�aO9�4���{����JOVڳ[2�f�vg]���u�P�z��v��Y�L���v�((6�p#� jѱ�%U٥Y~M�J�{��y��:�Y���$WNX[�cÐ�/<���������p�uq�e��X�G0��.>h��g0�1������I���@64���R�(�zK�)_Cי�8���pv�U]�W�#�v/~��\s�w'�5�����S��%���G�۶�<�����\�%�tF��7��s�t;W�sz�;�ϾX��$�|��r��8��iU��4�%mｬ��/����X���_��>���t���,��כ�Њ�� W�K?�rs�L{ ���uS�>�l�޴B	X�����+�l�}��gJ9����[�4=��ӛom�vߓ��%b٫��*p�q��[ڍl�EB_�x�h�>����Ї���}4��Q�\o���8�!��R�*�|�{]����^[�3�ځ��,���S7��{�XC�z���7ޜ��k�i�=K}w{>�v��S������W���K�ս�{�2���cmӒ�l2�t�Ty6���ʏ�LA�7#EA��ˣd�[��Vh<��:D�� ��(�"��R�����ʤ3�+o�}���2r��|X��.���I�-�#��:N��<�}o��_�_�5@�h?���t����F���.�L}��|���x'��(Wn+~�P}��>��}f~�w�0|7;�e�y�#���%C{�T��Y_=�RoV��}�1i�=����X�l�}<��}�wɯ��O���:�P+��H��������0�F�[��.����L��׃ĩ4Wqg��,�Vpn�$��5k,-�W�+Q���"���	�����{@��F	l�S���*�~=E�v�F؄4O��~�u���㣉w�XN�(�:�J�5
�ȋ�s�jm���^V�T�U{v�'�F%a(���C�M���L=�R���7`Uw~u�����WN�AB*�ͮ���Ho\��{��O�[ӰCk��Π����P�vC�����A
-��ͼ1�$BO�ޔ�(s:��I:�y?�#x�(�W�S���n5P������5Nc9��]�������|u��G݋��6�r���w�@�tL�T���0G���/�:.H��A���
������0����.�;:�V|��g2ގ���O��ݡ�R�U>�:��0�gt����u#����u��£�	�]xz��3�&���y.]��/�N�{oI�c�?:�y���7�4�vۭ��:�;�V90�kY3�[��=��epC�W^h>�*_�d�`;��2ɲ|�R^������KA��z'#m�\ݷ:^kؾ���Ӂ/JJ+�ڸ��ϕ�ɢ���=�oʨ5���ZK4T}��v�/��sr�_�I�E��rF��p�|�tƙgL��qF��w�YgM�\���0����n�4��I�����s�׺>�i"���ř!�w��$��iտ�n'��;��u@�%wu]���XFY���\Nn+�6sm�j9;���F���u^�26�������w�X�U2w�f� �r�J���P�6W�^<��lX<��|Y�W]�����c�����k\�{�n�裏�պi�A+K�E�=�Uk��+h�4���4���b�_[�� �F���;4°Ō#!��i��.�����<��5-]�m�	����3|0�~t��6��^C��&<�Gy��[�Q)V�E��n�q��eh+M1�����υ�fb�����*�h``I�e9�!^�W�efK�^�ec����4��gn<o36y?⻲2�,�J��t�(�_Em�_�ݣ��:��ٙ�\��U��t����z`Е�k�6�q�N?�Ph�b	��9\Fߛ�#�u-`�;V���
o��i����A�\�;�����x��]ݛX�����S���}҇]�)�\���~xՍ�m��2�7�:��t^���l'��_-`�5�T��li����p�F����g�;n�o�P9\��F�:L��!<?㲊[�����&���s)U�>�����[��kY�vK���Mݷ5����0ʷ,��tO���>_f�u�E5���cy	�m}n�3N���ϰu���qe%��1�Qho-��'�Yt��8��)�_\�����"L!�����,��N�.�f�� |y��Jۚe��U�Z�]��7�0�L=����V��?k�����֢ U��>���)姬x�E[��˹�_��צo|��׿���_��t�G?Z9�>8��&�J��I�da�ũ;�oX��a}�|^�ϼ�u�v��ώ?�������m��*�r�������7_�
F~���^]��ܜ^�6�*���Mx/u��9��æ��=6�lD�(��s�ѫ�y��u�uЁ}Z�� �B;Z�A�/7�v���q��Yţ+��N;m:眳�ڟwf����t�y�峼><�9��g��?��|F^��!�X��"�!�g&?Vx/��'{�7h����]~TRO��y��k����P	ky*���"��s�dC�~�T�}7L��� ��	�Nc�ۊՈ���� ��n��+�N��I�E�p����ۺ�2(���"�$^b������"�hh��V0�ƿ�/�lldy��{����FC��v��#�<��U�WE�����H��\@y6������7�ÿ�ji�׽���s&~����X(gG����f<�k�I�|E��q�����C��M'_CӨ��Vx��7��2p#��4�����r�?_7@=��61����K�u:�v��+'��S�:p:��skDxɈ����'�qo�8m9r����R���I�q�Y�H�z���;n��o����q?:��D�b��'^���]��7\�My#���y�,���/q}?f����Qg��l
G�������U����_J֌~e�n��8����y�;�u֙�*��[��}xڳ��RN �yKXw��w�2̺]y�5�-X��&��#�R���5�>ON���xC�0d8\��w�BT׵��Zn恖�+"�:J���~����h����C�:���m��疜��_^:gGxU�JP�f�k�3�mΰ��C�٫��=V�3BF��S�?��O���G�����`{��%�N.�A���߭���/[�k�����������6��*��yr�Aӡ������J9����SO9�����to���'��S�ps�f]����(���
)ﲾ�SoUWå�(��s��������il���,ޮ�ﶺ����Q~e�r�e; �[>0�t[�(��K.�d��������ӧ?���S��T>�q�Wş��+��.�<
�W}"�zGʽ�V�+�0ꄨp�݌o ��+�+������ϥ�^:]p�Qt��U
-��_r�t�e�O]tQ���Rp/�蒜�q�qǇo-_PF|��oe�&��8��Jֽ����>5 ���]<\|�z��Vv�~fz��Rv_z9#�_x1�G� �r:og��������-��O�k��A6��e~�d�k��+zt���
3b�fʀ�G�E��	�
�e(a^�ݬw��`0�֝`����&W�"��W�y7���[�k���@���w�_�}����6������
7���}_����N4(f�rVn�;�k���/i����Gy�t:�qb�4\
F�ݳΞ�&^��Vv�GXۅ�<�M�U8�q���]��
7�K�z�Vv�lk�]�����i�ӛ����6�s����4�|Z��0�Zю�a@'[<���/%���2]x�������?���r`I�x+��2����.�C*�9g����M���Vv��mP9��H��	���_�qN�N3/�gӫ|ʟr�:���в�9:��t�YG3x��@+�#�r��m�!̫�lJ�_ҟ����W\i��^��Y��ί��曦Gy���=iVi*��N$1��dw�E ��
��W�����i
y3��2�����]Y�N:���_/ڸ��##+p�d�Ī�ʛ�q���;�|��粡��W�C��!�ZJ��!ڄ���ъ<}�1Y��٘v <7����'��ۏdM�%��z��_���Rv�v��l�eQ�d��QLP����#",p��1�����R6<[���Y�Yk�Y������ �7YeY�<�/"���w8�K;#;�[�K��tb5ة�����y��q�7t�<���6��}�Z&Ksc[#�*��0���q|X���:������_���x���Pg;f��||��OE����Sڪ����N:y:�u|\�8u}�	Ӊ�n����-e��|��d�tY�3�W���9P�d�ٶ�N=-��K/�4V\�������j�o��C=$G�Q��s%��fvr,�G�0�f(�Z��g��a �xF)�����%#�/>6�ӟ���������Ү�]B��g�˱$v��1�C�pO�'Ļ�ܙ�P�u�w˧u��0u~0ȺW��IE�;�w	� Wԍ�;��;�k�.�k�����?k@4L�uC\A��d	]���DAY�Y�*��a��h�d؉�YθyF<e��`�Ì7���x߼λ���Ő�Fؑ.$�-�|���{�3M;��3~�c-Z�0#�.hX~�G�����z��Ě5�]��S�����#K�6�K%(Wa�,�=`�/�HK����Z��w�YA�gG�l�K�5�|�I�s�
�]ǔ:��K�p��h/�f�bwhY�^y�弳�'E���(?�ɏ2�I�J�U?Zsg[�v��� ˙Y#� �k<�N^j,>�Y�2Q����5���U��~�xt:�Y�˺�z�y$L��0��\�:�e=�y���ֱWB�pI=��@9�Yd�	�3�!���|ڨr�y�Ǣ���oL�����Rv�0bKoX�R��L]g�4���W2�re��4z�M����BQ�-k�>XO;������T2�N���c�H>��\����
d�Y��嗧��O��1��gl+���L���a�r꩙ҵ�s[6@=Ƌ[�qjz0��-�����!�k���t���Ĩ���B)�FYv)����[���u�Y?YJ��'�4�q��Yg�5�{�ٱ�w�y�sF��N8>���s���Ë�|b��f�|G�=��Y��ӟ�$�x�]_ϻ��ՠ���^K9�� e�kX���+^W��RuYWtt]���u�k:�Ѿ��:Y��u�f��#�����o˰��n�M��c��<`��Q4)j_|�t�UW���#�82��X��d�k��>�XZ�Ͼ�$L=r�!�a����̰���Zr��ȳ��s)̂Ӂ���p��W\>]~�Y���f(�_�%�H���[��X۫l�祗^Iy��'|YZ��l}�ؘ���uE�AK�!�x.��5�[�AK8Xn���������� ��W^�`e��jtϗ3E�ԓOF0`i?a���0�k��c�G�+��a��ˎ�* "��ub��#Y���{q<z��t����<-�t�K�N:�pƨ#�w�
�kE��방��<$_S�ݙt:,s��P��
��3j�&�u��� U��±���V��W��ϑ:�쟇A���|޳�po�L#%�#n?/q��M�b�.�5�J�%̪�;�(K�܆�#�r��uոC��9�q��ӑG��9��t6�˩�X�1N�H��O�=�-���F~\��t�^~ ϼ�o�E+���
i�K���U�6��u���[����LViw�>�R�>� O��ow'?��|[��?g�^���r������Wiw ���<�c��w�m����٫ڬ��Y�V8��`@������~ͳ�vP�ϬֵdL��w�t�w�=��r�O��:M�V)ㄯp�è{�4͛�-�t�h��^R̙*�{8�p�<��	���O/��R��-�����~����O���k��t����!�<����o�:���:�v�Y�@:���3��ӓ�_ߑ#}�f9�(��N޺�S�s�9~(�@��U��EzP
��k��vf	�su�Z���c�>�O���Y���˽W����c�?�T��s�r_��<�m%��T�u�+�Ǐ$�W_}%��?���� �=�{C\����^ʮ)c��8��"i�A�-�r���Yg�>�{�q<�����;/mɚ�G}(�������~��K	~!�{��|���К>*f8,���[o�~y�Ӄ��%�>�6Y�[��!� �O�H�){]��R�<�Y�����J]��+jѤ���ꠍ4F����H���4ǻ��a�w�w�K�x%�F�_����C�G3VR�ۏ}��ӧ>u�t�E��٣C> ���S�N��NFL콗�$���Q<Y��)��o�r�2�����+���g߽cx��p~뭮�s�Ǿ��/M��ǧ�֠�AB;����mI~x�]՗� E���n����W_�x{g�.��s���G��%E�;4�St��"�� ���-�唿x`�s���M�$�e�`�셾����J�}��2��x5��jd�0R:	Y�����l���` �+%���tX>Jq�Q8���R.EW8��DD�e���@� :�:�Ϋ�Tә��w��TU�F$\�6X/u�'e���ϱ�Qu�ѽ#���P`ʷNDGn�Ŭ/�eCX����e]�L�ZmX8+q�����e~���!�G��2��T��_w>���!�G�A��h(�9���N�!e�ru�:��NJ�v��i���`r����3���A�I��
��SX�ʸt���aZ;d�w�I'�8�ǫ��*VC�oU:�c��/�wS�(4�'�~o`ԃ�������B2k�	��VJf�T~�ָ�aNw3^\�X���k+_�q�k�*�E9��*�� ����6 =@¿
\�0,?�|+��q�g>�LQ�d�����,}D�2j�諎R/~s� ��?���SO;��;=d be�V�� >�c�^����ޫ'~����#~+��;賦�H��A��~U^ts�{�������N�bZ�㬩�p�����ZSB�@]8��};S��/�u�v=����ؔt�wLO�ӃVҮ��,�������ܞ����uv��-<5����6 !�ߠgfR�N=�����d,Y��:�B�¾�8%
*��O�w~�n˙�<�_����.��6J������%�/�����+����r,���(�_d&G�ֵe(�3������p�}�Wѧ��
C���[���sz���U��������K���zJ�ᐃ�
���r�j��(��B�D�u�,~�_��/��}�Y�ǝ�)t�C��,�,ű�qzQo�����|PD�ԥ�Y��]޹�,u0x-�`���~'��Ά�D�Įtc��7#���F�wzk�z�]�a����y�U^�[|���q�������a�f/���(�g�qf�
��V���!G��{�5��#�">�׫��e/���5ۅM�kK]D:�3�W�f4���/�b���WW��N:��j{�}d ��ӣ�<R�[�����`�ʒ��9�,�6v�YrJ[��>��~v��e�a8�u�䬙rX�t�D��3~��zV^�K_ې�5��^�������"���>�+B��;�+s��eH^��lf�nW�0�S�|���V&5F:�D�9��X�nDqL�"��5�2:N��4� 84 !=;�����K�+��"S��t�Ι��>�u)�L��#~�<"�%LM��Fj�Z4,qB��b�#H��V�7�e�vUW�;�����_dС��Pt���=���),����@j�"�(�+�W�>W�(��j�Ae��fp�:I8)��$7�P�Y�L�X��Rc�b�?��)���'���t�G�k�(O� E�-������9���(P��F�k�%�\;�Z�o�Zq�pK܇_[;|�T���V�ZIsߊW+��k��Rg��e�]�����?�Q:Qeŏ�*���@�v�Vi�,F��6}�*�����X��"ZiFWq�^},���2*S��v�{�2��¡Q��s�߇��| �צ/7�3�W�������U�(Xb��(��b�(�(�uͻRz]ci��\/�H"�%�X5�}�ٜek�]�U[rlY���{�}W�=.Ñ�y�_8hc�Mj��q�v�2k�)'��7��ԧc�da*d*��P(�ՉW"�}	s����ΰWo���2Bȣ�Q�E�R����w�M���s�x�B�O�g�'o�]w�2�_�R�ɪ�Qvg�T:�#����+/G�0�j�Y]�w��R��M�1(��PDXj�yhYI{�O��\�x��@��r�����s��O��ԧ���҇�N:!}ա����瀏?��,��VX�9��I�M���������pCOp��n�����%�~�ï�W,Ui������C�v��k�Yѻ`܏��n�0�G%M��ֽ~�	4چzċg�yF�.�.���XW�8�\}��O?3=��#�ǃ=E׺n�"�@���;zZ�X<��$�Yt~,gP�x��ki*���`|���}.��O�hKx�2����7�S��������S?�'�ƽ���\�u���1�~��l�Xe��~�´�����r�_���L��S|��ڏ����� ��7^�`e��瞏3��A�;L-�d�+��w���(��?P��(**��>�Hv@]t�t�%��a
�� F��s~o��6��P�fser�	�8�4"�E��z�5�L����q�GO��o�?ᄓ���i��B�c�9.�Q(��}��(�'�tb���^�B�%�2�U������84�e��.K5*=n(����B�u���y7\��?J�����NZ�%����:�m}�4��_ҋ�(�AX�
�n��J�\7��C0nt�А4h�z��ru0���� 8�f7�i6���ϝ���0;�.�xx�t��%/24](��*�v� �kX������� �L��ܱ���Z�.��Q�9[|s��kr	c
���:PN��kA�NƱ˘���R�ԓY��{&�|�`�]����vP;��ţ�oh+�\��ڊV\	�V�\���V��}�����~ܺ��FS�]�a�,�����	�k�#��!Qiq��E�BcNn���@��r�n)��r��Bn��Oiឬ����3O���	���<eA�t�����[�7��%_K��,����"ƈ�p �{~)��L_���"?u���({�cкgN9��d�S%��UO#�����Z����Loc����g��<��SWO_��צK�Oq���iʂ��k��,[S��)���WO	�NG�'Z��?Z�Ⱥ���Y��K/FYP���t퀿���3�L���,�������e?դ��L��*�M7�g	�����̧��|�+Շ\��ɀ���ig��c�=6�WJ+�:Bo�7<[8�n�(R��?�f�?W8�39���7�KMW)p��3ܘN���o�xn�(W/7�_>L��¬d^��� �,����%f��j\p��I����� B��O~:��G?�~�ӟf-��=8=��3�^��tW)���r�t�7N��w_��:$�c|��A{�����Q�� =]2ᩧ�>P�����z�aQ��X�T���+]_�������.eU��K���j6C�3 <G.ث`��e/�33����D��s'�0:&��zn~��к�i_y���?�]�{:�y�^�:B�ݭܱ6
 e�{����(�|���~�B�s,�ZF5Z��*���f�T�y'� �Q�KcH#x/���|&~�x�������^�^	�$�1e���@5n�և���
n�`u��'f�ؗ���%#>�aJ�S�b��ݺ<J�<�x�y/<v�}fTt�=w���X���H�a���h��'8��+�n7�'�	-
M۵�a���:���<=%�y�^xJ;�+N���xɽ��l��L]���8{�[��=�"��NF���|��{��V�np.��jtO����8aa4�6�:��u���K�:�>�lݑ�g�z�����W)���6h<ӥ��X�9X`�m�E{	�p+ec�d�r����x�;и�6���3�$41:'��R�������(�:ۍ�>�����f ���`��5��چ�)�ܸ�B	��c��ܮF^��ޣ��ׄ�������~ʽ1dØ� ���a�Vnr�}u�ڀ�K ?�w�E�����Wy�%ˡ3X���E)(��7���u�ٜ|�v��GDek�Pn��OrX�����?�~�7k:�̳�� ����6�v߽��Xv�5��ݶWp�<BG�͐�B�t�l��t�>"���ߎ;���/�N����E��\��m���*�V��/E/x��@�%6����Q<^+���s��3����`���uG�R��R}�����M���1��0J��ⰨY�!'m��,�N_��h�;�^����ߞ>��OM=����,w7��Y�E����r��@Ա��A�K>�u��j@op2@r=�O��'�S�!d�����p��Gc��xn�c6o<�e�W�4��No�}�c���@�5��uo����[|�j6����L��,�%$��\��3ӽ�t��b-�/�N4^���A��U�����N"�zt�2Z�g�wo�ܭ�J_Yj�_�X�_Mt@,�W^���,�w�yW򵏂����?�h�x��lS��Qh�o`�33@�~�p����9�f�}Q������M�g6���?�R�\��4,�!�д�᷽���Z?�n�s��9K����U�?�������O<az��]*��3���w�S�eӮ��9HUr��60I!#����M�8��g�90�׾��,`��c��Ϭ�V>
đ^7�j`�mԫR)��-t������&�!kP���q�Ơ�X������+�HG����5�1�'N�UJ�����u��ݴk���^���o����g�]��+�7�<�(���j�
DA�Y'ؔ�15��M{���g���Y�&b^K�]�TGxx�i�.��ޡ�u��Ns��Pt+L�5N	��\c5�|�����%�s�{� �N��k�Cj��ΗZ��+q����� �+�	��l�q�Z�+�)���M�IhSW��L/�)�����:x��7Qt���3��t����!}��;��g�3�����Et�ݝTu:x`���|�{��*@�c�C]��_?XJɵ�NRtm��s4+��WP�%�<�ܸƪ�w�Wi�WN���e1cq�Ȱ�����.'̀�u�<�~`��TvG����/8�V�|�䑸iӭd�Y�țVvg���� ����t�N��r-���oK�e_��N)�UϬ����~���N�<��ś�0Ȅv�M"�_��.z�w+����|�������g:����Ipf�h`]�����|������X�n��<���g�>}��G·a�N��m����͛���w���h���^��#
�^u�6Y�����?�_��wsb�zH�+_���w��f�Q[e���؟��gӍ7�P��R�=jGpT6~�<�[�[��/~i�����O�2kf���>���n+�]�Q�x��[-�Ꮮ�����ƚ>�I���u�p�	-�)����j�Wr
m��靴�f��'��A�qȳ�E8�𣮰S�5�6�r��v��R��n��%���:,�[������h�(���5����R<N��Z����z˭ӵ߹6���NDP�,��[Ƃ}�ٯd[���y$�<�L�����g�}N)�ϸM�����7Վ<�L�[�Iq�� �����Y���8�c,WQ�{�^���US,�f�͜���0��{�v�x���������_}ﯦ?��޳5�����_��Lo��Hխ<��G��?6i2�ʏ_9�������O:qzᙧv��j w��{�w���`��{����0^�&�q ���E��>K�vg�����/����ǲQ�#��(T�0m��ћ�3�����A781�����T��7�:��G?��������W|�����?���l-�����o��r�Y5�w�鑥iE�h���
��y�o�ʈ˹���s����~7_�q���H��7�U4�u����o:﵇��q�!��	P�FC��\q�OZ���ݘ^ڽ�����KH�:�gם]h�.�|v������r�Ϯ o%���y�u�]�{epD8���Q^eůkʬ@/\���yn��l~UW��XE-��N���Q|D`HO�<k��b��Z��\ZU���r7v�1@]�cnWF�hA>��sy�Π�	�WK��n1�e	Q8i�˺I�-����@܍eQ?�7�]r��~���)�*��;�H�*���5��fyXA�<�,�ʻG�"��⪻�z��:��6��L�--��Z-����Q2l��R<�b��ך�1I�.�N����?י�C�E�a1�z%��_*�A��n�Àd��;rS�e_�v��/��~�a���׿?}�_O��T����R�C�y��G�;n�ez��Gc�����옣#?r��We�½QJ1���8H?UW��dZ�T��6�U������:V&�2�`y}�)�&������9�֩®�h�[aW���׷�׵��������	�T|��_�~�ww��s�T���T�}�����Oӵ�^������W� /'�nI޿���2�w(@�����N���w��������>�#G���j`"n��w�x���V4��MR�Bx�z[l]	b�*Ma��J��t�������inTv;��C�t�f]�<
</߁�1Z�pK�5]�<�yo#:�M����#场p��ǖ��>���Qt��_L�]w�tCd����#��I�Ly�6Ε�Η�������g|c���q�$����h�=��/��H�)��'?�I�]���W_�_��`h�u-MK�@���λ��50c�:���ſ��ج�3B����������@�A���!�3˪"��}f9��Y�����?����z������Ʋ{�=���jT�]����@��FR��
��AJ��6���Sq��# ��YsO>ɗ7���xh��o��:.�o�"�z�kG�!IG#�axg�Hp������������~��������K.�"mrX	�G+yq���dJ�FHH��x�ۯ?-�E�:0�L��n׃�o����Jc�M(�M*-D��5&�ӎLi)7��S�Mo��J��8��>��1E���.�Wc����m���z'�2ŝi�Vv�t��$��1��L��B�0�k����rAh�w��
��:�V�PҬ���|�^�����:�_�
�q��U�� ��&=�ԝ�k���f�c�=f��*�V<"�z|7�N���>R����i���%��.d��`]c��[�6c�_:��Zi7����Ug�q���Y'k]'a%=�jӛ�S~}��~�+w��U�Z.�������v#���;����V ��C�:As�BVx�2�w���7뷦#;bڿ:al�A��2�y��p��:K�4����%>��9����� ��We�ذ(�����,���n�2ͷ��fЩ�fC�Ҷ~�����n'2��#�i(�ەa]���'�4fY2p���m���7��YgW|�Nu���=������N7���鑇�.*�T�@�z�צ�ﾷ���ӥ_�Gթt�k�]�u�g�a-�^�Rvɳ� 7A������Z���7tԀq�&#�������]=B�Z���?���a�9�K�O������t�5��6�G�=����R����of�<@����ar�dӿ�W�*J��GY��������?�O�i��_?2]�oe��
i8P��<g-|d��l�=���<e�6B�β���o�Y�fʁ�t��k`[��<�s��ײ�eC�K�(\�N��_�g���	7�;�n~ql䷌3��y���K%Y_���XK�x����\3O>��t��Gd���G�TYe	W퉌��hSfFn������)����R��#=���5��~�ʪN����f��Wf�_|ᅹ�h��n@`l������ޞ�.��g���ӗ����E��'�zb����_�i?��r�q�`��ˮ��ǡ��E���W|l�G��N��|��³O�z��F�4�g�}>��i�:�f�@���կ�J��f�ԩx½��:%����k��ڎ#:`�cy�ŗ�|��֑8��Q,�*�uM�}�:��4
�-�q�N�!u�����f�K.�d���?��A0����ޗ���rL��;*�<"W��J' ��{�;�c�=.�p��Cq1��YðE��s}1O+�h��MS�HホE�Nf�L)��\�B��O�td�t�_Q00��/�Уvu\�
�����b¾�Z@�.K�8�����Jcy�`x���F���ug�5���
=�|��nҶ��{��Q�(�6T^}��9"�`1E��3m�O81g�����^Kgm]1w҉}5�9��W��-��ΦL4����<�Y����>]�\^��<�:<\9me7�S��^ҽ�M���w��w��GZ�^�ߐ�,|�{*� W9���,��򗿜o��Y�}����,,֩u������_~Gս���0�C��g
L�,�s��j�cǗ{�����ȟ�����x�UE���(�E^K��,;��C�������Lo�t�k��}du����~��v�i��׊?�x�����@_�~���/��Y�ړ�4�A�j�������ӣ�>=��SS_�������cOT�{�x�A�����a��F��\2e�I�:k�2��L���Ø����ZX��ɧ}f�ӹ�D��5�C(1��G�3=���6n��s��|��)#޷��1O���'��L�-AY�ʈi����wz��5Ki�;h��~d±BR`�^�gR��e�����k�}F_���S>���d��x��k=&\o2-�T��[+�CI_�N���Ít�]���߾�n�<�X^۹߭����w��y�Y�7~�V}8����'�,�Iޏ1����A�K�2��v�P�uN1��P4񶶣~#w*�6�o�:�g���,w����c���Xi�E��ߗ��c0t����NxJ0݆�ŦG�k�{t,�{�lZ|D	����'�L��֠!��c��:y�Q��S}�y�٠v���7v��"E��Rx��Ab�8�`D4��l@�#Ի�X(��R���nW�s֡�>da��~��N?����@�usHE���Q�3�
�"��w1��~�Sq��:������d�_(������SO>��	�Ĺ��A�t�sZ:̣"$�ˤN��׺c�Y8�-�V-���vYH^�Eg�5���W���:�1�C�T�'�8�m�����g�$�T�Uk=�[u� C�p�:�؃�o W��<����H���̠����|�b� k��Ӫ0�u+��.u��!A�R�x�XP�2(���K�첚���ӱ������Z�sh�4�����:�6�_������ޔ�YKv�9�>�o��2�zP,���Ő���:��!	D�� נ����e}�f��i?�K��6��1����c��Gm��CY(�d�v�����d��K�-Y�ZT���uڬU�9���F�8��bv�:+��qO+�����l�o���6B�
K�۶����Ι��UޚL��mi�C~��p�g���ƨ۩ �^і{P;��
���#L�{���*�|~s���:�*�
ﾕ�KVʮ>D}�?�uN�I}���g��u��e=�p�j e��mX�s���=��(�� �m���%��%�p���P�,��]
�Y_a������'�.)�2�Eʠ���� k�='�Pv���`�9RPn���(5dͨ����fh�|���+d�!��R�����'V���R�͈�������)�^�a�6�T�����w�o��nKC1N��{���å�:��T�3;	���ִm|�;�X�amv�?�G�o�:��3pe��{��E������N>�(a�\rqɫ>�Ω2BJ��7����-�,{`� ���m
�d������/�X���O'?�(��~H�sLW�On���9�yh3M9B��R�+]}^f��,Σ6�.V�_�;�!zړ�9V�I|���Sq(�6�|]o���7����]p4h7����k6O�7�BW�'�E�C98'�|��c�����B���nú��4��m�m����+a�:��̫����)����D�U�o��RitK���Rg��V�/w���ʶ��F�u(*� ���A��h��2���S��)�Yi�p���﫩<�A%�b�t�L�lcx�F�r���-fp!������&IK�f0�%�+�m��J�J42]�/����4�����Կ$����w{��Ά��� �V���֘��� ��<0p�2ɣ�n�6�X�K��dCI�s��u�M�s�'o��c�o���/�7��7ʩ��ߘm���s4�Q�p-m  m48���M7��AkH�޷-�xEGj)#l�����8Vj����/Y�7���4�o�7�J�s�eàAᦽ���+�4�h�s	7	��'�������������_�vv;��tv�t�!)�?��䇎��Q���  /.����#�.���t�M�g�ptr:�tzu͒��橷ٍ���S��c���)_	;�U�{��2����Rj�/�?u�TB_'�ٲ�+Δ��x�S�E�F٭�r�8���m8��0.��[ʝ��ˆ�=H��Oxi�W2{�e��S�ڃ��ڞ�YQu�>W{�	ǥ�St9ʠzv��v�Y�U֍�f������~����T��2�9mIx@�S2t�x�.���=�%p�w�tk��E��V}^������s����9_�s\����K��t��Q�)1��Ҥģ9 ��%�<��{�tL)f��]��vt�<�v�'�ʀR���� �F[���7h�S��[�ml��b��p��k�D���j�Dɧ,��V��1�u�lEk�t�l'�� �����W��.#������r7�����hl���x����q�t��7d���qͼ�{��<��Z�b b���p�th��S�Nht�h�a���7s�=wO����ӝw�Q�o�X�w�қ�(�h�o�F�^8'5�?�[����W��������Po�VDFV}��g��Ǟz�Ȓ���'u��u���Ŷ�~$��y�;v�������]�|^�P��C�MU�|(-s)3;�
�����{��dQ:���@ۦ�+jM�
�)�?�I���F��_Ӄ*��q:p�zWX��щdAumUasG�Q��F���F&mU��Y��og/]�8y�Z��V���N�2��9��L.�d�!>���6Ǡ�&�B��0��y��"d�6�U��&��ʣ���b�R�s�{�G��5
�pY�7�uM0�꧃���)Pa1U,C�	Ee�r`0�5n�[ ����x���Íx�����a*=�0�\+��
�m�_*-�� |��gy�7
��N,,3�5���oџ|�I�=x��Q&u��pv�B�2^��}{�J�J/B���O���
k�*��%܇3�8����%����54���k`G�*%C{���L0�3h	F]�Z�ҕ�tໄa7�2��m �M��M�\���!��D����K�h�?E�,d�c�3kc��rJ��c�����p�	6ݻCV��� ���n~W
?�.��V[�y��H9<{g�h@�����dvǒ,|[d��:��ë+�R峪�+ J��x��V<F����)O��.c���"|��$;��{Ϟ�DSJ\��X@7�mPʮ�/���͂a��A���q�U���{�;g}�Z���?_@t|�M���x�I�ӡ� MP����O�t�?�� 6�eW�9b���O��/�8=S��Qy�}����3ԯ�L9�
^���I�k�e:J�/~���J�R�F�p�Ϊ/���w�3�|�Mi��־#7�z�R�KY�Y�8�XmZF�;{ X�C�-ҾX�*��՗e��]�o�y=3���DUl��j�$�S�PRf"	���1��ʩ?����Ĕ��n^���̵������o���r-k+.���c�Si�'FiHk����\F0�+��m�+����E]�=A��o}V�.�93�C��ߣ?=�q�U�if)��6X�)�f��?��V�C����ʣ:����v�z���X?��O�9�i���{��,ߤy�A6������D,�<��2b04�:5�X�`}��Qr[�O��3j��mm(곚o��l�2��3���}t���N=�s7����D9����󁯋.�`:��z냖1 n>*Q��R�e�Կ�cT�A�VtݮX-��E΄�����u�)�C9$̠r�U����b���/o�0ar���[�M��F�OW%F�-�g	%|S�vXu:��k���5B��)b0�i� %����Ә�@��z�-9-A��T�5���*�m�T���(�8��9w�]����Y����O����5�F`}��;E��s�)$�@�T%�+�F�TTOc�t�d�z��BuĿ��I��[	�,�
C ���W���rp���:�N:�nXa�Գ� *<]�
:��ȂQEIع�i(��t^GH��'x�Q�f~0��
G���, E���y��:��G�׀O+~=�F�w�1x��S���[��v�����VJ�\�Ѿ��E����ȷ��Cu'�|u��W��o�,���������F�,Exy�}{Ìe4�B���h���'����@����ъA���4� ��Hv����Y��:u_i��}ױ���N9��霪�cګ�U�A&\p��ӑGQ�}�V׾b��Bx$|ҝ�g�-�V�(��G}�Ϭ��e�_ӠhePʺZa�fj����)�}�t���20�ܶmoU�<�j=��Gf�M��rғW�Me�6Q\T�+WqDX�Sr� N\���P�:]��3/�0iOs�����2����*���'l��Y��S��A����3�i[)~/��kC��?����\�B�T�-�͊e
�rd�W�@5EB��ɫڑ�����dˈ��`�e��&]p�Ў��gJ��KۡT0=Y�����%�MW*����|�N��c횑F����s-Gje���{6���j)N���۪�y��mp���d\
�mO:ח<x��~��&?^���2�d��@s��O���K/�?v)�.�˯�����H�+W��P.Gq#���	�X������X�8۾O=�>I(���Zym��� 9�5)&�N��;>��p ��J�e����1��'�^sغ�+�L�z����K/���ԗY���6� w�2�1H0���r_=���d0�Yb)������{�����K�<U<j�b�(�ӟ|P�1��a��M7ߜ���wh�䃁�"k��7}��,�%}N����Y3�tVEK��VX�j��)W�a\r饑�*ĩ*���G[�� q��+���):m(��/`�8�pt*��6 �3��^�uwew�ڥv�hFj	1%W�����g?���h�*S#�@���o�3
���X�tb:r�ȗ�4jFLNq��� 4^l��C>�S$0"��>�@�o�zf~��r��31F��@�Z4x�՗C�I�ux�P��i�MQf_�+��XV�*����eg]kƔ|LQ;�a~�G)-�47��)���@	Q��ڍ=�"�v���}���O^�v�?9��ˁU���0
g�b٩x�?4��ʟk+��\�u�F����<���k�i�
1�[Ó?��{a?lW�������<;�$���Qg�%hS��#���G��#h��M��:�sq���Z�7+��q�Y����]�J�r�F�=m���U�58쁛u�}��z=J����l>�4o�Y]9tǏ{?�Ǯ��Ө�u��B�X�zX��3.U���SN��%��w:G�W�.���*�ٛԾG�2pІ�Ti�?�.O.�R ��N�q�|( �r�y_t\wХ�U[B_��Z��VF͑m��&��4���N��+�x_R�Y�'�����V��k��8e�H�q[޹U�9�{����;a�.*e���%��x�^Z�O/�r:?�y��6��hm��2K(��:͍�n�h��v���zh�v��[:��1��]��賜��<w�w��Ԟ��K�e�D�@��b�_�eF�l�~I�X��8眳sH�M=�綾_����,����!;���t3=\e�T���)��wi��O:��?��q����~p������L��١U���~1�-����(������=`���^�u��T�
���?�9x.a!��aa�0<���cB��lE���%ب�r����ؒK�����j���af��[tT_tK3��ͬ��8��x�W�}-�Gf<_���c����җ@�`9.��K��)����2z #���+4�ْ^��/��,6T_yՕY�b &]�28�{����Zvy��b����m�l��K�&����l�Q7�����gp�ѳ�bi{{UY,ˑ>C�>�C(�����t(�k!2'պF�.�67�3�A0��}���/�pg�=1B���O\�$�PS���U�v�aD��=EL�Fs�>�����qe*�hC�YP�dĄ��S��#�����릛~u���#�Y0&�(0�� X����Plu�	k����a�MQ���>{Wy��,e��-)�'p�b[�ӓ�t�C�4����:��k0�H׻��y������kg��OW����FX �"��!��zZ�� \4B4f��X��^;�3n��q�8
�5�xZ��*�� nH�L�JC=�#�n�H���Sa��U���Su���ŋ�	pQV4������@	�_�ʭ�%���T�>��%X���������\	,<F�վM�luJ:��;;:�۝�r��vnйַCຑ�
�,yھ6i�!!��uT£��
�W}��l�$�L�f���+����뙕+a����H�adP	�{%V/��������݋ˊC��{��W{��
b֩ڸ�K�\�k��:1H��aY)~]٦�4��].��'�Ŭ��Qr%���rw��v�U�t����aV�~�&{��?a���{?��pXv�]Z��8��dm�יs�15�<!Kڎ�w�����|J����j��ޭ��V��:o�����Q^J�Vˢiѓ���g�e���N�N���?��KV~������Ыe{�Q=��0#��Ȧ{�?�ɖ�٨Դ6��)Ew�e��7}B՗�Vy�G�P9*L�Aeϒ�W�/^�8S��*u5��z��ɍ�d�[<��55~K�yg��]��7TЄ�GZ��{��:�~�n\���s� k<���z��2��`X�x�-v,ѻ�e׺ۥ�˨f�,�j�cәM��A�����G~K����O~���h�7^���_Л���l�����Ea����}D�+�G_D����g��l���l��/�xe�)�<]�V\m�r|�e��=��[μ�s�@0K]X��]�ڧ�O}W=�}�|�A�r�2�El�F�\���s%�qH�d	�(�#�:Ù!rYW� 2sܱ�F�5�!��,5�tG�N}�#�}���R�#�8Y�̚Ė�}�[��u�>;�{uhF��Ȏ��\:
Ǜo�Q��Ř��_t&�uQ��7�8�ꗿ�)��",Eה���٦6����-�6�`�Ȣr�.�����D�*���l`�`��Hϔ���F*�������R6�9�c1m+�ݠG�F�a�q���S~@�����Y�@<:ܺcm��
bwjs�'��B�A\i�0�뎊�:�.C:�a'�r#��)��]��i�����g�ơ�Kؘ��A�	�ݏ�vZ:8ǲ�-��F��8 f!���"�g�_�ո�2#R��uU��������>�J`-��_��/��A��Y�l�4h���>��#Qx�Uw�a�:��^b#>�,út�|����*�uZ��%`)B�R��>���W������/��@�mզ��t�E3Imѡ;~���٬D��e:��8AN!b����5���Qůhh��J�{��@�XQ��)�M#k�6��w�~9��`
ݭ�3�~��f�X��_z��M���?����5��5�Zd^w�Sz����\G#��K��Y>̼ �(/�'�,�!*�
*�Ƹ�G�^t��%M.���F�\^�M����t�,��M�<�΋?����˳�Եz��b�M�ݦ�U��[�����< ���5,�`q�����T�ʓ��Y�p�Σ���Q��!J�����s��!�}0�T��5P���{r����ǰn�e���h��,u���#-3�f�c�*EWr��j�V�Vn(��%�d�yh��*�%�u���;�nJ�z��+?���:��>!����v�̸��4�O�u��+�>���8�׭x	���z_NZ��@��٬���7�,�~j�������S�d����hx�q�����[x���Xً�>m9��b`{�dH���_R��Ot��Í�D?����+�So�w/]|N=�����F䭾�|���l��13O�һ�K�~tv�|ݍ��̔�r�-9��pH����\�s!�<�o��#��~�R�#�8*K%,?������K�e�`uċ5>K*� L�U����#�~��3:�
RH#�|&�*�4��_٠@��e
7b7b���	�Q(�5+'��|���.���Т�:�(��!(�����K��m�ܽh��g�_��������>JH�4ŷ���ѕу���`@���9Yk��T4XS��+���	M�1��Tx���NI�hӽ_(\�Gh�V��XN�����h��3�]w���^h�q���A4��;���u��a�l�<�4�2���l7�t8�q�-��L��4�A֫� x�{gߞ��32:e	=+��:ݽ�S��:�ͱ�?����`���k����(ݐ���Eh%��Yo�?$��n8@�6m��bq$�X�4�]N'��g0��4n���X�'Pǔ~�nM����[�ˇ�9N���^�C�n���"a-�� @�g���l��j�f�(������m�~��<�F�*;��B_��	���/ϖA���8Q��19�ԮYWZ�������M�
�zs�]w%��{4J�����㎍�N��@ȿ|0��=��~G��鵑��k�z��S��y����΋��?��o��20:�JG�w�o^H2.�	7��^�֒
��R�%�i��t�i�x{�{�'�T�jwx�Ff� J����'�S�w���_�w�����ł���P���^��S�m��q~5+�s�-)����n�,���ʻ�\�?ijs�p�Eӻ�޽�a�2KWm��:E9S��6)3w�yw�1P�mp	i�%Թz#������+ą?�;a�K �|�#�^�T�-��?�~���r"�Ur��N1[�HK���V��9گ�\=��
�tM�5�����Y��>�G�����$\� ��VBi��
�[�|�LgJ���2���{L^tA�]�2~f��Ag`�2X<m&H�t�al�V���2�ы�ՀŻ�4t:L��8�����ΔC<�aIt�6^��쾨�̗�������?/������;iI��Z�Q��M�.���]r��Iӑ��z��,:S�ݢ����rt����y����M1Գ�v�������-�`;%�Jߚ¡=�
"��P�/�*���|
ePG�0:*H*(�5e�0��r��Vc�4-ZgY#$/8����M�A�'���a��	)��4j�4:��}�����?��Ϳ�7ӷ���R�oME����)�Ghr��y^E��ʴ��؅ȩ\�La.�8TO� ��,-�[IT�:9��8@K#.S �N��Iz��X+#jո�m����\����E�+l6X'�A�uG�rk%m��fh�%\o����"�)���l[X����
^�yo�2ͥ� ,
��a�K#����7��N���@�i��:T�eVA��7C�C̮[e���>�|D�,�y]�J��M���A�gg)�SMb	.~ˈ}N�[m�Ԏ���6�z��@n�(�E��(������Z�S����~�����Z��͠κ�6��.!������n�h�uI���W'*|D}�ݸx�����zᴙ��{`���;#P9SfKg�����&����C�
+9E�/�g}-��lx���KQ}<k��J��!�%6�<Y���Ԓ��	�CqD�B���� )8
(��f}_��#G�䪺����>��%'͆�WݪN{�4�QYEQ���m{E.^ۭx��C���q#�5�/����|!ua��m��%�����9	e���mo�i/��N��Y~�s���p�Ү"�8���y��6gTN֩���Ȇ�}qα}pv�s^,�}.�׌����ڞ��Dyo��n糃V ������&�^zb�������rx�X�{���~��tn�j���נ���x���-�4�x}w�X����z6�_��^��5����:5ύ������n��+�A[�S��v�w�c#�(�⊾	i<=C�:�7��>�a����0����(�� 4*�Ŀi�e?�eť���K%�m��^��B��ϩr�/q�����}o����?N��ߜ��/�b�~�3f���c�=>�4�0��Xw�%跽���>:n�%�=�-�h�z���&;�P��7y�������ӟL�~�;ӟ�ٟO?���r�������K��0ڧ�h]��F{->s[��z6���C�2��"���5�A/m�������҇,���c���[�P6|ӵ� mXS��kH�%�pKL2�̣�ֵG�=e�����F�QaR
���U� 
�Ѵ���Ԭ�GTʦ�A̋�&���`�� ���Į��ua���ʉ��2����36e�U��4�S$ࢣ�I�5�f�#T�[u^�K�m�B/� ���42�V����\ů���47X�*���U�`�ě�\����f�S|�ޛ^l����F:�p�Ӡ��X�yğ$+\�s�[�n����:xH�GS:ta�t�$ ڠ�8k��S���*�����Qx�+yJ� ��W���p�?aQ�T]��(�\n+���Tg��?�/����{���c��V�����4�n���Pz���"�M6�:�y�Pt�����oZ�UGYa��ި��;��v��uq�������頚W)(��!��\	h�Y��SOff�Bj����,!,{6�tg���/<��w�\�K�:#l˱��jRN;��2m�,/)�������G	^��9�ݒ�x�Ɗ>��i���ƭ��l|Y�djWAԫv�_�<��֋Թ�r��_���?��}�u�Vإ<m��V����Nm��v�#������t��9�;N_��,����R(K.��7s������1��t�xY<�Z�n��t�AYܮ#q�����:U�ڞkQH脯�9n��/q�f+y�/n���ѕo���]�/�@	Zj�h��k`�(���5��S��J��ܫ��rf@��\��oP��R�ș���|��c�_�&�V2lſ��0m���p-!)�"�a��zb��z�b^��7sZ#=�u��S�2s�W�K7@��9�;��/af7�7�o�B��hG^2�~��r�+��fo�E�>����O<�Q�f��m�q�&I��l0��:��̳�>�RNys�2b{�$%���/�q�D��L��{��0�^���-����0<P�/K��A�1%�Wl�L�W��g��~�`0m�ʻ����wi�HYp˥~��i�w���@+rH�F	> P�$��9�0��i������	S��@�2�01�W�=�)VK
�����),�v�*��",0?��u5�����ý��*���ZǸz&���b����#�@���3aSa��Ĉ�ԡ	�k;�𛕓�A"yʋ�n�&�=Co���в��`�i��)T��͚����Z�(;\0)ņ��č|�fXφ�������KOa#����=ZP&9� ����t��R��Xq(��,�}�����a(����Fh!E¹���S^We�������A��}'x�Ծ/(�
�� Il��];%[��3���R�6��=v��iG��'����&}鞱�X��b[&)��DR�$� A �P�ڀZP;
����{�y��*@�{fb���{��<y��ɓ'O��{/:�AI��c�xO>��jwo%@Ǣg�;�`�&_��Am�
8���ʂ�T����:=m�Ü��^��/M�K �g�$xu��$\[�i�����#v��C#���/�i���?L�=A�I{�Nu��zs����`���F +�V����c^Fy��M0nsF�����Bo�7^�$;�rj�&x�j���ŷ��:�e͋�G��2�
�_���2�#nw����g�Wq8��F�C��մ�?�7}�Mp�n�*_B#�&.Yu�I�A�߱���p�s2I�P�����_Н�X���W��c��{@�V�W&���_�Q��E��*׉��ײ��(���bc諌'�Ǒ�N_����������������{�}��e�?�è��.�m��h6�;��4V]LC�*c��S��E9�'��5�UL���N$N��Jn�ސ�#��q�ja��׸&ކA}}�]� ṵ��:�� [ʫ@Y��C�ԕ����E����$7���r)�?_8�2�~< �+�g��M[���G�-dL#�E;������;�l��~�k�����]Co�W����I����Ħ�q<�[S��P >}g|�l��F`Q��?^��B�Ь��Q�m��~�ʪ��ݕ���m1��E����_�;�)�t6�)��� �:��%��xN_F�ӯ���qF�&ta9��4xWQ0B�O�q��Ǵ�/G�FA�1 (-���۶o�l�<\w�5�L�z�3�>-����� ���J@�Vφ�܌>�4+�(�9�͗���+>������տ����������5-ܦdņ#�.J����/��+���SΊх�5nf!����
�=w-D��xk�(ś˗�ȣ�;+/��<P/�+��J:y1�6��{�2�=o��euzi���[io���8�ԧ�-I��^R&�ԇ=��M�Z��-� �[���� �1e(�,��h����03��;uc��DBu[�:^%����^/e���g�p^Ss��,x`@�. r�<2`�^�x�P�o���)�D��p��к� �)�3�Sgt��(ш�	��5����*ͷ�dw8��o�
���P� ���Ӵ)-�J�����҈��ݑ��?���U�5xZ���ڟY^c�[<e���j[�zK�ua���kpn�.m�W�Q�	�.�
jFFb�&�ܽ��ts�m�V�|Cضuآ�F��W�������s[�IUp���i	#2I�~�]�`f��B�投��G��	h�O"�1A�r(`�AWУ�����k|�����y������~�7��T����-��x�;�I�o�aj�m�� S�G�nzP�B�7�$���_�Y��ർP�n�Vi�?\��A�!d�vCdU����2C�&�%;�J�����oZ-xb�<U�m��O%�/:��Eߩ	xY��3,L�
��mh�U��圲[�>
U���Ā�:�g슲k��0"o|Z'�L��y2�n�[-�Q'��⿰`�"��];��n�i��� o�w�4���^�u�תN���M����x����w�>�|��v�)�I��k�)]R[sǌ�|�!oC��@��6E>�D��X1n3F)Ԙ�ɟD��En�C,�0���f§�����:.�nQt\ s���k��@2�����9e��OA)��i]Z�@��n�Ԯ�T�$XʍP������+/����R>+�<��,K�R\W4�U	�Pm���f����N�A���H_��̤�����������n��_x�������1���p�JH��Z]dC�%&�[�G"S;T�?�"Ê��:G�T��|�!���Ĳ����Bh|2���wtG����1wH� wV=�-C����2���М�7��?��F'�g�wt�j}!�N4_� �oE�b���/�:�^b;��c���)�/�g�8��֮�l�l��a��z9M|����`L^ɔ���R�SŬ/c���mE��y��|�9����T/}�!��l��w�m����-lN��fVX�lޭ�����W���4���׈�n���λ��S�w�M��o\���u�.���>���![^ϗ��S���s�@<8��w�hߩA�f?]�޶l��h�v�m֥K�'����&�:Ow/�3���$�V����19��)��$o�ؑ����T�A|���F�n}Y�# ����̫ �.�b
�+B�Fy"�Q�)B�r�C�>"ǒ��ۤ����k9W`���)]�E�u�y�X6��햣�98棁Y���4y�npt�Hq�x�/�眽�@C������`h�㚻1����il��_����m�ַ���լ�r����v��9VԔ�}�ȶٺ�O;��)أ[�B��ҷ�E�K`��0�
�9�T��'7ȱ�S���Y��g����N��jM*���}m |Ҽ�G��]u�[Ac��yv�zY���7u�v�� �����Ȇ�Ͻ��y�����ȣ��pH�Ʃ+��M��frjF���l�bB������Lϻ���{�8y\�j^&[-����
+�'�ûq�g~f�ٟ��᳟���я~������QrcC�l�!L�>����9\#d�]�����e{�WՙL���x��h���N\߉��X����
����ч�3��w��
�h^�m��1�?��B��y��Ѡ�iS�)�VB*Ǭ���% 8f��d�|2���� ��rK�Wt��VJIg���������7��GXe��x��8)|T �`5�71����΀�ZQ�����S1�V|]ç_o&�Jc0x2p���*dU����`��E��¬	y��=�𵧫�\�.O��T&<�X)X��m�9�TqJ#=�SQ��Ð-�ː�2���K��V��L����N�OJ^(��U�y �ǡ�A�w0S�,G�rN+n�s䗭�O�<,Ag�UH�S8����� ����
�{��d'�[p YѠ>̖�ZÌ�ʫv� wV��,��qE:+t<hz���k�r��9��:GWpp}l���>y&�ӫs�ޭr�p���]�Î���v�m7;��Ox�M�y�7T;"�zMZ������stll���Ձ�S���C�Z������۶o�W��:d�3���'�u8�'��d���j����z�[o��+<��g�	��v��	|Ϟp�]w�I���w�kH�����8��NP>^��e����W�tӍ�~�O[cCn���a��r���o�}i��L���R� :�<�H���*�2�Z9�~K�A��O |�9H���&���B�mB�(�CB0�ܴ*ȶ�K��/~�E��I��ʇ'.UR���m�(�
���l)�U��!"���k���8��
��	�:�h��@5x	�@�3/P3�T�U�y������GW�o����]��� l8���EGh!��xE��������� Mv�x�ԝ���I�/.S4�VQ���Y�e�1���=�?��ȶ��.&�حr�l{�x;��9��c�'9����R�<����|�X�P��#�����D��vrt�� g��Y��y�Ld@>��x�l���	>��z�5��]�I1�6g�N<m�F�f?�����|���<�ϻ��#�i�����N�h�����7V�y��K/�hZ�r�ɛ�ptqp������C=d;��C��y�2.|��E�񁞒���E�8���Zn��uT��J��w�W����6�[n�u�W}���^�hښ��yc�Z�[�c��#CX�@�LF7o�d�(r=��KEy�.�d�+���4 fER��FiY�z��:
l�����}*�m'*���~�Y�������
��#nVHqqP���3�a6�~!VFar�F��u��Q >��er	�շ8��Qԭ\�<<�?u#��F�w02S�LV�x�#�u�ʚ�Vψ#���K'/g��@�uPee`�qg�'@�����C�o�*�|5�Ngd�,$[�>4:��a�4�F�}�ƒ�y6�P� �+���{ 5��D��y�Mg)Z�f���:џ=̮��^�>�/K�P��B�H�!���wݵ׍���o�E:x����3��&ti�N�̱ѝ����֪o�Z)x��Q�ЮC6z2Ǖ�s��a�㘼��n^IR<F�WX�('�+_rt�ũ�[$��Ub���9(��^z�E�ݳv�J��e�.�\���:M}Yɂ>wJ�@ڳ׹�C�E�ӏ�Y�生3��g���������ǡĩ?r8{�㭲9w�q����M4ye�> ���'�cc��3�p�du��E`E�kv�����0�?�k�U�N9�;w]��3A���kة8>�y�i�����w�.�\�땢�ru�y�l���&��s�G�k��1TN�'Mm �$���6�j�l��t���?e;��.��Q5=�LV��M��I�8=Շ	 +�k��ؿ�}��Ýw�5�w�≲Z~�q0���缑J���j����!��싩��������^s�F}��������*N�
?PS4)G~�S��%GW��e�BO.�'�1V�[�Z����{���k~�z:g�i#V�ȃ��UO��'!�z�P;�����8��K?o�f�3���؀��
��C'�1������RM'X�s���]���G�(��x��I�u�s ��G��?QTڤ�E?�)m� ۤ�J �������i��=����o�B�H��O���]����-e��{'{���-|�3��X�,	<�
l?���d��OSc'xg7N%�<Ŷ`Sx�̳�%p�qX�� �����?6�w�}����:Ω?~
Go�=�[o���/�]��+�߅<�2d�����1�6��ڞa��X��'����LpY `+ٱ7�z��O>18$gW�����T�sG98�N��c�`�l?�+.�?w�u�'	�S��z@ˆN��qQ��
�>��~F+J�.0����O�2X!h�$Lf|x�_�)%`�3����,+r<����r4 l0s�<:"���5�O��>LBe�GZ8�쳃�
ﭑ�H�u`֓�`�Z'UY 1{Nb�|�F�J�M�Jy"W�����Q�Jrzu���(��Թm C��Y�8�ϐ}R����$��k�!yj`�N2�G\�E��� �8��牡��T��Mn��>U.@G�	��d0�&(�jp�2<��Wq6Hc�(�o�*�|gh1��ځ�xF��sK���ݫ|~ ��Q&N�K�X�>��M��lP���K���n��w���,N/F	��y��J�%�D(H4���,�	
��>�$[(�l�(������w[�_�C�3��!ߢO;����]����G|���]w���씓y�W�f�"��q��ț���>L^��.LX�:�w���6l�����|��&�]+���V=:��q�N:�ML� dvVNH#���sp��C]"B9�-�)ދ�﹟�[8�7:
^9#�\a���ck�9�	�?}W�K���[g2hQ�y�s�#@��F`��;'�ZG����;��2��[ؚ N�c�Fz�+d��T����'���N���[@6luxG��.�ByĀ�k�ײ����~��t$T�8Z����Ɩ������p��&��<�蒗2�Î�p@x>3~^���jǁqI�.��)���`�P�-�##��C��A�8g�ݢN�P6&���@9py�D'B�Mp,���14-��(<5~#c��p�/�'߅��Jn ��:)�H���L(�r��3!���3^������2���Ч�z�[��<	�O7sG��|؁��,�pg�9�ǫ��*�^��|����\�A��o���,�x;�"s��4=��C�=w��z�ڕ�(���n�ɋp���g��2Ɛ�	:���=j��5nsĹ���nn�Bʫr��;��ӧ�#�@G���ȳ�#�wtpՖn�j�	���۪et��'}1�E8����BEY9}Ϳ��*� �T���G�#��^9Ь�N�C� ����[p~كȀ� A9(3�/e�]�"����B�O��ʈ�|H�q�i0lc6D��6�+�mx�6�����̛��/|���P��]���3+ɬ��F-:�_�p���q�)�}I�����Ѓ%�����>�6��Gz�;:�n �RD�r �B�nFL�'Z9�r͖CX�MdP�k⧼S� ҦP�Leƙf�B���F+NrO��[Y-Ў�����`�n�@����n���)�mr�p³
��X����Y�<3��k��U =fu������jK�ƈ�zY� ����`���g�=���O��gb���1S�u={>��_��\�����%�A)wiv�F�@�`�P%?r �� ��2�L9��m����3�ji0?�Qq�E�c�;R5Ж��i@��퍓P��eo��d�O�//̻�ؐ�MKF%'��@�:6|���6��|�{lN<������ۜd&;j����8@��Co��~�0�� �xph�/G8Bc;+(�.�H���+�ꨀ��h/�/o�a%�Q;4�������p�ː����#���������Q2�^�'�]%<�9�{&�j��:�V�z�4��~=�f�K��qiѷ��@�dKŷ�FJ' ��l��/���!o8aE3���]Qu���a��$���<�N�����2�R�雏�A�C���n⃐������+���M?������G;��We ���3|��%wb���P���N'X��<����o|���_���O8�q�T�u��o�M�(w6�5�#7||�򙠳]
|>?\���r�����UH��'~�<0|���y����	�}b�^�c?�#�}���;ڌS, P���c�L���5u�O�[0����;l�bр;�i|�)���+wXNH��
 G�1tMO"D��w��26�� �҅�1 ~�wS��cc�ٕW�l0�d�^���4c��c�$-�&7j�e���q��f�������F��gi����8��q(�Ѡ۶��&+ʿ����Wϫ&�A!0���h\�e|f1�C�XeE��F>;.r6����0������'���:֞]
@���>:�N��z��yw"� /�����d3\�J+�%1���
z�&���c���v�1�9��u�"(\h��0 %C`���K^��rz�~ё��Ξ*w"�=��]z�5x�By9b��M�-o �����J>�un���? ���:�IE�%v j�N;�� �U��W�����~~`F����y�u�MM�"���q��od������J�%�E`^�O鄴!�����A5�)�5ϩ�S{%��sG��oA����K:m�^L���nPsn�1[��t�jf �~#��s��Q����ӫ��)�Q�E��	2�-د7��˝��_ �?�W��c՗��3'�{6���S�3O?�s,i�`FC|F���JS>W������?;�n;�%Z!������kEE��y�Mp �q�@��Ka����mj?r�-�\����t5��9}D#�X������;![̸���o}{x���yl��1�@��,�]e�ޖ-dM
������K}_T���\L��#0�X��xƖ$V�~��/}ɟ�fu��ua��@�8m�4�D�����5cu�~
N�7@յ �#�����M�Q�$��#pH������s�#�j�2�Ʉ/�~mW�H���B*��;��N�U�ۖ7�)�|`<t\&W�6��W��M�t�Nx�.޼���e��������F�����;ܟ��*{��]�Ë�ˤ[���~M��Y���ӟ��WwYXÞa��t"_�"���+�+wl���
�q��Ƃ���3�-z���]��1&���_�%��O���S�X>����^ldE?�U�ea	?��"/����܎���p-{�!���x�����bp��[�9��]D��:WSR
u�jdϾ��J� ����2x91�V�"@��9����Q���ʀ�����r�p��W�\{��'∲��/��E��Q|�Q�G5{��>���(̍r�w\y��Yc��:1���m�WN+��k�&�
@%y���4�{`S����]wr+�?��>->�̋����;�" �ڻ�H�%A��j���V�h-��P������e�SG/Ђ;�u*��+ ��  �Q��˼�C�!	��D��a�;��e�c�%.�kGꖛon��f���|�Bh_^�����¾��О�}�ծ�=b����<�s��9_9M
u�����
��4�L����?r!c��o��P�9�Ug�֮8�;~3 z���׵�����?9��Fg�PK�; �ן]���Z2�ƀQE�����#mI�΀�Zy%\V��w���
o*�x�Lm�l9G��6|��j�.���w�xPm�>;��5a���˽j�ڠ�Qr��HWp��a����g�Ǚn�m��U+n���F�'��U��G���:+[�No�7��8��#z�"/��d�s��>{h��)�%8�]7�T��V�	<x�����[dm\�p�<�4���� �g@��q���&
����,�,#��1B&+j:��&R��_�����/��7&jLb,�٦�l���wa#^������Bh5�9o0��F��8��|��	���8�������/@���&}@��o�%�C�p4]�*$_�gr�Ex��+��=Vo�s��#�&4i�������<J�r��Bl6�p�9w��Ipig�(�DՑqQ�����V>)��&_G�s&m����Odfq����q�Chc�x��/F�+�l��˚�����3��� ��@�����G�sr��<���ɾ�^�A��y�����8������5�>"���hV���GYu�+o���j�d��*<m0��bh|�od��rY�f2qR�����첲��f�����E���M�őܽ ��9ʂ�C P<a�"��83Nf. �_��Qa�`�@����۷��'��l�Fp4N/�G���[3����g���^	W��@%Đ�Y(���8����1��~���=SP��B���a�F�aP�����7n��}{�]�p��V�^1<ppx���<��d���(92���3 �3�Z��Ȳ�!�(�;�҃C�o�ӡ���H;�T:p�%·�c���rP8�.Mt��C9��6�=�W��29FW�i������t�w�)t���=+���p�8�5��+�amy�[i�t�@��zZƂ���_��xxU�4��8S��A���v�p�tD٢cGJ�&U�pt�~d8��c����|-��^��^S.:�{tv_�Է��}�@"�t�����o2�L�Qt�.W@�zy���#��\�X��\\n�v�5�٨��'�,������m�q^�� :Ǵ�^�<�A��%���|�ZmJ����x�ӣx����♤3ɡ��ҡ-ܞ��#m��B�Da/��!��ࡃ���ڋ֍j@�]n�&%i⓲��\?�{D;��A��d�+�����]���jg&u+ڸ�C~2���.m��̓�-�B�I:�5hYך��r�s����?�,z��u��y�+��o���S����r^s�Þ2ư�Ja�u�2w�W�"��Ipd~�?:��9�-rҵ~ԁt�(��}co#��V�c�|�	�rl��}��Fv	�5m���H1M-�*Ng�	Ӻ�}�8�
8���������A�RW��yC��{����i�Ny<�P
���u/����7�6���������.*���Gf}}yg`��4ꇞV�>`���?�36��S�=g7��L�󶨱�֑#^a��M,B��=&�L�/���<+��#~�>�g؂���'}�K��۽�	5| ۼ��-Vg�W�����ه����������1� +�%��결>��&	ڔ;�L�)륗^���_���-Y�8b���ܵ$�L_Y�^}]p��k�ӯ��<�U+�8��uv1�8��퓳�z[�ՠ��ؔ�L�Z=iLZ�!0��R�j�W���ipb�C4,C�ˠMeQ cF��)a,��)Be���O�1��xй��֌���G�wdF��'��F�,)�=�4<��@H<d��Y�a98u�r�e�T43^�,QXi��~��a}�{O)��~ʛm��Aayo�c�}���e��W��	G���Mǧ�@�>e\��82�zVO��:҆�P(+�D	R|��y9��/\f���a�C���� �� q�f �y�z���c�7�N�G�T�8IB��A}�'�9qЗܤ�l���5� O84� Y�a��f�;�w��#t�M���+V�G|"�=ᇏ�ȹ��c�0�0�N'�j���|��}BT�kB�9*z̴��5�Ǚ}Y<��f�/u@f8�T��ݯ�k���˻�:���I���(�:w���i�(W��s~禌!2lv�aj�����]�ڪ���d�w�����[n%�p.1ԬZ�z��n�]w�����U���4o�%�,�7)��0{�xM��@��`�i��j'z��-�vMޯ�v�_����<��~xۆ�s��ܥz�v��s<��m:�	�z��?nn�c���� ��y����J���=p���5��i;�gd�s�xk�U�5(��|�����[N]�ٟ&��S9��pn}����jo�a0�a���m��?ʧNY�����jl9P.�I:y8������}¯�b� �j�ɣxa��.��Ok�C灭.&�Y�ՠ,<���$d�r.Y��9v�|�i�MOH�x')2�.�Ƿ����+_���qi�ꁯ�yŻ�`�>y�e-����h2C��C���'�Bt�S3��hU��i;'�z�C���(��<���G6�+ۡ��V&��.|�2���(�G��~��N���zP�����4a���8��y�ڥ^��>1���1$�+���I���m��6mGt�A�i����$x������~�'rx������w4����`���x�Σ�^|���={�_�{W\q���Org�@�R�4��4y�N;�<$Ǉ-8�mD��p�����/������S����|T4���oJ����o�结£�ܵ��+�飏�:��vG��3A���`a�[��t^g��?pHL���6����@��H���@�Ƙ<%΃"4jSލ˓|�ƩEP\�^SV�t�����p���ʞW���p`���L����8&?�c?6|�S�򠇣[�r����Xf�E���J���rÜ�mi�;��	Ұ�A`�A91��aoil�`e�W�P&q��}�ߚ���'0I׷rT!�H���t�Rt��g�+'E8����y .O�MQe��ÿ�+*�G3�ņ��u���� p^z1��qV�k.�/B�O<88!��~��I���c	� ���M�`���u�]OǞOf���p����#�Bo��F�c���,T��k�����V�Y�9wNx����}pй#G�x�}缌�o�+x���+�~�sP4�{�������:b����5XԍUd���ϑj��m���e�9�n�f�u��"DR�ye���Dз��x�&8�����D�j�OtC�?&�|I��k��r�W����?��LZ_۷W|k�q�WDx����{��v|�鼳��'�����_����O��@���裏:�7�����������O�~�;�7��m�=���~�����W�-��o|c��׿!����`��Ŋ
GV6�mt�_�������e��;ʥA��8�i�À����5�	t�	�����c��W����>zy8�5a�'[��CM^�bGQq�f�4�a��v����k8��,�3�P}���(�����#�J\�<�IӶ���N,��k m�5}�;&���wx�!�@���K���2�9�\oU���P�ϛ��d�6`�����/�º�XC��W�Ax�z)��|˹�#o;x��t��]��JqcZ��0Zܨ[D��j��q���D�ʟ����N/hZ~:�,���s�2�<S.!���M�r[0�g0y���	��\NQf �(k�F:C:��<a���?�rx���p�KiI�}�k�ܵ>t�u/�1�`/�@�X���P�U�u�S�����O|b������?yj�˿�����O����.�H����Et������!}���^A��R�2�p���x�A��f�8ĝ	ޟ��s	'�S�z���?'�9<+��7����Klg$�L�&���,Y�@���EM!x���1�� �CcT�P+f\Xkq��c�fbb�%.J�1�I��#�(lt��#NBaoﳽR�����Ҏ/J�����،����P*]��?�Ƿ��m����?��?>�#G����k�Y6JD>+��/�q,Xi�qx��.(<3K�С�(��V�u<�=��ǝ��,����fAHx��xL'���6����n�$��
7,C^��ٰ�0�!$"�2OiC��O3��I�P�eL8�rr=�E���l�Gg�8�h���i�<�kl����C�<(eĝ�����V��7��7zL��=�K��")�h�w���k�����ޮ 'e��5�CHy࡟L�|��:���z�%31�e��@��Fϡ�#��
��נ���gpvq �*`�ۓ�TޒK��s����� ��	�����H݅0�_�C��rv����.��B�����M{0�ܿo��j��N.���={���}i/K(/���q��A��g_|Yvp�&M&dY�g�)q�C�h0�a�Ƿ���3��!5&4o�����U'����3��&{����Tv���~����t�.���v>m�Pm.�������8�5Z��U4ic�1��t)�������h����&��tѧ(�]u9M��	�Łe�~E�g2��;�o�?���.�+�әb��Wdpf;+��S��+��[>��� p����ѝ�3D|$]i�V>�w~x�5�t�l�G@�Nȴw��O뇬�5�ϡ�۴�u��+�����>���|���,�$阝K�����^u>�i��b�Iz�% @�Y7<O��!ѽҷ�����Qh���Z�
�sƴ����D��9� ��Ҭ?,ޡ�����*D&z5�����8��3�ںe���L�UW�m'�=�C�/x��C>8�v�m����sz��/��<����^^���(��f�L-z1G�?� �y�.��!����-�JLm�~k�Nb�E��"�����ǿ��m,ugBWr�	��?㮲�g5�^R��٥o�7��^�q���1���`�����O�~�q�|��hҀ�����p<q0#�J�-�Zu�qY��B?������nk�
.���:&��5�B�����Cx���F�})���<��ۂ�դ8VP�'~¯����)B�yAF���W�R�u��b����'����pĽ:��p�#F��}^���|���x��e9�����d��}��a���������'-䆑���>7����Q�|S�pl�"6���x�Mb(���ǘ�P�>ݢ�����
]D�Ꭲ�Nh�m���G��W��N]�2Ϟi:;��0�=Px�3� �h'vf� oa<}�}"��ҏ���ç?���Y-�����d�С�����H�A�ͷ�ч|=-+�ԕ}Qg���9��_ud5��I������ �}� ���HH�/f�l��-&D�'8�%&B<������j7�m��g���7�'H:z��X���(0�j�	�����8w�`�M�w?��>��O�n���e_5N�3�<=|�4<��SrJh��+y2Qb�`�� {3u���S=]o�7��c�6&;Ȕ�~`k�J�0�ig����c�\0���e3�-��V���#��	l}	�mY|E;3#/��}�]��~ >�f���A����RN��b��2B;}brV+-oY(�����Q�?��`�7�Q��)�Bh�N �p�J�|�q�/r���K����;<���W�Hȁ6`A�����1_���Ӏ��:�a"g��߯�	!�����r�-��\s��k������f?5_�b��:"����9zf�W�./���i�`��_�����$=�Z��s����g@�S|�Bh2��y��΍t0}[���Rd�L�g���)��z�Njd�����j+��h�:��C����xE��/�h�ҷr��C�74�N=�^�;×qt�:�������9�B���*�Np��<uc1�����Mh�+Z��_�%/�1��I���o�~x`��) r@V�ǎ���6�5>��&·}���1(g��� >���!�w�3^h������>:����ϽEy�++�^\�|2�/�ߙ�N#�!�";��5l2Ƒ޻�5;��F9�g\��gN�.�k�J���5U��W2�.�:y�yz����g{�����/��p���ï:���
�w���ǒ�sc�K1���.g׍��bMJ(�&J.AKX�{��������`T�C�����3��A,�Ω�(4`̋~O�4���ש�����vr�ˀO�G�4��3Ί5/ufŕ�/�O���������_����*U��f�xS�?s��ݥ�v�W8�P'N��w��/��/��4"�J_��<���-u�]:�x8w�����
u�s��&Ȋ�J�8蒶+��#`�]����-<�.�E܊�8cy44w B�ʛ�C�0S��N�>F oCpk+h�ݜ�5c����.3��|�������T��#CU�/t�-�}$.����]n�J'd��n���lG�
� =�n� hԍ��d�n^Eѵ��40J�5 S�����^�n|��O����KrzK�� C Oߊ�^Z�6<r'���TX'$�����˿dK�lh�'l�W�^뽺��ħ��R.}���>����g�"�k��:ؿO}r�탃�d�F�����j:���2�*�u��?p#�R�;��y?����a��m�E�s�&��!�Ⱦ�|\��]���]�e��=��#@9��O�i��C�ħ�S�Ό앤\�io�H¦GBY�)_h�JO�M�&�+��V�yMh�7,�oyBm�q6.Ν��W�(����c/�Hv�ң۔� �L�6}� z�y���S�D^^��ϡ��o�rM������A�W��B����6���K�Gs_W�i�Q��r���^�QH������<��'&{�!�-$�b�UPm+���2Ȁb_��S8�<�C۹��Cƣ�t4ӊ���m�H�S��a��/�Z-�HqM�A �A
z��������ތ��9�gʦo�FR��R��鉂O������LZsv}���8���k�nh̶C�Fg�Q��Y$
��̙ d�A��Gt��&||�<ck�\G�{Վ�}�J~�-7��[x�8$;���u�1�Q���r[�E׳���B�Ya�'>юW�+���=�^��^�_����桴�����k�5��*O���o��ƊU��`xg�ЩM��`����������@K=���_ȃO��گ��ަ�~���.�䉧�{�I?�u!g7f$�ڔ]D)�󀗎EeU���y��ლ��V�Nd�.�k5��|
G��fx�d����e���+�������UBz[��a�cd6���ï���4"�����A9Ǽ������{��y���ȪU�a�g�Ue3��8�n� qv�
�r�m�%f7�S�8�|�
�����|ex��|�e� �錜[��4_���Y��bfc�Xq��n
��R��s>)=�Dtl�ب����("G��)��1�q��1��D��c����pL���� <�K�+���th�+>\���d�9��3�����Z�pvY�����y����B����SET;�W8�]�;u�M� �J���Y�<P���<��ߢ���m�52>�/�<?#���Y�w?0���7����O5����"2���lrv�@�,uK��HB���t��b�b@�	,�Lڇ>ɀ��{�3���f�S�J/+|���o3H����3�Ȗ@E�v��z���S���y04/O��ٻ	X�Ƞ��� ^��b�
6-�Y��2?�|�&g����`Gp��{؆�}�s~�L���!�����W)ϓ�F�3(Z�����&������k�@y0�P�A=�_>���&m�	�xt�>)^<H-<󫣝Ͻ�c���J���}�-��l��\��&�d�ܜ���ȉ�	�Ŷ�d2 �p�^xo�'2t]��|V��{�a��+��֮�3�N!+�©/e�3\���5�\[�~���}�R��o�w�蟼�:!#��z`� ����qN&@	56"�7�%o�"��:�c���_#�L:A[�<��o�C'[���Wp:���B]���4���ve~�o(�	t�R����]��Wۨ�k�/.���A;��>E��-n�9 .�s=��m�8��>���Nd�Uɤ����U�ϻw׶	r3;:O�ȓ���6;�~�=��P��	ߍ� N�<�>la���q�(�O�&N7[���� ��<!;6.�IG�ș�t>k_}f�捶�^�|�x~ǋ���淼��&��ʿ\6�umP�g�Q�xX�zӾĻ}��]c ���]2�=� g���׆�o�Hg��v�?�.�Y�]�1���SB�cw�
���504q"n��f=���N�h��@��ƫ����`(��ܙY8O�e/�U������;;���v4Y���:
�wx��G�|�T�SP���Ԃw�Ńh`83���<0r˂�63[�Efo����\f:������L�ɒz�.xA�P��V4�M��WP�O�ۈV"b0|�n=0�c�Y���{�[���3������&>�[��t:6E�ҹR�����7�s��<�HUG^
�7����1� �/g�'?�SÝw��}���e\{�5�9^'�u+����)�'� �C�q�1a�"������U��s���I_ҥ��&��@�h�s24ʧ����bt,+����_����'�~��Rۙ��m�����&(>�_��f�ob=?il�ֺ	$~����~4^����7�n�:M�y`퓟���-M�ڵ�5i]k��F���].�Ʊ@>�	��_���9q�
�[Aѓ�!2�A����<��KD��v⸝n���3ˠ�;U�V�����������~�}^r�����|2X����T;T���$��,�vv%x%���U�AzM�Sd�9�=�Gx��8�Y��פG���>�A�}�q��]ɷ��N2��tu�T�xmtR���Zaޚ����P+�=��[�qL޸3�yK�2�rǕrzw4,�r��v@��5"�M�_��3{�ؑ���>����a��W=�Qo����e��v�c�PUK��c�<G�)�*"|7ooc�gY���r�S�Z���Lv�l�\�q�7t2�)]u��L�qKȑ#2��͓+q� �Ep��S\Rc:}���ccʤ��&���5��Cr�>Wvr,�G����`�	\��x��;`��ߡ>�w���az�'���^~�����r5������D���	6>m�4�lR�E��,�1��>�HC~��NN{����<��Qvm�YG&'8ݯ~���
�~H>�.Yfy8��Ѣ��<�f�����f�F�21�ݿ�w�-���y�]���^�=<���-g���\�T�XT�137�y�7���=l��~�A#��T#�yH�/3l�[e�3���^x�yu�<��~[���*@���?��=w߫��S��.��*��|�(K3A��������~=�!�����ya�84�2�݃����`	��2j��3��s�Ω'V�̯�(ƭ��9�:�W�B�<��7��<
oʳ(��)�f���"��
6|�	�.�e3|:{�%�՛�s� �~�o����Ȭ�2	c֊�YI�0m۶��S�Ӄp�R���~f�8�|Q�z$ctJF��:mK��G|;]�O���*M�\�(+�쁤�x9y^[�A��9��0���������wo�Y#�<���BLK.%�����5����q'n�|�<T:M��n���I\�ۻ�\�v�zx���[�o�A|m�>�l^=CN��ֳ���-���;�t� ۈK��ں-|ʧa?�?2 �p���gb���������#cۛp�_�#8�a��&�k���[p�������Ss��!��SrQC$-�j�tɽ���V0�kY �V_E'+�#�I���UG�S�)>k������|�S8����dĎ�A� {�v�L��k#�� >���kx�d���8r��[�	�$��.פ��z�F�N�ϖt�~����#��c�-�p޵�û���V��<׹ej2Q�㩤C �)H�Lq��]�Z�F�>yeX}�y�F�Ц�&���Ʊ�_�H�S�ͷ�z�C�
��RMhQ"�Р��'�1 �=���A�B�/Z�.[���ȽdY�?e�W��W��l��߆P��'&vȚ�Y��;�YdA���aױ�îW����ț|�'4��7k2B�d������~��^��_�}�NZ�,�qǂ�3�?�+W%��k ՝7�x������"� ��چ6�P���Vp��l�p�n�������o��p�]w�9�~A��>Q��s��A���nX�v�a�!��`#�P�++�*�"deE���Z� O�2�����@�~�
��H�|20(�ѣG��˾XVJpt���Ճ������(#B�B����a�W,�g��-Hʄ7�l� ��ƆG�� �88�����?�s���)+���(�� ��ԱzA.��;L��!
�P�L{�'͡]Y>�5����?�f��^�!ņrr�@��,�/�������a��k���ɹ��^"+چ�qpׁ��%�-8G�z��qk
�\�d�>џ�5zG�S'�.��ʐQE��Q�:���5@`ԠE���)�#�lq�M���,x�<������"��[�/�X�M�n�w3b���
��<�,̮⅌3Lq-�x� ���<d���6$ޝ���.�-X��	��P� {Xq(ؒ����05p=���Y��[yR�>*�6��k�ҡkθ�E<W��%�����ƽ�KG����o�3�.,+��C�΁�I�,D�͹hx��z��|l+��o馯k��!��Z[��5�	��fw�GdX<U�Bt��yB-��\Gu�^�S[�T�F��|�~	���J��4�����R���'<i~����,��kla_0Gt'��#޸p����mӭd�U�GNK�!��N�e<+G��矎����JU�dZ@���j��1A�\��G�uD�ɨ�j�	R6y����?�*�
p^x����iB�P��f�/�� L��F+�R��_���>|l4�ԋ_l}�&o�����T�k�W| ��c�F��f�`kp�	�=Y��'�F�_l���X�4�Bf���~�����8¶�rh͇�h��a���v��ich�H'���g��ki�1��DO�g\�;���xVt�+�5�Mk����/r���=Q�nW|����'���쓗�~���ꡇ��8�������٭����Ta����pl�$$_W��Eh�IJV�����L)*�H�C�б
��!1N8�|��_��oo���A�4xзAUC�3�!�r�2y	���ϝ �EщsgR��� _���M����ʗ�2|�s��@�B�>Gߖ+����o�����A.VJ���(�{��2��Bb&O�
e��q�R��/�?.�2*_�)_D�:r�Y;w�\zw�4_Δ�A_2` �}�������D�r���d}`Ӯ]W{O7m��1�a&釖��*�tF�-�Q����}�7�8j��dب�0 �:!�Z�5YPU���M}hc��_�C�[��^s�}��ة��_|�ɔ�'ot����έ�:�1� �z���z&"\c/��)n.m�xPn�]{ݵ޺D�a䫅�0�w�*9�������l߶U����jz�}9�����,�@{d �����s0�����S�U;8����g�@���n�G��8����1>D�9�tJ*��VpJ�씟��Ec�RGh��?(.er�Ν�0AbH�u"��9�=���hD����e�* U����!29G��`t��?�K�/$��W��S��&^�&���ߥ!Mm�C��f��c>џE��dB����O��3��_�������Qy�A'k�rr��rjth;t��p� )�������ے�	o�|0��+�B�ël	<U@��xf Q��a�;ʡ�	߅O~׭�g��ٔ���t
��565�ԓ<�o�{�QE׻p\�]���\t(~KW����~�p�o�Y�*�v�#�E@�O����gx�^�ZŸ�Mc_:�R�4����8>��گ����z�g��c�����+�D�m����8�;}�T;���ҹ�ʞgZ;y����]^�섳�ޏie��?C�@T�ֹC�L��tN�e >p`�_���X5EHԈ��4T����0?q�J'�1�Ua� ��ܞ�̆�C�%t�it����x�����rN��w�S�mG�G9��M�P��S���O��|����l��~�k_���)�N���Y	��Qz���\b8����0A�Iwg��+;��K�N;���2�(3N� \f��VAN1.�f0=/u�4.�G���AԿx[���'�2)g��Ч-�9y��L��@b@�@8�l��C%�aH�}X�O�e�3��B�p��o]ƙ���iK�0Pq2"{ha��g�*�{ҡv��fr�K�m@[=�e�	=&�{wY	`���7��d��q�c�i�K{[�M6�WZ`�՚�QF#O��Rh�(X�.���8Υ4<ʸ��]^��gh��a�|�lӰq_�Z�/��ڹ��LpX�ۊx�*�$؎�g�c&�E<@�<��;�5��x�"����>Yq�I�m��W�ʟڃ���p��8�����<l#���_HR>���K���G�c�m��Ѭ���tS
��I�����ڠCqq:)'��gE�m�,P>i{x �#��������#蜯B���5A�]6�K&�Lx�9T �M��(�,����@���"ì�`��c�j�94~�R�4�z����E߂'�������x��mjϰЖ����p)?�2�ȭh�]��˔Q�6ь:u���`���c�p�K�-�&S� ���CU\�c_|�+w��� ����I�O;��_ŅO��-�&�4�ۤ����m|�\cb9���+��!2�5��n���y��>A�#��H���}^=�yH}�||���Ѝ�z��bB�WՍc�rN��vH���npW��,�%��?�I"?��G�_ڼ|Ї����l~XO/|��fтW���J�Dچk߱iiz��,9�l��˘�5wک+������$X�Yv�.�̽�ҫÓ�{��]��/���E��;>J�� ��C� 4��:��]\yՕ�X���)�<0k�~ټ)�
3�PvVQY�'�FDv(*J��2�͓��Ny��� V���Q6��P�o�)@���h42��#p0X�eec�,�K'%�`ϊ0t�z�Y��|�Gwb�Q$�{i�	�s�2)����p9���Pu�J-A�����;�ȬV�K��>��,�Dn�
 �T O�y2�gE� �{<�I�p��
9���
H�&+f�ER��%?�V@�Șc�䤣>��Po�_7���{[yp����E?�KW �H����Hh'&D+5SFg0D6@쯢S4�0��A6���m&t�����@y��[�iK�~�Aˬ\�;���-9�u� Wx���>0�%�o>!>��D�[Uis�H�6,�f��8h��Ǩ:������A��(��_tY	�s�Wɉ���k�+��!��+���s�ݼ!�G����-/��Qf�Z�Ȅ�ɖ���nV�ɇA�qn�!VpXY�����Lol��
d��Xo2������co'�,�4s�<�2Q~��G�%u(�Z���ʠ��W��3��4h�'\�er�rCڼm�<�q�4�K��M�@?���������SF+Е���T��G���X�,Ԥ��dDEZ��QQM.U砷|�G���a�Sh�#z�~@�,��"So?�+l�m>�#� x-�r���\t<x͖�*{��p��MJ�u=	�?�jo&!DZ� ]机��<�3H}bo2n�W��v�Mt�1�rz+���?ѯ񎢓"~����CXu_J^"��?@��v*h��\�M�s3q�����y��>�V��s�/���N�f{A��p�����B� �:��ZՕ@���uw/i�Җ��a�"�䴾*��G;F��/V����gGꎕ著��슆}�6�"���T�n��������P�$�<ȍH�͈r����گw�~����.��}E�����_��l���H�ƇA���@�����!0F
�E�Oe1�e�B�W��;�(\�!�:d6��T��-毤����Fqy���߅�,�x������p��d���Xs6W<{�p�X
�1A�{�0���<�5�Cf�p8ٳ��,�n�3���0A��u������Q@�X�"(�R6�z꺀N�ū+mV��]���.2��p9N4sn��y�ihf®���0<�s��| Z����cr�(�L�ή�h0�q�zͺ�õ�\k��0ȓz�,�A�����Ww���6�e��=��jL;"w�� ���I�yUm�=�M/<0$��㈾sM�E�ⱥSg�[���S'x-u� ��\6�;m~�&lo(�t�8�mp�2�)�~�AV�V{,�F�EXP4�rE�����m:&h�͉jD�	-d�1�$g��K}��g�Fmyβ�J.�n�m۶ݫ��Ǧ��٥�q�(�8�'�͋;Qđm���41����(�G��l�+���I?��olM���9��-񃓀�x#zz3�-�
B;AۡO�W��Q�rI��}o<���d:�+�IIM�7�V0[�������|�(��NQ��@d4��iP��)x^`P�"�����.K��},����z��9���_;��B�da<S�ȃ������st�xp�@*�S�E)���l�%��ށ.��W���B+i��ΚL���B�Q�㚲J?Mm,3@{L���v��kJ8���c��C��s���;5��VzhL�qO��U��iТo�
��$wx�3�
�,;�v�#����~-{.u[�K�qS���6t�2���&y,*�'x{�O.S\�&Z�A��w�[�}�V�0Fmߺ�c��V�+��+~�ؑ7���1���ˬ�~��]%Ui<̶c���0xqM9R�Q�,���S<Pt�����)�#4t:;��c�G�s_����(�� "\L�gF84L�:������+��T�]���N��@��Up�i�� �ui���u����A�	���d�,n�Ҷ.[ec�������a�P�(-�F�V�=���3�����d�/� h�����v��A:��� �uji����Y�8�d��u����߇���Ȅz�V8ȅ@�VT{ �[�#t����q�dL��ލ��fd�<����d��N���섉�ʕ�9���kTċ+]�Vxh�렗S_� �s�'<�a���i����e��uV��7%/�����X���#?��$�vL�y�n&G��ȑIn������I�b{�r�Ҧ@;�l��������2y���,9�j�w�����lh���]m�P�K:5�(z�]
��OCH�'B\!�F}�>q�vaHw�	(o�d��b��q�^��30�;���|V��������yg��)o�M;PGo?R atv5�((��<)��3�bK ��O�T�6�hb�hS=Zy-m<�s�*��9t�8ڱ���|�+��>�	��1�_��*�<����W={(~������uv'�yXH��G-������<�ט�ٗ�^��
 y��Ů��Y�6�Y<�'m��>�6�����,=/9O�x���4م��LS�6Â�ѵ�rv�W:'������6��� �n�e�q�mx@�����-�m��8���˿����{�.�Z�_�3<��]ߤ&����M �Y0��S���������ل����8
�ĕ�e��-w��L>��+��Z(�9�}$�H6|"�K4�F=��14�A��۱���w����B��ԡB���d��t���/��b���Z8�M��G�|E?!��|96��#t�i����Gh�$�O�L\~i�	Ѫ�Z7�g��峑�*;�ā�n�~n-ِ�,�`6o�A �ǫ?��hK��L�p��[�A�8,8�̓�L]���jх��];S)�8%��������1��a�@Mz3j���Vd����T�q�;	1�A��7M�˂��p�B�"s,@���)e�����UZ&��_ƃb	��I�(�ȏv8wV��4�Rv�v���[����=��nGt�K�a��KuR����_�Vq��~�?� 9�جz5�s� 4�K�@�L��.A��f%����&g�����¼���]�5�n����L}p{�2v_-�8�>����Ȳj�3˾[�]lA��.퓏� E�C�r)�5���HzW����%8�:��C ?�,3�T��"Gn�M�E�l��+�E߃܄��1^��w�Y����к=��a�$��vd'\�%1F�m$����]�p�8E�R�Y�z.���#t��?f���r���\��r�]����n��7�"�8C[y�eڄ���6�|p+�6ٱ
��K{+3� �c�QA�˴a1y���cRi�rv����d���;��?��1�[7�M����l#�,�`��Rբ���͛��X5���5�둣o��q8�{����W�������Y
�WN!�yS��:+/E?F7�\�rLe�yw�PYȋ��Հr�g��I��"�e��`�V�����,|�^��m�dP�e(��#=�N��� EmE��	b&rɵi�3���#�P���s�
��q줡�^.����E�;W~P��H[Hq��+R�N+ �x:�y ]�,7���6��#C�>�'f�|
r��-];�8��ke@tf��>8kq���r�J5N��{�V�Y�.G̳j�*g��af���M����[����C�C.�d5e�f��b�W�p���vКꁴ>���5�i�5����X#N g�-,y��N==A�^
�Wi�L[��!7d@ȝ�K��[����kθv���<�z'[=<�+=F7����m��r4��8�UԿ�-��`C��UdJ���!�W�l�n���O��."6����9�Ƕ'z6�-A.|EO����U�O=K�C@�2��Du��˼��NtۙC�PP�U�RXi��L :.'9#הit˒��g�'�3s�ӟ��,Hk�-m�F��	0^s�MjY�x)b�;o��29'0�U�l�$�#�ѵ����m�?_N����������Y��W�˥�U�bW�Z{H��+����yZ]5Y�O���&g7PmUq�/r�'zr?1,ު�]�h��e�}��҈ær��lc� ��?�[�Ae@���/�P,%�h��l�F�X>��j�"��+�<L��+{��=��P[��+�C����Es�8k�<�FA�b@���v ��@堍ذ:����X�������qb��Q���m]d�J�B=�c�V =S�8����\��H-�Z�^+���=�R,V��q��1>�W��a.ڥ$�S4
D��3 ��"���:@�7G�(3�*�ρ�⷇3ކ���8���	6�����c�
; �@�0q\�2a�J��2�#'m�j��J�"qǹ&?��خlNT:=N�t�^qB�:"u{&ke.oy����E��|qmC�
n���ik�U�C4+�O��f�r\��y��-&M�C ��m7�/ ���Ȇ�53��M���,��2�R}˽D�3��d�zQ@[Xl����+ ����]�����'\�]uF������W�3�ť�ۡ<�/�]z����؛�Hڄ~ϑ���3�,S�3�R�zF��K�^���i�b�3��n�Zu�'� �R�%8���^V�Ezڐ�Pw���fT[7]��/��'��?r���
�Jѵ�]'&NM6�'z��M��?{��W)�]T[-�G���B�x�y�ƍ�� ���,:L�Ѓ�?���}��S�_�K��Gʠ�Ǉ�:5���o�vZ}��f�zA����rS��zF��Z���z�O��u(���p�П�l���E�r�ǭ�y(�>�ןEt���k�7���З���w=VY�#/tHW�Gl���ѷ�=�-�7��˼��o�-�Gc���gNO�O�V����0�7�K_`��_��Ї�s� �Qǲ��Uq��)����P�xp~�������XK^C����j���_��E�����_�6�'�xb�٭0u�����3�)ݓ0��s�`	F���
%o� �W�#��*M�Ey�a�-�V��(�6(Ƿ�sI�T����`��x��x���"��@7�6�:q��z�]*�$+�p��
��n�:� �P�i>?�<�u]��G�aQ2���Ո��%��Ċ<�o䬮�#�tS�S����b^ua�гV<��"�S�����;�vțΟ��8��40[��Na#p
e�dE���f��Ϣm���:��;��ue�����_(\���N��L��4뺗����8�����_;���ݔ#\���u�_���Q!O�N ���9���nfgf����'��Vd��-^r��Գ�@N�}G�n���)}4ĩ;�$C����X�/Z�gǃ"����m ��!sIhѢI�mmm�.��>��
� ��~v\���OG(����/}U��[�J�vf���K�&�ѿح@�^�Y�*]���V��l`נG�ߑ?/�	K3A�ڮ��T/t9�+��S�ދ6.xقҜ]��ur�D/bӊ���u�W��¯<9�>� �s^�Ն���S����'y�M~�zI7(Qۅ���W�a�kZ#��ky���?{^�|:�4f�0+��8�Pe��5f���p��{��doۊ�Z%u���C��B�B�5V�U;����O|�.5�̈́�l1}"����wy��I?����Z�L7[ݤ�АŹ� ��i��g�>G�p�&�T���G]W��; Gw劥�.�Vȍf�hR6�vN/:�K�FX6)>X��Sߍ�M����&��+�N�l�n�d �y�������v;��nc�a���#á����I~��>*Q�Y?X)��yFr݄�3�,���c�����eJHz���	��\*���	��1Q��O����I��y�\\�_� �]��� i�:(��X���Iq��8���y[ e�>Bd�WI�;8����m���n;"C�m�j����p�6�: pU0=�n����wttJ���J���H'�p�Q�Q�^�T\΅'�M�Hp�"]G '8�1ν����-8�p���m����9i�E��!CvF����|�_9��*Gܐ��
��6��O�{?t̳h(��)�E��C&@�O�e-�@F�yX��O�Ԡ��2�K�����0�s,rk���O���y��o�u��i�ǒ١�@ՃrrU߂�%M���!)����Ѵ8O�㊏�q�&�2�\B���&�?���v%e���|m��v�T�`���Hׁ���PM"�u?rޖ�ELe��jjҠ;�6��A�=ri��n�ʓ��$`����S���p�z����������t��Uz؛�8O�Ň����	��ڟ�	�I��t���U6~U�᳕�B�w�x>i��F�|��r0�M��y���A���}�����W[�Wo)����M���� {K��Ҹ��V1�Z"��F��22!��l����HyY4�M=��{�1|u}�\O��呎�=�|B�	իKhDV���8������(�k4�
��,���,��`�*�:�ya�۔�<e�K�vv���������Fm�L��x�G�W\1���Wvqp�{�eoc��|�vve7�,�s0Ca5� �P#GG�H���'0[q�yw��� .��	�>�_K��x�`^[,�<?X���D<�1{ޜ[�(H��:-^��\:Ru&ڈ		��āA����/��px�ǹ���ȅ��>R���(��R>��3��'��y�bD��}���X�{�LL�(	t
%�	���t�2���[�}i&p���	�"  ��IDAT����"ou<�gg�*�=�P��,��=�ui0����SU@�]9d⊺�9�HC*m�	��k̸�g���ڀ���Q�uǵH]����K7�2؇/�8�At���GΛ2� :]q����<׋2���(o��Iޞ��n']2�N��r�M#gl��ۑl2�>Б���L��
_q��E������%�KC�hX�����sөy��I��U���X�e�]^_��sv#�f&L `�����	�u"��ۃ`����|L�,��n�����	B��Vm]gQ��,�� 8vT���X
͖od(��T��8�ex�	p�h�~�'gP:�i{��.�Q���X�n�0�Z@�ԇ���_c<�گ�j��w�1�9��u�4`>�`�w����m�so�ˎs�|�)�+Wf|a�c��ݸ��_�f�T�9�u��%��t�G��ɗ\5N�P�[g�Z�u�qFcr�(�8Vr�`�
�~���&})wB�� 8լS�3�۩�ϕ׶�vW���,��7��q�#�I/�#hpj�$�EY�����F<D�?˿(��Z>�/`�_�2�g&�l��J�'=r���>Z� �-mey�ڿ����p�w���z~g�����/��~����'�|�����
��*��Dk�[,��c��uB�`�"��ĥ�.�5C�	��n^uD9��.U��`eR�cٮ'2�
�\(8
�^��\f�@��z�5[ Ȅ����gY���.���
(��,���FA������8;L�8�v.�Oy��+?��n|�h�Ү��п�s落�zo$� �#`4�/�Ry�)`���r ��� 1@ο���>ȹ�(�0tWi���e���Yב1y;>�a�o��Y�N�A�v����C ��@x�]��!eA7W-�4&m	=�Sg�+����0�+�<)+��4ȁ8x.[ ��2�Y2�v蒖S��u� �>��ӱ�	�O�*4SAtխ�{P�mu겺�9S��µO��˦��g����ۅ�_F��ܓ%G�T��&0�cp��%8?�ć���,��MPv����7:���ݜ�Vh�q��r�{~賖E�]i���a)��쒵0����m}��-9L�n�+^�_�R��j^�e���N�#?�-W';���5�U3?/�#Y��^}�'\��L.<y��09��î��W�/\��>�򪨂�?2]ڸ�ؖ���f��\�F/�η�='�YZ�t��"��+~�I�{��d�n����^�c���uv�x� }�VvɃ�x�(���������@F��f����*��c�v?t��Cɛ�_�w��묇�7^}���s�_�5�$t�Πڜ7��5|�u��E� �.m����˄�9�B|���yp�cQ-���׮Y�%lܴ�u��� �n�X�,��B�x*��w~ی� �['�y�7��i��n�\h���ď��;o^�sgw��Ë/���'�z�_P�[��2xWF���O�v81Y�rt͸c�|���s`���b	�G����X'�3B%.|���j�NYC�<4�B�s~�ʫ�v`23�s�� P�_�YƧ��,�+��:�E���n��Y���^�zzg'q@u�
)R嫁���sĵ� �ygX�nud!࿍~��]��M���g:��,o(�*_Ǆ��a�7%���8���F��	4��U@�u1��6�@Q��b����^+e��ʊ���4�č�+�64�͘;-r��4�2���B��p�x!?��̔yX�Rf�ݠI�Vt����5p���K��N���NwF�n�8�8��u֟e�:3��=W�щG`1S�,���a�~��(�N͜�Z�}^z�@���2�7��eOi�gd��;ϓ��uݺ6��ϔ�����:M��.�`an}j�����b���k�3��#?�(O��q����~W� �Gnѩ���� փ������;��,��e�X!ٖ��W;X���;������6�ڦ�Y�߹s��N��s�Z8�<�Z2�\��}�Яոq�Wq�F��;��a��e�w���jN���_��&�If�G�7 Gh�_@ ���;���gH+;k>�D������$�����Q����lE���~5a5��k�۷m���:�u�]�'�T.�9�����������t$�������&ʞ>u�"ڻw���`���Kj{_��>��� [����U�1	�޼*,}A
�EN��?�~l���<����?8���I�6n�5_{��|��<��.��Y�O��=�L|n�=���˅�,�E &�[7oi�nVv��?��޳���W.��}����>�d�]VvQnU�B"����Rx��>N�/�4<+�� R;E�f��x\��.2C���M BCR/:{�W´�hŠ�G��c#�x�$fZ[�mU
OT2�{kX����"����#��S��`�!6�Y�8�?y�o���霕�����_�N;��	�b�u��5����Uw�����,-y����n}����r]8��q�Nx)qV�7W�뺷|�?���'_sl�xT]^����Ƞv���A~��\,����N�9n�ڌ�S��>6���AY�C+�%#mK��Í��rZ��j{&0��+���V�	V;_m�}�:��CGh[�z@�./\�d��/�PQϳ
��c|X1�\���4����ڃ�e��ѵ~�l����2&;=�&�	m	T� ;�C&�)'��s%�E�TO_�S�_��:*�wIa����W��n�qn�X�NS\N@h���<�����>�j�>}��ݖC�Q7�����:�����]�mNPt�z3័<���'Oőn�tJ��pE5���=��q��z�������sva�xHw�W�]ɗ�zB?��'�c��ҥ9�N.(׀�`e70���$�sl=g����݉uθ�S���>�M�ص�M�4���ė��G�s�jE�d;Ҳ��G��[k�⇃%�?l=��CVPe�Y�o�_0�+�#Ttr��-A�vU����q��*c2��8n|�����eeWN/�{0noܰqعs�p��k�a����M��l�/y��{�vP���~d8�����s��sϛU�Uxx���'�����c���=����cڙ8��}���8�m/���q�� �PW���;tlKԶ�q�W�G�6�M�h�Y��5�@��8�T��<�Y�;�Dp(�yx�c/:o]�k��Py�E�l߲u��ee7����]޷o����W�g�}~x��O���ݱ3|�_�Y�f<�� 9��k F����_R����h�8 -�,��ī$�� N�K(�j)�$�c+��]����P��1��m"uxp�x��\��d7���r��g~�3~�Ӂ��ïn���{>0|�����EAE�r�	XfpR�HK������ ܓ'N���\��騼f�Qڎ#��uYE˿���y�Ʃ��P4�N�*[[��XVʆ,��pL�o@��tp�\A�$���K���)�v�ӆ�����V�v��9�r��;/2m��6ӑ@�l1�P�
�I�U2��i+�����πp-#�jLD�}�G�u��?�"�e��^�Rv��x�+�{�y��j��aaEG����*�M�
�5�}f��3�{������᠌���N�9;�y���w����I^S�� 3������t1����kgW2CN<�<6�t�'2ia	D�e)�(^�����r�	����g�F�\E�6�y� ׳Gg���=u�$����,8��1��Y��۟ ���@�f����z�v�^�6y�Φ~��&�<�q�d�f}\ =�����9e�uU1.�C:d�\�Ȁc�jǱ���<P���.�n��a�*��+��ɇ/�O���~���[4�s�2橬�/k�n�Y�Z�}�ȝU�ZJ�~k��L[c�1�c���i_xMYi�	"B����Wl�_�W��0#?�e�c_�^��5(Ђo�#�����u�珣�p���.�>3�_�m�8E�Z�z��G7�g����_-[�6�M�6�6v���ާ���r���q���_��/��7��N��'��o��w���/Ȇה���x�)`��M�U;��]�������<:|�[�^޽{8.:8� ���@璂��zr~�d�_�y�8c~6Ƣt��[�� tV����"b��O�3c۷�F'6�̡]�h�0���>��x�z�`�-^b/��|�K�B��m۷l�[����ĞW.���s��h�������/�:��{v�H��w`*SWe�e��1��q�W�NR�&��dA)��I�2Q_�v��tr�;�_���� ���QG����҄O�q\.��������r�]w��/��W�v�~yxG���7�2�.��*G����L
ǡ�5�L����G�<�ۛ8/��9=����Q6���S��=|C��QsK�:A.�;+��!OV����4 �V��i �Ԓ�z�2�'������N}A:���Y�z����c�K��+ �;�M�B�E�l�K�q����ņM�<#t��0�Kk8��� ���(PD�|�Sx���m!��v��� ��I�<�����e7n�4�Kڏ���>|��O>9�!���C���~�9ZguL���7y�Md��68��W�?MHS�_��r=��K���i��O񭯪�j�3K��?��r4/}�ԝ�\��I�\������5���`�d�t�1�Z����� �����_v%x���u�&ib��=T;U|l�\&]�/����:Z�c��[��_���S�L���+����[����q>Ç�����Z�ގ ������W�W�M6��XE>d��l��u�p���w����(͋�1c��
�[kt˸���ڿ�{0�¦�0��Dٺ(q@>��@�lәlw_~9HU�Ia���̝Rw�pxY���ݲu���G�#���~�v���8�;�V|7l�s�%�ԇm�-<u&O��Z-�{��d����W��}���sÁ��o��t������y���_�O~��k���ry��[v�,:d�`[!Rǌ��{hr�U��� v=�'���˘��N��I�s4�@k��:IU'�a����v��5}�K+W����S���)�b����W�opd���������}\�{v=hU7]��C�G��V	bQ�	�Ez��(���5��R���al)��^����8�P���S��Oi��W]�����|$�r�ObcJg��=��3������s�/����\}�5���8Ǐ���_:B�_	�R2dI�&�V�2��3�b�mj\n_�_�P�;���U�88��=�Z~�#�L�d�G�p�|?&��F��t���ӱ/ߩ���Pr\�.��I�o0��ׁ4�[�ވ�h�L2"~����³�6��W�?�.����l]��?���'0��Htkp �Q�5��(�L�@�2��pPF�[\t����,^ח�d՞'sW[�mu�*������L<8|�+_^ݳwxu���O>a�#��^hF�U�P+�E1m~s~����ˁ�X S<ǥ8���!��_���#�ԛM�����U}}�i��tpЕ��QI��Kl<(���3~��U9�)��5�]���C�����\gx��q��[t:��$�y(��
\�0�����͋Ꮖ���2�Aw3u����h��q������'�AsAz��E�u�1��
؀82���qF8����	�f�!.��~e<Q�H���w��v,G���"p��~��%��w�^	��X�:՟|��<y�az>�>��
��8�*?�n�㜲H�~]���{���G��e�(�$,v���
]����,6�-p�{�s5�;v���nި����9�������m�ׯ���94��_����w^x�E�����y���|���vvU���3d4�/�E��"����˧�+�C�͒o���5�q�	Z}#۵k�;�2=?�*z��]+���s�@��.�M9��Uc��:����c�ٽ�����pv_{m���+{����]f�ƀA��e��-Ɨ�"�(2��a<'�W�I �>��T٤q�"D����s=�"�6��E[e��Af<p�F���M�!0
�@�v\�c�����_�;gx�W�����6l�-
�U�}r.Μ:m�D��]��uS���+��q"y��ꋓ�K&��A���ŀ%����>Wz�P~@����\���%��}�&ظa��4{���o^[4��4�ʥ�Xm���;wV'\�YWE�yLOqt:��|tv�ፎ'@��O��'�PN�k�uT~�qԭ�.ޫ,�˸S%�ǙӐ9�'Ʒ��a��5�-{��\}����n�}�H|�_�y���ݻ�g�N4�O�*�8~�c�.^R��[�'R@�/�,�a��g�|����c���P�y�P�F��K\��tp�Z���$�:O�]�sΖ�˥���x�<⮲��v&��@�κ,�@tX��滎&�=�-,���$�������^խK�������L�E��߇�;+]������k�/����"X����H[�>k?R�� M���!�W��t2��n��fؙP>�p�saz��ؙ�_��A����a;(C�Fh/�eS�É�9�a��R�A�C\�n ���/u�1}G��
n�MlkV/	�?��V�m�u��%�z�{��+{����0~�b��Mù��*}��e�V?W��fl���=��۸i���u�굗�>����3��?�����%ȩ=
�7�:��'�^f�B]�uN�m$��B�돽h���	�]������$����ӧO�X�(��8���b������=�ᘨǶЦ�/}(3���=�ʓ����p���_�$A�JLP�.{v�}�E;���?��>ofk�sv������)�X��l%+��?+��;��S��G�!eUA��,eU|�< �1i,�t0��)��V݉[G��\_��7o�<�y�]�/��/x����[y�o�n\�N���CÛǎ��~d^J�S�[��:����e���r`�����*'�m����:6TђCG�h8���f���3����&wЧ[�>Pf��D��@�gw�#�4� �+�:"u��:/��nM��3+��8|@�q�ky\��wsv����/-�< {��Y@Z^х�)Cq�-��i�s������L~��2q��%]�n�����p�}��v�o�8p`�����{�{fx��W����^a��;6��7���7��Q]�l�9��U�Y�p<ǥ8}�⭎����@0WmRy��<�䫼S>H$M:0&+Ҵ[��P�g2�b��tg{�66 OW:Y���%�[g��q�x����j]nģ����m�7��E���������(\��K�7���#�0Bц��R���y��h����tzC�ҧE��COcٲ�@d̖��tݧ��7t�������b?*���6�.�O�.pJvEw�V�3��d(v��MY\��![ݺb�K��h9gNk%@�Vge��"I�>x��R'�z2�1��>����t���#�\�����#�8��$w�y�!�e�f�z9��9��:�S�G�)��x�w�sV圓�zֶ�؛o�L�y3D�L݇_h�<�6�@��Sz*���`�ȇª1�5�ë:j���ڕ,��O�7~�No?����|I�:��vt�#2VJ�U��G�,��n��z����a���ݶ�ٽ�[��.�|TA0��.s�z�)��
CQ\Ɖ|�г�������⒮�4L�a��Q%�) �t����%�O���4��L�AG�d�Ź��c�p��h\����
G�΂���V)
�׾�Z15Y�N�F?��\���.��)�O��[�i��
*��<1d�|����×��eEgsRx�����U�$c ��b��:�Z�\��|�E9GӤ]i"�#;����P2��fh��m4/��U��ǀ8�iD?�^��N��K
tZO�<�4�ґ���~���G�^�o<Vy-C���Hi3�c��9:�ӊ�jV�}���&�)��hO�8w6��n�=c�Q��l��m���=A���jV�h ���	��$;�E���ǻ0�˩��=Ct�����=��p*���R��ߕ�'R�N����V?G	�ߋ�c�M�Sx� KO�cx�(0��;�U���,ǵ����!w#(ZS(��l��|��r�>`(>9UH/�8O��'�u��*�?l�X�BU��e�n�M��C����~�������qEÁ2�cB�_5W�!<�����P�����5����1���v�ӟ���Kǝ�@.L� ��RdKm�tEU��|7%������Ե�ʶ2� N����#�{�u~�-�r'�����c��#����?�˶1�x�䑣<Cqpxm�>o1;z����㍬��^�M
��5�7��aæa���~0��uê�k䘮V����*x��g|��;�7m�bZ�Ma�����퀢��?�t��@��C�,������]s�۳���,���dt�'��%gU�`[�t��	e?�_уT��|N��l��:@$�uD�	P�|�=���]:�F�}���L��e��_����+;sI]q��'��n��}ʃ&�n�%/����'d�
4u&x>D�z��ɔ���9eh�x��%�#�?s��p������1G^�tNNG��t��y�R�r/�Ki8�#u6��T��l� s,cO�i#;�C� �`uFN���D���(?�<(�o���|���Q�:�y��C�j�p+�kh�S�-�ZV"�~L��0q�]���('|�iQu0����5�ė)}�˗x��C�/�2��L:�a,'z��jZB���v��W���9�m����S?�i�:A�N��ɣ�Pu� +4pǆ/Յ��<V+�#2ƫW�6�ߐ�6��Z>T�^Fh�â�@{{����K��JF����^�3|#���V�'TS��K��L��s:��Ta��@������k��+�G�u�a��|�0��.�X&M:�%�#Y�O2Y#yq-�:r'!-OD��d[L�#+++�N}n'�F㡤�A�#9IcŬ�K��;D&r���?�ACɣ�����ƌ�T����GC��8����`gg�g ��8�8���(Iq���O�,�[�q��D��MR�T���J�gqI�YhA<-�C\�h�V� ��:�����d��=dƫ�X!���G��Z
�6���\�K�p=�בx/@�Ƴ��u�nc[4�~����\O�6g���* ����fO�˥��B�5�:����3���!a%Tc���yK��.W��Z�p�J�_9�|��M�7������Maݺ5�j�I�º�k���z�;��;w[�m6o�:l�~Ű��+�-�^+�����y]��t������+V���y�Z6E<`��C1���7�
��o�x���V�m[� �|��K4�.���e��ԙS�����xN�#�j��q�Q+T�
���Rt��䲂M~V�`^���M����;$�.-�Ѫ6��^�R�����@)d��z�\\Z0c�e�/ a/�х�tʤ�!N�\���<�z}'fe�a�^ѷ̤Y4�K�N�f��
�h�Y�=�h��Ij��=��"���f �	�N1W�Ŕ{��g(�|+Ɓ��x��y������Gʾ��^c�I�3�v7���T2�g��քG�Y>�r#����A:�e���,�v���������/r]ћ^�f�_H^��Vw�0}�_	�%�l�U����A���T�\G���׷��V%O�5��ͨW9l^e��e�UA�K�C �[�$�6�
kF;�d�k2��Ȣd&LLv�M�|/��^����5: �Pc�L���P���� ^�.�֗����Q@,��Y`Q�?Gx>?P��2ae��y_�I�q��U�_V�Z�~��G�^6^��q�葓6���1�8�=��a�@|�Li#0���u}?�̥����ß�y����7��G��7饏8�ͱ�D��/�v��ЩB��y9/P.:໰+��p���UW]5��q���F�|����r�Q��fk�zX�5�����^ .c��gM�ꃿ�VV�Yh���l�td��q��*����1oL�R�X�)�[�+t��S�bzU!� c����p�q��<LqI�ѽ��h���%]L+�V����f3�:;\�`@�z�¹ʚ@t��M0��6��� 2ϓ�R�}�~@OϫV����rGЩ%Ѣ8�����*/�ܵG�e�����\L� �����\z����+��5f�)��X�CK��'����m�?��>��O?��?9�������?��~���o���G6��э���E�p�O꼮��\��M�v=�%@9���M�Ss�����2/Z���kʓ|�q���r�*?y��F�Ae������;�+��ҁ�[��a�ի8��������4_ۖ��29� _0^��n����"�8����&��F�s=Fܖ�^��B�ב�h�z��R,UyJ�v����O�ottn:���3�{���2����gCC:,͓ �#��0蟇g�������e�Bϧ���-'�|5n��5����m��y�nG���xn�Bs��@� ��,�K��ǅ���p�� ����_�X�8�|3�'��\��'mQAQc )���
=���ud,�-�tp��A$F�f\�0��nq7Г� ���4$(#��O�wt���qi�ē� �(�S��.�O��S����D>P}�t��+[$9p�`��Xf	�P�'�y��O%�
=�e:�sU(���ڀm������"H<t��GY���˷�P
T��y�6����0��U�(Ĵʓ��p�&߸��:<0�#/�������[[U�f�8]�POw�v��K�S^ɢ��R����ѝк4`>.!�z
qzkoٲ����T(�X��˅�ֽ ��.%�Sն�	��R�*<���@��Л��V��?��G�����~�gv�����z��_���������Gy�3~�:ѿI������ ��^3��m���7�� |��g��Ӛs��<`��E80I����ǘc����P��|l޴E��a�;�k��n���[�;n�s���ۇ[n�u�Y�7�x�p�u�;��5��*;��jd��/.�ّ@��b�&���LZ#VTx5�'T �#tzY��m}�����k��PMS�z�
v�I�����J�a;���3�Bd0�<-���[�q�
�<f��Ƴs݃Y�.�*O������#R��������I�(�m&;����͸��� ׵	ފ�>�x�Ϝ
���-kM�Ls]!� r�c�H&��ɧ�q��k�ݖ~	r�>f�C�h卭q��]*4����h+��7�C���.3c�I���fC9���:#`�*�)�hM^��G�.u�A��h�e,�Qn�狀�3�"�m�� ���t7���2tJKr�I YPV��0m�>o��
U)K�cp��T�����e��"��c�<� ���I��E�GC��NP請g�s�Ӯ8�7�0���Ýw�9�b�'O�s�gϜ�R`'���;3�U�y�{�g:N�=��\xO Ihs��t�АZ��%�>6Pͱ�o�0�46�Y�s!����*R�����E���AW��a�	d(�wuz��A�[��\s�?��d���`�p�z��c����|������U;�0�>!*!z�'�}������H�5�F���\X��d>,���d��J��l�2l۾}�"�u�Z��ᰬ֭�0�x�MÇ?����O|rx�ᇇ����p��~�ç?�C�O��O����'>�qٕEc˰a����=h]N�T֌�X e�����	f��,Gz�#���"�B>�څ�(��P���>�&'mr�k���d�6GDav���`�_����x�1,��:��L����ʸHX��N1�k�i;4�U�8_u<|$�$�XFy��nȇ�c�- ���������2����rA
�a�Y%�/ׅ���D:���� �`��� ���qgC/sx��V�m��zq��
�-����Q���ױ�x� �{��L�p��'�M�������Q雎q����瘯�p�ۃ��7(�y�]���ن8��,�Y0~É�c�CK���7�pR��c���$(͕q�h�Tl>�����N�����Txh/�3 �E��w��;�k��λ�];w�������޸`�5�`�Re���c�O|�??΄gyL�ꓺBo�	~���:��?�v�.=��x�P's@����<���#�ƙ%���s���q�B�/'����-/�t�@�0�ur�q�s��VF_��И��E�ra����&�R���Շ�&��W�St�ƭM�b�n�m���%ǭ[��V��������ÿ���~����7�a��}�h���JF^��B@2}Ŗ	������`ę�U��/��{���(;�EYHo<ҧ�0��/6��_z���������]��:��ɓ�E����[n����p�&Ɨ_�j8u��p�ț��o�)���}��Ï|d����[�=��;l۶]��ی�M���h��o����p��9;?��i��$�� MtƲ�D ��۞ByZ(yC�Bt8�:d ϝlB��i���Zc����WT)�����X4���I�d��C?�P&I��Lυ1��C�5��X.~�RGV�<N�0���>ǎ��>�3�
�A�J�s����B;�����[3�(w��;����Ǖ������2��Ds�
�ָ�:bY+Xg��OtlBަж��`4�����������
�l������AZc�u��5(P7ױ�!/�ʫ��c�9P�y:v��(�\�$�F�<��$��:^რ_���;W��qd!�#kGSzT���o������F<��'!��kRy`;�0������vIY9݌Oy���m�Q��+��MѮ���P���ˋ�Q(f�Ev@����tr���Lb�(�ӑ��`�#L�-��n]/���	1��,r�VDB��β?_N�\���8N�_�����u4 2�hVNC�H�G�q6tb�G�W;�m�d�J�6^B��Vh|Tw�39�0��||� ����Ǳ_F��y�p�۹�CL�(�	�܎�3쵸��<6K����v�����.:�U�=x�R��-�'�(u׋ i��WDP�K|�ѵy�#2�{8��8'��ҋ/_�����������_�ʗ�*0�W����d9��E�����m�?f�wD⌥~��̱[����?�ɣ�������3(����B�����S��ec���2pV��߾r�7����ÕW�n����k�W�ȑP�;�3R6��9Ѐ;>�z�U��G>��ᦛn�S��C�|�xf�N���TW��w(�	R��2�c/*��x��a�5��EPy�i�b3i���&L�A9��ji�^[D�3�`�� ����E�����O����q@��P��LBʤtd�ݞ�7g.�;�:�����Gx� ��|\�Q9�'��6p[[;p�8|eB��6t��rHz��<(�k���y¯���G�G���-���N��:�����'�fs�L7������~�HU��U�1H�>��Pq>W(��յ��tȃ�r=$��� ����e������/&�$r*��jmW�Z���p���t���B�����2��@�E�b���|��[Z\w�=l��|(�gk�X	�MH��0d��\2�jǚ�KeA%_�g
b+IJ_`�VE *f��3�����t����IZ|43�P���OD����-���[�f��LiΡK�.�WY��&�aL���DϠ�'u�r��hp7��#�DCX���G�  �2����_���`��9��$������2W�,���R�I����PX��l�aAN�+�熿�2�z�A��Mݜk�]�D�����-(V��z�uY�ˇ'v���[q��w>b�&#�Int��T�W�(��z���u�	�{c2�z^��դ�/$�Y���C�Ňm�Aap�ݚ����lAV�xJ�}�<��6�W_�3���n�}�����џ~�������7�4��/���_�������w�q�ߗv������ʱ�P(۷��m��N:� ����6��ǃ0���3��Y�|�'�V���E��)�3�WY����6��nЖ�o�_��)��QA�mGq�I�p�ZD;���&+��u��I�!g����e�0'��%So�c�g��ů�-}b��1!]%�CVѵ�Ff��]�������� d�����^s`GH2B&ȂOǲb�;P�&(J��$�,e�+���.� XZ=s���������0�mY6,�t��z�
ٕ����>���?|���i��A�B���d��<��TrN��!ۡ�c'���mym�(�zK����R���>o��g���~�璙��\���B��K� >��n*�ª�Ԟ���������/�y���_����/6S�0Q�FF:hqf	Ɩ��*��N�:���B&\s_���.EZ{.�
��?�(�iXt�q�A��{�>��O7�t������yI4��m۷�P�ౣG��{��%��O}�'-�I�����Q'f���y�o��f`i��>�e_��,Y%���0����e�B��CO�3��/N������p�V�H�����!X�jn�Y>����ό���Z����x�!�ˆO}������p�M�Qa���^zi��~ax�ɧ�j��g��z��������+{^�ӸR���?������������{�
\�O���E*_�_ ����ΗȤ]��(y��6��G����w9:�Dr���俍5{"���+��'�����Rn����^ɒ�j9�칽�
ޛy�pŎ2�y��f��5#M��<�O����/<;��#���7}w��[lI��g��C��#˖�J��xUȃU��b8����4�h�-���z
q⽰��oF�ʏ�6?�ŎV;�V� ����9[lp���4;��������ک�<��ҫ�8f8��Ϝ�Q{cC��]r]Nx&}Dg��R�O�4��ȫ�C���4'Y1قW�0ｶ>6��W��FG׭���ki'��~❠x�����z|mmp��CҽW��^2㫌�����s��އڃ�(�����DS�]���
�@(��n�iϜ�0B������ȏ�*�+������Tr�f����mh�6�y����O�Ψ3�Y2�$�s��f�i�K�A��ڤ`�F�8'�ȉG�F�[I�K�J���_r�����ŗ^�y�{�I������Ё��	;�c{�;�?����� �^��I|���^����CL����$���"�lCϓ�e�E�r�I����d�G����}װO����Wqv_x��n>��+i�J�͈-C�yt^}~b�a!?��Q�|ꑶ�M�,�6B�Ĝ��$����A��o���Ly�e�P�1@���'���0lݲE3�m�����-[7�FA��=x��mj�@�Q�O����̱a�N�G����qq`�yr-��R��G������{-S�-�,(��.a9�g��h;߂v ��-c~��2_f�8�}{���2`t{X��~��n��f;`���>���駟�JO�5Ҙ��ym���~�C����/]=�=�����p�9�c�KG1���_��%�P��|����� G���2��s;[��/�ɉ�}֎8�����J!��/yg�{��~���⨭��X��2�A��8���$�B��_��B;����áC��Ç_��yT��i�i|C�P'�t	u�)rA�Ll�-��q6q�(����Jl ���Vu��J�@ɽ�����]l�o]���0P1x�o;4��ƛ�����x�A~���l�ͯ@{t+J��>9��ݫA��a��C�a8�M,g����쮜yH�M��B���>�U�'�Pή�a��^Ƙ-[���r�p��*��
���ȓ8>V@�?�ޛj�6��͵�.x,��G7��<��s�_��_��x��(\�c��	��m�?N�I����UZ�p�|tlJ�����T� �O(��q��@�}��]������vԄ����%���&G���(k޹[��J�g�dhs����q-|~:�?U���s�ٌ�M`R�ZG�쪝�C<�lgW��:}jx��g�yF��	�a��Om�~m�]3y(����G�4{qB��٥_��ޱm\/|�s�>����~@%ӳL���,�[4~�	|����p�]rv�^�ٕ3��ս��/�<|����|���J��> �ʸ
��!W�f������uL~Bp�W����q���(�\J*:�z�+�-��1�'8�~Vt�8�S��>���;��o�>�9�V��γv�h��9,��g8x�ov��%���1�����*��@�s\s�\˾��e@��[;�"�qa9=��2�ز̂"�������r:�η�Hq|�Ƙ�̗�6v�ހ�g���~��7k��ћo��՚�}�s�pvYm�+=8��>����G��G>�Y�?�j��?����~���#G��`�>功yP�����٭�\�Gkr��P�"ݷ��&� _���g~Eϊ�N�nd?"�����b��ڵr�����^�Ş�5%;2*��j�{K}���iЃ/��?"q�����5{1OzՅo�=|ط���`u����۽t���Fq��#_�c��o�Q����Y�J"�b�0�{�1 2N ���8��S÷3ͪ/�dɾQ� ��&?�#?2|���|�A����&gwi����x��8�{�ԏ�i�o?�������}���c��v��9�����p#2hWVvqnXmf0���뇻�[��S�}��g���˜�GqFݦ���5Rԡ��g7+�)�&��o۶mx��� 1@ο�?��?~�7�_��'-�]�8	{�Y�l�Y}�t���^�^�C��]�a����{Q��4�m�k:?�.�8�N`�+�
�7�A��/�r�crvM`��]o�H�o������}�0%d�KG@����f�[�H�pv_�����f?��4	,�;�M]����� ���02ɤ6�Q���*��m��S�+N1l�f�6��/�7V�>Q�ټi��]�i���ٽ��;���������ٻ�59��/�����O_��W���­F�Q�x����F�-���%OXI�.��o��[�&�(!�U�OE��͓����9p���ѳ3]C�5;��7���J���/��Sq�m�ۯ�N�x0b/$��+d<(�СC����o�6��i) )�M�&4Em�\���hPGd�\s��Bwj�X�I�\$��⁹bg�����(�m��.�E�+�Y;�30��ў�E��L]B�D�Oh�߅|����m,��<0]Pz]�*!���~������n��ˠȶ�����U�~A��1����=������� �z�㎻��O��u��k���/|a8&G |���
qf�g�/}h9��E}j�:_�F�:�4&�?�fp�V�G���+���8u�����0�.O�{ P�Y���r�m	labe���Q��Q�a	��$���ى+�5ʏc�������ɧ���V�}m�WtϜ�5�	������7���L�׬�sM]��8�8�o�}ֶm���� �M�C<�6:�ul��98@{�� 4����%�Wd��c�Kx�m5�͟���~�~j���{e7���4XId�P�,O���N*`��_c3��	FmE��w��m����W�\O��~��~�H�8a���d�����Pg�׻�6�,�+�H�2q<�x�wX�ʹ�2�����'?�k��q�.<�c\v+?m���Z�3��`�������}�����'ȑ���\�wz�c*�s����w�Bp��|	 }|�%�h'$�	�cd
P_�i�����|�/xE�*��s��E�G�NP��K�����*g�M��8Ѡ^����r���G�"w�"�(5i��6o���3���`��Wy/S:����y�|��g|��c
����@�Ђ��C��h,ٰ~���_S&���QwꀜY]F��Kݰ���¦�/�\�!c䍞��~S:����������{������]Vv_ٳoxᥗ�'�|r�җ�4<�\�]d� K�T����X�:5n ��g�LG��C�(��Z.-���X�"B|:w��U��2�s'#�B�p�B����4[�̮�@�THce��~�G�*Vvq���g�a��UW�p!��|_�x��<];�H9(g��H�;�i�tc�׃e:a�0N�6%��|�4�4���=T�	�_�[�y��{Yn�+�[����G���%^�^�AȠN�ѹ�`�:�0k�n� d0�D��?�����>0\s�u�J�{v��{x��g��G��>��0F{^�3�Ќ����?�S�������_���@�g��ն�Q�Y��yFϗ�m�&G+׽<9���9:��:;�	��h2��w$��-(j�e )gW�\d���Y8�>̀�-�m[��8� �.\�^��jrf��Υg^ȟo�_{��~+��<��ja&�������^~�E���;2�v�O{������KtL��K~�� C��L��o�U�F�Q��BN���S����F��J��&���Ǿ�H�'��N�W�tD����_?��?2�z��!�ڷ;��fE���Y?\ɤ�� k�RL�)x�~Mi�c�������^7/�U�C� S�0�gt�yg���w�=���%�J�����,�����CnA�����|�-�m��f�a�k�i���2�0�����ns�)��"��{�ʸ#G��m
����}��>3���~��?�g���Ʉ7X�c�};�F�x,-�� ;W:���7��s��<V9���I�N�j�������:}�i�v>]7��x��v
��(>�W��M����S�)�r�e�ێ.�B�_�I2�^qɄ��U�œ��{x"E5]dơ	ϯ�x���3��]	�N���������mO�C�mQ�yA�Li��Ek5q�>���gѥ
�Sll�w��(�4�BdO?~]�S�k��0��q����6�w��������l�E8�����|j���@�YR5{�4F;�P�6ʺ��3��L�PZRn`TH�уg��!�_J5?���n%WG��Y�����(�STH�����ď��f߷���*��1K�z�UÕ�`j߁}^�8�����	r��]���ڋ�ݮ����%8g(�8N�`LUT�;u���L��<=9�#M�(�\>�ϧ3��Q�Q�^&>rs�_\{��h��֎�mQf�6������8����]Vy���^���������@pC���S�X�e��?�������Gv*00e��Z��g^�7�L�Y��=��[�������<����J��c����!�ewz^�Y���S�E繎í����~��������+`���S&k֭�VV�i��k����췤�so���TD9-y�RO��Ī��ԩ���@�;E�Ic[�9A �E��%��F���2��%ے��iT�OP��k �t���V�S�J�oC��xc ��qx�#�8�����tLȸ�遐�Sr �+�����|����A���my�$[;h{) K�c�Ԫ]��貒J%#t�%���,�O琺�>d(CǱ���W^y�������g�<ȁղU���j9�rH�X����e��D��'��(r8\8�[7o~�o�-o!a�_��>�.�����"k񗺄oج�Fju�*���~B?�.���ߩ�e�k��Z9�?���?��'������0�L<�+gW�267�08�:�!uߋ��}=P����z�	 �U��R��_� ���7tή�I-�7YPt}�ܾ�\���ȃ���8���=������z�`E��E�K�]9���$˦-�?i�3~sUsz̓p6m��mV��ar��˹���hc�]�Yo\�;����rv�G����A�@'f�|���ሎt��_~��L��$,�ƈ<�0Ak4�+�oH�k�;!A�_q�$7e�Ze�0=�uM�g��NC�h��P��@�>���P~�vHz�PדK�А٫Ċ(\��=w��*x���5�0��ׯ3E^�ĭ����G����N0�"�ַ�떁�q����#�'�zY܋ �ч�QƊN�g��q*˘��\(}\D�Eu�q�@rS�����q���s�N�ã�r[���<���ȱ�7��A�� �҈q��ڲe���O}Zz|v������9Yy����9 ���2�;O�K�#]��ա��B���q6�vt�Wq��e$����#+�;��9*,�o�۲e�_�S����&�vÆR>����>��?����;���hV̯����kv�\s��	��6oTI���A���˪���3�.ߖ���1Խr��	y�,��L|�A:6���!i��>�0U=�\��Q.�z�f�s ������b�[��ox�#����_���9��*�}�}V�4��� ���NV�3!ɤd˖-r"��M$;v���q�pŎ+��v�-�1����[����ܯӄ�=Y��1_���ߐ@����s!76��|�e�M�f���N8����t&U�ǉBF|���Tz��
������ʑ���8?�LrX!�EnL�p�W
�ƛon��6���?�s���
�C��)˪�0ߦ�O8�C_�`�'r�Ex`��B���6.2��:��K ��kѷ䵻�t��|��d�O�J_1
�Z��\�#A�6�x�n��|�����ёr�쑮ϱ��rP��_��[��h�2��>�V�����(�*(�6�|�H>�F���뜳\�0���rZoE�;&(�H=�Q�\&��Y�-N��z�ȉ�[;�����+�ܡ�Nkd{O ��UA���\������d蹱{���'g3�o������;
2����b�r����L(u04���	�ߊՂ���k �】'��Ձ,�ޗ�y:7�].,�*�K�OХϐ����`�gw!�Ә	�ׂ�T�{�%����!8�v��
��ګ~�nv?�-2�����^�k��=�_�(:���2 f����@G��5���z,깽��0�R�b��X悓8�|�AÙ�j�%��^�Ѯ�eG ���*����?���22�I�/�@��K�ଋs��h��˙`��?mO k2���+o��f�0|��{�{�{��;���S�ۆ�o�y����]W��mz^w�ͷ(�6�}��w�y�p���y�$�[(8�����A�$�IN���h1&򹅚��@Zu7����>���-��֎�} �8 � �>��È��q�t[=�XE�m^^Ƿ��t��:'0 ������rpۑ�8�l=ۺ}�'w|♶�@Nq9�,h�S�s�;�����J�� �T �*9ӻv��I�u�*h��D��A�[n%�:�z���o�D	}���ۇ믻^e^9�c~�7
�����aǗIm��y��pƩ'i��������Y�+�j��d��c!ힶ��+��p��-�,(ee� �)I��H��>��[�H��h�I/^[�u-k�zW ,�r~�-i�F�ɥ�0oX���w��V�KP��+	��X��U�2�$������|,�Y������j._��y%[�NT^�'�8�<�R[�̣P'�	u]�V@�;�ވ�T9)��]$�x3�1@S���Ra9�ѝO`�mtRZp���p� �"(W��ep���7%ki�a��ķ"�?N3�8ƪS�`�?։D���Y����c
��$۹��E����B��/�������8�h_����|��hT�宁�?����8u�t\u���ز�Ŋ%�A�d�s}�O�Y���o�������#�v_~��ĥ��d[� �ze�� 3 �Ճ7)��-���M
֬��	ܞ��6�|���S��u_T�A�m۶6��a��mݍr��۷m�n��L8Vy����>���=�����l���`�=0X�s�|�m�6��U@p�nq�pf�w���m��|J��̊	�*(�g���5[7I�ޔ>���|+ڤ3�q,|���ڇm ȩd᜽�ܵ`��<��l�<p��I
��Ā�
[=(��Ia�E&H�E��P:������pL��\�\�p]�Oiy���VpY�ݲ�o4�#=�&�f�UW�v(="�+�-����k�Q4q|w]}�p-δ�c��N���۷�U�Mޓ���f�f�e�FD�4���0a��!8�ic{!���~-mEh�lrJ�'i׌�%�)�,��O�tnh��_'y�&�|R.G��Ї�ׂ��0ў�TaDǏ��{Do���z�����"[uD�ɩ//@[�P�;CW�r;��9��!��:�y��K�L>��Wj�J�����m������d�C+/�g��:���wЖ���a�k���^~%��ʟ�UE4�Y�yPx fZǞ�|Q�$t%��_h��d�)�D;�����A��I�������[�h�d�=�PR�W�:角M��h��L�i#��ݰ~��ٟ��f�7��n��[3�~���7d��8�8����+��_?<����J�o�Q*"Z>�6����P����[Θ��r�ݕ5fx���
�:|>W6�=~A������#3&X{��<�P�pD�8A��\�q�tZ�����"�W?8�<��0��g����n��Fƫ���OO?����������|�oc�1�)���<��pV����7�t�����?�*��������v��\b��MN#��JΫ-����}�]��#Ex僴�>��i@��Wߩ��y�I�����5k�y%�[n��u����w�z�����+�l����u�D�2���3�s�U^����ku�ӷķn�b�����x�`���r���F�p�n�=��v�~�<x���ྭ����ls`��+�w�^��d�۪8��lpxg�m��D6��E:�2y�c��#�NǴ}RDC��X0 ��K�%[���u�p�jb��3�K��K�<������?pyl�` +�۷��V �.�Ĥ��UY���G���b��r�x�	﫦]1����k�lU׮�)J�yG���$3�:�)ԝ��i{A�LON/MF��p��fNoڼ������q��u��z�;jo��;zl8}�-��+�f��-��c�[��j�#����=	c��k{_N�:)>ŔێZfO1~�,��y�,��2Ѣ]�����l�[D7B����M�(\	�>ӵ���'�w�t�k����*���S�qp��,�O�����|��+�+�w_c�ZM�I�.�Ť^GT9�no����� 洱�<�v����b�����yn�>�8^���%Ǉݯ���x��O��[�����5c���~y�m ���,�\or+�����'o�Y����5V�K`ڳ{��{vy��؛Ǉ#G������~���4PP1$��T2�5OK�8w*��>�Ց
����B����O��>�t�I�+�΀Y���Ջ�Vf��Є��B�NJn�~[ޱ�L�,oJ�<��30y���yK��wq��I`�K�m>���@|���N+��냱9)�����ł�^��x��<�`I\;YR���Hiz���&���{,�o
�� ��V)+A~-�+�믿1<��cޓϠN�3n>��ӯ�f� ?���8�/���_Y�~�'2B����X	�0ɿ;pN�>������)4 �d4��z�k���4iݹs�W Ycŕ�U���ȷ4`�={dy��O-�%�{dhY�ñ�&���2��(�lu��l�g�0+��cb���&퍦���( �q�h�qk!{���6cK��c���)-�ױx��'�©��Ը���#�<NS@n�`�&8l_��䴞�8H���{����YI�z��~��ᑇ>�wm�v�m�m���7��'z��s�?��c���>�$�8R�9ɉ�'���s�L�I�_y֎��e�p�nq��&>�`	�-�2x�.��#�6syjK���x�W4	�P鹞�D�e��ᮻ�~��x���	�ӎ/�%�ǵ�];�p���6	�; �=I�"y��/��y+�-��͸뮻�������j��xn9�J��#hk3t�t��}��������4��9�<�W����Թ�[�q���-��n���z�v�u0�t`��1�uI��e�@�L ����W�5}@a��m�ߔ�m%�!�Hq$�>���]��8_B+~OM�b�l�ao,�f����+ Tz�e��tvl97̈́�W|�ʤ���Vi�Β��i+_c�l��]R��{��ҘǛk2.���b�3A_HA�☗�P9�gt
�>��<F�d��u�dz�/3�&���Du�x��%#��`�0e� @f���f\�z;��k�`�)���|S��?�������:f]���j���Q;����y�/�f0�W`�^�ɚ�"z·Qx��k��yr�[�J�����S}Q�oX��s������WQ�.�@�Vߟo�L���*��.G������Oګ�8
8������8L�e���p8ppJ����c˾3;:��X���8�8���ցU+yO��+�7�|�t�	�����~o�P4xn��W�)�v�퐀���x�_�����s���km�
�/d��-(c=��,��_eT^#~sh����n����I@f��5�x����|�!?��я>2|�����z`��Gt�я?�����瞻�������ofNiuԡBx&,�߂�I��dr��6�$V;�ȏ8ˉؚ�Î< ���{���=�8�7�r�t�v������o��n�n��;cVȡOy�e� ��������?���;���<s�>W�����vn?�꼃��3����������w-^�F���Kn�S/ڴ�4������n�61R{{��#2g�����b��
}ge��<�0���`�'�ܩ��^�D��rٶÄ�f�eI�-C<���q���=lݮ]W{A��s��ڼ�\��|���Q�e�B���p��7�ҝ����w��]Vt�k�;r��p`��vgew*"J�3�vn}�s�N+�;��+%Pi1�T	�=A<|�;�jr�4�Ai��
k�.ǩ�εL��L��X��u��U�G���/׭�Ӎ��}��I�NbJCǫϪ��%r\�h�h �a,)�B����=����������Z'�BuL���e]�C���RtÁލ+��6|7C��}�Q�G��J/�,O{c�O��;��:��sXx8c�6���'V5�d��f�2�fU�`���l�������)�b$��o?���1�_c�O��V�{�1;��_w��KY	l
6g���[o��O��?��Ö7F��D^�	rlQ����0�6�,2�e�UL�]�AGY��I�^ޱ�w��^�7j��x��I�y�y�"U���.���C◧���9F&	�	Ƭ�Wu��T���F3���~���޵���~���?�������o�ѓ��9� z��+��g��><�[-�^�u�g��}��ᥗ_F��A"���Mvv$�7G���B6�/�+��ci�QO�̶1�⅝�� Z�~i���\�K?d��ۇ�����l��i��sV2`���m[���wH�Wz����������'�h��X�z��r��c��|�;�:h�{�]�\7��E�c4m�����3�揺r9�� ��O��@0o��@ǲ�oӟl��m�뀟�|��©`Q��#h?0��5=�|U��K_ݠ	(ެ�5��ͧ��%�_�	���[D\^��A?x���U��o����#I�#�Zk�	$��P��]]�lg�^#��k���,{f���Ə�p�h6�Y�Q���6kE��XZAk�R!��Z��{<������M�D5�]~_#N����\t�R����i\�%~X�>�{��f�����L�����է�Z�~�i��� �Ô�*êVNP7��U�TbS�Io�9��s����2ɯ,F��/��fvW�bf��xe�����rр�+�JD-Q ��nB��&��uH�佋�AK���7O2A�W�{������ALGT^:��񍀡8�7�jq�1 |O�����.t�k9s�T��!>���Buڙ��!ZD��Z�@F6��0G�>��t� c`ty�|��o�+!�z���I x8
kݨ~lN�^��?P��`P�]��x�����;P^c���хҔ������r��a�F��=�0�3�a5�x��"�	�+���2���g��,�g_�u G�V��/g�x���p�m�ڶ�۽��Y0f�(�l���(���lq��s�{�� w+�Rf��'���a��X�A��^��=��Y�(���@ǑK��lEg�2/�3x��Ǣ��B�O:"ޘ�&]���͟W�,^�N�mU�;f�<�2����:H �Y��<4��7��@�a�[���Ӱm"�Sv#�)��@��9�G��в�e�V�%�~�ZP�>���ѥ?c;�K/�X��QZ���N�8^�������<aB��Q¨<%O� ��u�0k<ȉxjzv	���H���(M(��ݥ�!������r
�2�|X,���7�N3ی2L��F��#�w��Y��?#�B_����&@{!]�Y��j!��C��e��y�tb5����@�p@7�<)�޸\�����?eP��nd[1�:�|�]d�Ã:��P�O2]�zǖ%�&"�����`�I	�=�����)��x�[�xG��yC�e�_����]�bE�����#Rly��rq��g�E#�.GrE ��({dw��j�DOց���2�I�jnۤ���d��_��K9����2��3�G�����ݻv���V�g�� �ƌ�;�D��`��	5J���wF�F���>|�%v:.�d�nw�Q�~T��V��t�2_����h��54��Vv5p��+�������1i�d	DM��އ/��.�! ��8'z��2		�M޶.���D���p�������4����&�[�t0�o ���	 �]��I�\�`!����j0�����]:1[�M�/T]�h���:����~H�XZ�d���#E���!���H��Xfey,:��
��¥�	�ʿ��=a���F�Y�K/�22^�PX�7V��X	A�GC��� �p��%���^�x�
���q�ϭ��RtY>F�&���!v��}�Zqg�(�g�'�Qt�1gPQ�����3��B9=���ɝ��o�q#k<����H wl�PhX���ar��[9�� E
ݏ�%.+��/�Vh�?�ܗU�q��7�'�I�W�a&�N��t��_�F�Ga����^9��u�6)�o���}�����R�6H���l�2��>d/������o�O��g��%xl���T�t:T��z�O�t��V@Pd�~x#{*�o叕=�r3��� �$�罕��S<HeƐ�̘D�f9{.Y�`������E��M�� 	~n޼�|���HA�e��A�}���x_㵲s�O�P"�a�=�՟i�B(Q���!�g]�!xa[Ưv�9^Ux0�?�m������l�����AV`��qVw��]��Y�t$^� �$$,������W�ٽ�r����:��B��|GA���s&�
_Y��약�/a���19���c�f۔G��Ydfk�.ŵ����&^!���������X1���"��J��]d�7��.m�����v�80����D~����&�� "p���L)���b���I�]	��K�ݽ�lk�]J�D���4&��DO�Ͷ�v�����ǁZԷ�'���������0f�:���B�UR(�?�<����\Ì���z�˙�4�q�me�Ν����3"�t@��ˎT ӑ����y�P'ڢP��k��k�;�c /�=�a�K ��PWF��ԇ� ��8"s$ɻ��,4��U��y6Vz��|�����!y���tZ$�8W����F�fA+������r�뚛�`��_�z��7�Q����V(�Ǜ�%���_���e��S�����<�F��#J4ޠ�:	{7�������~!�)g|��mED�
�~M����J��*ց}������r��������Vf���zPoR��tBt(M Z䤷M�Ǡ���$�:JҦ����A���2��R�8�a��e��YB� Ow�tFL�� j���/QtP�c�G�؎Bޠ��t��b�|af��J�a&*��.�pX(��g�������_�Ƴ�Q-'�~�qV�n�&��RQ]:�x��w�b���Ivt���(�Tg̵l�:R^}���ҋ/y6�O�o۶�J3�|'�r����o�|��`ٻo��ˌ&�!���$-�-�F���>f�/3�����I�i��Y5�������7�Ɗ������y;��4w�hH;4�;3l��<�>��g��=�=iǮ]�k����M����9��U��blݺ�|��e��뇏TH���>d9���ץ���Q���]jB�56��kt4rs�:E���^�0 ��x�4bG�ږ�ځ&~l���ۆI�B+����S�~HHO~o?v��[����rf�e|&RR)k�ដ�?�Ƿr�Ψ;ɛ�cǧ̚�&=���
y���cG$sb�JZ����(�Q�b[�?��:���W�S�ٖI���o߾�wWs����������c���E�[�4�b�A�������FH��=�Lr;R~���O�3L�gf���>�.��<T���b�F*��hd���&�� 	X�G��w��&b����V'�q��) L�E���,�y@����l�.D|T".����;�KJ�}��G+?�h��λ�׏�9��K��3fZ�_��Ơ�gOK���lK
�>/ċ�S�����F�j��X��~�1�V��w��a�ϻ>��C��i��H7`� �(� �k�M�ѿ�'��� �36�[ٕp�6��J�ݿ�`y��7|3���<c�X|֖�4��Xq"��X�"��3e���~�Kpm3�̖��R��\�dq̦����p��i��.��	V��C�+�j�3�ϔ�^^������>'�,��׋/�d���]>^��3C��y
l���
]�1��g/�RBi�̲����G]�=2�A9[a׫H':���ѣG�{f�b�2>a�_�|�R�K����m�^��_k;¾�Td{ �<P���Lۏ�Asv�qx����Z�� �EgfQ��!�(�i�� �z��sϙ>⥬�%���±��?r�dyƉ�&��m:j�9z��M| %o3��WZ(������N��^�e&卢�ʮ��ԛyȜ�[m��W�Y�W�_�� wxaeWu�~�?�D��/�a�};~�����w��x�Ё�����<��������F�E	��'=�۴ic��u��1�Qb���;�_� b׎���ͤ�(���&��=�^��x�?�1���A���{h��w�/`��ټ�Xu���|�m���8�D�"k�W&�+�,��F���+:�y�K���Na�a�:�l����)<�&=hq<�x�咷�(}L´?��H;�~��xVL��C]�����g�cYS�� ol��nӦ�+�O�\�P�C��d��+�u���Eݢ�1A�dP��#�xuB�Mmh �L�gjൄ6�������
߿Nc8?�s��ON��;�:6j/(�W^_�����J���{ƘP]�;�}u(��ef��wI�dpE���pe���	p{|�����GX�0�#(W�ADP2Bf��%���(�.�<ga�e� ���/�0�A�^H ]KnЕ8�װ�����߽k���U|�
x���ˁ<�@�;B:�gVJT�=���E���o{�j�Z��ۢ�3�
߱�҈��R�p� �c�Leò!3���!;�3{3�,Z�%F+|��N"\�b<��C��:�X+�����'~���8�-���L�Cb���"��a�;]X?�+�����1
���\l�6���=�t�t��IQS
e.{��.1��~�I�f�����+/�M7���T{�����)��Aƪ��Pք5_ ��n�w������C<�-ɗ��:�xN��פ�<f���m��{�纊�4��X�J3��i����Z!��~I�!��L�0�E�{s"���V�́�	Cg�D۝ ��0}�aԿ0�U�qБs@���Q�`����Qn(��J�r�hFŕ��.L�ڲ��.�ܦ���@�z@�QG���_vl�idU�zK<���my���"�MH�7V�X=��d��Bhk!�E�$ćI`���Y��o~�=��ܤ��%{� �Q1� 3I6 m��o��	9��'������J�=�@b�ج�|�
oUx���|�.�S��㏷���|�l�����j���i���y���M��3�r�
|�б=Z��SZ����D�-��K��\�t:�͓+��F��9�YǼ���J�g�j�b���6��^8�/%��i�P�r�=�5ڱc��G�\yꩯ����_�j��H Y���,j�a�g�@�����mE|\c��u���`���0�h0���)
#�f(Q��p+3�̪Z��Pp*w; >���	�m������LO3BNO��1��Z�#g�0��5�=j�X��O�Q�Ι篋�@��:H���֯��<��iI��|5�ы��|@�D'��	�vØ�?̂�� ��,���\&\�,�S�C/|���d2����V+�|�w��E��^d�9�t���YZxE��n��g^����	Ѥ?fys��DG(�m�`kx#��{���o*�(�1�~�3����TXg�=#>��]ᏺǹ�w�mc��3l�́����qǎ��_,/���:{\����t�F[o��j���8p;s�P��v<$_�n%&`5Ⱥ,p\�}MN�Hh�I̺�U�f;B�`�riV�� �\&M�Xغ}�Z��t�-9#��-��u����@qވSV�ȇbU�&.�2�c�� )n�!��3���j{�6���{����C�Ц�r�t�LPwC��~��mx���_�%�]"� ѨZ��ڌ��;_�'�8�?B�B�6h�N��#:}�͛/!�tEY�����#�����5+��Ԯ�r%b�߬�lW��e*�v
j� �!M�D�]	�M�s���
��at[�,�c��[�o�g�0*�8�#3�O�L��4�:)�7�x�B̾�,��f^Z��X���E�,�Hp#�� �|�6�^L��(�����6��zV�)�R��I1��-\�`��(X�U����A.���r�!<���c(2Ǎ���Wޑ�t|�{�#; L>:Nd�Q��x������%��c靎���we��|��ha�	q1`g���%|Zw��.��;v�;wxv�Yn���p	��9A�z�5f/�Z��N^Hq�M&|F����[:���7��O�ܮ�;���{���HI�j��V|}�y)����<��8��2Cu*n%��d��W����w���-w��@�OK��:�����*�w��V ���ϐr��� vόW%7���~��Oa#] ���0U^�P"�G����[�[�����2��/����_�W_{�J/u���#J1[��/��cP3�C� �ߞ���'��N�7�F���`�bV{���o?�qG��'g0� �_:�ˣi0/��u������~�ܿ�zI��&�#�dҬ�qր"E��Ĉ�;kFY�$V�� aR�/�2����<ԧJ��'$.� [��q�a"7&Y������9���� %mb����	�1�u��4b�3�% ����y��HX$H�Vt�p�������=Q���i�3�
L�Qn�bT���P�9mڌ2_��[o+���}rw��
Peo�AO��8��М�g�jd�*
M�(� 5A��A��x�����X�G��X��=��ɺh>�&xD�C�A`����`��*��Z�p�Ǵ[�


J��m}�,f�h��I�bVe
e⩧�*��v[�+w>k��L��	m�o�u�|��_5[��'&����Q8�}�r�����̒�I2��W^)~�Y��A'���JG����=e2�۟$O��`v����)�ʗ�1�/B�����1�S�Gz+����M���ò��A?4�G凛
�Y�D�=(��AF��z52N�3#�Hq|�/�&d_���9Y�|"�.P��+:�����������ϑO���H�d�&��ə�Θɬ�L���2�}�̟Ƕ�E��O��W��t�*��!��g^�T���c��v}t���2�i�'��ͻ(��ŋ8��2��6g�]�ԞP@���#�P	#�i���:�Q+��(`(�l[آ��oR� �3�(�B���W&��Ӯ1]�>�ڤ�b@z�B%"��M�
?���g�';3��>G�0�!�O����S�a3 �BӘ�2���׽��/v�Y�=�T�F�c0L��쪕�"|�B����"�
�&\TR.K�6{�y�?ڝotP8�A{���^�3��Bߢ^q���a��}�`��9�zD��>��4��~ժ2��]��t^�IH��%:�c6�Auo^c���$��C�E��p[�{�����#��0	��]��D��
F&�a{��l*y�-t.�����$#>�-�)*�#� �[����`����h���u���f��޲p�����np�s�4���AG%�k�f̘��H���)崗�cv��*(�#6�����%L?�p�z������D���c�	d�L@���Qݫ�U��6���o]:|*��UG��,��d$�Etn(�(��g�l�K`�����)��wG�L�pE��>��b�2)T���K|��,U @뿂� %��5\~6�zE�q"3,8W�!P#N"����;�_z�J��?��쎸a����!�����#w����
�x/������2�L�����9�#X&����;ZJ�Xٕ_ ���Rf�Y3-��-[��)#�4b;�߬1E�wV����e���VW���|�_*k�jp�r
��W���2K�`��,}��J�ѐ�eA~����2(�čt����We���V{�YVE�eV�3�z�	�2|�ӏ�2[�����`�;����(��g���Κ2�l�T9�d�8���n�S�E�:�]M��mW>@�)�y��9ު��#?1hb`ɬm�r�1kK=f���G8�QHb���^0HE����9S��=8�~�M+s-H�8�5���՟�WN#/��Ac��8����<G:�P���HK0��L�  0��N�� �2��j�A+��N��f�C�f=�_J�顏�}�:a/e�v&%�"`�1*en�x������F[�β#�+l�b�Tl]B��Eg���������L���2Iµ��<�p�Q}�\ţ�'���n�.�)���Z������?W����]���+v�#F�/���"Z*�a%
3���	e�8A�v�=��a����g�uGN#MAsNB	��م�xI�Ob��5�B�02�\�`q���5���(NC��=k�:����!�+U\��ቅ�G�C�O�y��(��۫���~��A�~���_��D[��w���QdQh7\dΠ�Rt�ܶ� �0���5 ��^f����~�B�C���Ｋ,]�R4��Z������=JE=�B�M"7b����ĵU�=�(̤�h1	��(�L�V0�,1��R;[
�9�zok����bf1��|���2��P���"�W�a�_�����e˖�,�c�jP�B��>��/��Ϻv�������@*j`�Z�)O��b�z�꠫@�ɀ���v�(v��.C�z>q}�
0iS^�߼y����rx/�"̔?n����^z��?fG�p�Z�X .�5�*$m ^"���b�xm�kb������(�N����J6ܷW��>�4A벓A�H�S�s+��^��9�f�� r������w؆i��c��ZC�޸�WLh��'�[��qۏ�KuF?�����ߏ��Z`�r+������}����fU]�p����Ζu��ߣ��L�h&�Q�sD~/��!�`
� �*��D�A���P9e$��$��.A�5�%��ݷ�;�w�}��%O�{�)<p��=���{˽��#w�n��a�Nn`����`� ���r.7^���Y��D4m�0�X��8��c9�YcyT�Fl��[��}^$���SNxfwϪC?u���������J�BI�0��/��<$R���~y�_�Y�o��=u�:nvף" 1��A���f~ا�}�6+,��_����_�^���~ϒ��3�a�
m��H���wHI���+ݮ��\v=˜�ǎ�<P�CT�(�1�3�(ў�Iev�Y�sVZ��m6E0�I�ˍ ���%I��)̓���g<>��w9���r�ȤD��,E�QN����f���|do(ޱ��9D�<&o1K[g������d�5����en�`F&�i�Fd�D!щ*at��濗��#p����d�Q�fT94{�#}x_(#��0���~�Íp�?����
.3�/��b٣|3k�(�1�5y�~����1��@����	�EbB�y�O��h�A�߃��a�p�O��9�������f������n����@��?�=�ʻ��ХO}�@�A� ʹ��F�����GC�$�Ӱ�3dp"�Vh��(�,�M��"�O�����!��?�cP�!5�.΁�)������A�&?��n��gC�TD�NܩN{�~�V��"��K�d��v�B ��ỷс����/�F�+*�"��IL}�]�A��CH�H����m�����|��'˗������կ��~�ǯ}�����f�ַ�U���o����o�o�w˓O=U�����%�SչpR�>)ȟ���_�&�5���D�3-��	�����4����eٛnZ�8�J���Kc(�<��T<F1(\��a��Y��A��#v8?]�׈`y9���B��]���S�.�O��yv��Hk��4~TOY�#Dp��1h�-[<[��?��[6�p�/+n(9*���z�`�����[��c(z&�?ZZ���h��~I��i1�����D�A�BK��³څ� ��`r�/O_�R�g�gC�溷(UE-��ٳQfY/���y�93>��¥��*�"C���]�����{��lle O���a����� {[W�X)��׻�$��J1<y"N^3�a�6eŇ��KJ�{�M��*�[�w��h?���8g���eNՙ���ۚ����\w�N:~�y�7����R_׭[W�y�m�F����@��2Up��b���ԧꆞ<\v.3�S$�Vt��6�F�� yv��؋͇a^{�U�w�M�'�6�SǬ̦�v!��,�*�� �"�ɥ9���j���v�=�j�Wk'�P�G��˳����Fۯ$_Z�,��oK8\t1��G���'�l��ҫ���^̈́6��y��rP�����(Y���7l1b%��)�M�̆�b"eE�
���#�v��t�IfgO��a��<�G%���4J�S�s�p�p�KoG��L�F#N������,���G�����Rp��S�|�o�?����
w�&>�����G���(Ǐ?��7��":�w��h�$�'L����������~��u��f2���u*�g������B#7�pc��U+o��8LS��7:��A�ݻw���P6��𙳧ʜ�������Dؠ��Mq ���/�x��XMa_̂��ɡ� �C����c��
����Q<��q�4�.�ϿZ�.S_��4ͧpY���,�྽{�k����[���������R�=ʒ��+�d\b�?�~B�EğU�(�����T��ľKh!�u��K�9��P���v���
X�ٌYQ�]Re� ��|t�1��A�ؗ���4x�fx�/���8G����|&���ǀ�K�u��q*]��y�g9��������Vr�_���I����C� ��C$�c�=��Jn�B�<d���	S�N�����s��w�}��[�}���z?�t1�9x �X6^|���u��~�L�a����:)0�����[����[�8�\?������L��={�u4�<~�U��H��L���q�ƌ�\�5�:g�w�o����Nxo��v���˭����l2��03�9���*7L�O���$��.�N9O���V_��J���Å��R_QrSѥ�'��)��_J?{�}�[|bKWFѧ��W�H����4�	����|@e�iT>A�|�K��{�1��x�.1 �`�f�)f�+��Fn0��8m�;[��~s2}�i�ث)rC�H��
K:w�^رF&�.�;W)Rɥ,�3���?�[F��%�,�s����a���K�\RX٢��ć?�T�5>D3W:N�%ȋ/0r�*m��
��/�ͱ��=�V�/�V�/B#Y�W�C֓Qe �P��yfk�G%4����Ȥ��"�6�H�(g6=+?z�`�����N�+�n�y���\�J�2O�=��si�\��y��&:g6G3�Gر�
rO��Uח܆0mF�?k�+{�ؓ�M����I��B�w�QUe�����i���oY��,��D����4u�������٥B۬��f	��R`H�('N2�u��P���Pi��Y-*2B�FAg�	�/�W
AS_��`���>�@)QO���]�f(jsf�=N�Dл��Z���B *�W=X���{G�c�h)��j|f�@f�f1ڧ}9��!�c³g\�t�w�x��|�2���65 ��x�����i ߷��j:u5�k���9�6ϑ��縊�=�yf�YySq�0��� HyϬ�Y|�u��?�:��_�$�f�y�P|�Z�%�y���ț�uG�A����,�c M���y���BP���iř���Hv�O [(�e&��|=����g&p_�rU��`��622��9��n�g�Y��W���7������k�>/C�ľ���>^3F������N�r�ù(�z�}�g�[��Q_���S�1c-���@�2#f⢃�t3�J���\.xR���
�����QP�+y�ʁ���_�� �W���	�E�d�<�p�����[�=�	�nܬ���v��\ͦ��]Rz��w��+e	�p���Y�g�͇P��9��kd }f��]��2���"\�Ȑ�_�q�6ω�(�$�0=t�*��=�u���5�.͊	n0��x
aG��/L���/~@ȳ6�x���?�^
"�D��	L�����B;r%)�s���I�k�BM�Ȥ8'���<yQ�R�nETj�		�竄�}-���ܯ�Z��MDIL ;�У��&DQ��$Ü��-�%����#�BU�=V8£�-�"�t�3���33S4�H���c?HtH��N�%C
��Q��	D���p]�|�OB��qx�q>rH
��n���KpU>N��b`�Uk��Ğ��ӣ<)�?PoDC�����>H��� d���5 �;J{�<���� �vmOl�{�-�BT{U�E9ۼeK�@�_����6�NE���h��z��m7���Z­��r�N�=�s-�� ������ُ~��-��h�=�H�)�P<QJp3�PX̗H;�F�R�$���X�t�p���q74�i*��4����$�90�����r��^a
��`���c����";x�p��9�
/eй�wV�؊�_m�/�xo��+�L̜3��c��ù�O	�s�ݞ�N��&n�����W3��*y��E�;��� Z���,E�'�@gy��!oE��w���މY.W��_���u���'��Q�`���CY`ࣔLib�2��(��;�﫺ae��b��钾�A��d��\1@��l�?VY���#.���&Q���Svm�Y;xD�� Ei OTG�����x����}��_���{��ND���f�	n-�_�ܧPm���K�a�F>Z� m��������0f:W

��������3���À�D�2Y�V��:�7Е���Z����l��Ў�3�QnAcyKIr�����@��p�u6ܙ���PC��Sf#� 3��/.*�EcMa�!lU��Y5R/)*�t�:d�M�����n�b�"���Ũx�<�$�<�:�8�P�L�m
-
�����Fʭ�%,�[X�ME�+`(��3�Iㄵ� ����T7��_-l���
ԛ_���sO�Ξu��Z5�r�����R�T��c4�e�\B�4��?qLm��̌��Ō��1�$���oo	��aeW�����'��c�?�޵��)z�4r :jܑU!�'�4a��<G�2$ �Wn�`/32��}�x�*o�"�cG�I��#g�4o�`�@6-�h[��t��)�I!�Y�1�<�8{u"�鞐���f)�l(+˥�G:��3ki�Pș�g�{����eϞ�e����b��%��
�>�i�f��Œ�KE���;pTQ��KC�w��� }��ys˒�Kˢ%��d<��#�B7n�P����3,�;?�E�B-���0GV���?��b�i9�3(aT�,�TH:��

���'���m�v/Y�����6/�6�\i`��9�<"�Y�FX�/��$\9\�� H���<���?��{���iA�h��`�8�6T�#��;]��P6�g��l�����O#�46��`�#����&�i wtA������3a�ð�ہ�q��D1{��N�*��03A��n����q"$�Ä�1�LtF�)B<Gc��$H�h@���D��-h�3'�60���ły��j�|�}�3�P�2�Fטd�4�޸�e��O�� Y@/H*�t��YM:z��t��^q߾���Q3�`��K�.�*NLu��hM��Ì!d2P����]�~�|7��~���	h�B[(�WA�'һ�x�0\w݀2D<E��B�����`w���mZ��u�&�,�[�Qٲe��`�S@qD����,��Qf��LY�GY���E:[fЈ��G���+Wy/<+.�,�|���<r��{��ܙaE9�g��<�N߃�I ҧM0��Y�9{Q�r�e�;��,Yd��M
E��Ǐ����?��պ�g�w��	�Sn�7dJ
�b�-���w)�LY�����'�g��q[�q�Gyf��� ,��U_\�u]Y��zoC�=y<�������!� `V4��,�al�?9���,>�	�B�s�g�٦A}C��g�Y-�{��o>n���& ��AK�7�ԇ�� ���r�	�OT6`��	�C�	��Ɛ��k0��-M��]��:�V>�ѩ'�1����"A�D{T}`፫W���(
� 4�G\���Rف�n`li;N�r��Fb1O){���x�)�su�U@χ��0���X�����v������ad�3�xb4��D��q�vFވ/���3��{�'2���I��`��Wd2YEf|�rXM��c�݉��#�53�[�p��)��T�)E�EHmٺ�|��G����o�Q^~����oz3<#�-�p�)>��c��7��30س��9F���Y)θ1���׸
��X@$ (���'8�0����TH.R栉g���{&aˍ(��K�+K�!P���9�4E�\d��Z' ��oR��X������X���aV}�Ae�VgF��>B���'���+uB�Nq ������Gʽ�ܪ���L)wF�^� ��Uޣ�/��-��t�!1�Le. �M���ɥ����
Aͦ�a�N��C2�XL�!��N�>է��-_R�/_\f)�Ї���5?�,r��Ck����gw�m~1��ln�#���|��w��f�P�PV�	�3��<�������D��U��X�)Bmř��Vj���sz(֒�l &8����k�Ω��E����Ԡ������:H����u�C'��s�n�z9��g���~���
�oW���`�rc�;�[��C��!�n�Ŗ�+f�c�ۀP$��X�<�Zb�4L���	��n���=|d;����?�3��Mf>i��f���˭kn�ū��m�q�QV�����I$�ڿ���pǑ�V���~���y9��0Rv|��%���óg[��Dzz�pȚ>{>�w��6�1��6Z������KA�.c�m�Bs<9~�#_(�a�Y���C�:H��Wdu�kWW ԻQ��@bD�Z6��*l�u�	33�&఍_�C�2j�T�ܼ���?�A������?��(��O����_�Uyᅗ�#�C|��˫��R�y��̳����C44���\����_1� )u �cH?!i��oܩБ�\�D�e*!�	鱜�L�;ufs%8Vvɻ�`��5���9�B �'�������;cY�z��^	7����=d8�T�ӆL�Z�¯*��D���j^T�mQ��%[��_�@-���,p7,u��J�����d[�gpg�� �W��=��V�+OGJ��-Bm#Ow ����'���Y�y���}���@��B�h�~��Eag5Gʼ�(�G�M-�R!��kls:)�Ġهʪ�
=e��W��&�])�U9����z�P�pc�e%e��_�۟q^'B��|!��'�;��xC�f���'���ڲ����e�W�y�{���6*�n��z5 ��#W��g���3V1��c��e�1��M?ܘo�7��%���-�{�r�:�K��Sm-�S�#ʠإ<��o��Fx�*�2<q����h�l\�3f��Mt\o��y҂�e�K[����0M��1��4�m���A4f�|CI�_�a͏��ߣ�$]O:��k���<�F�xn�j ���c�#�l���#��}��b��'Eyȴ��?�����+���M��Q�S�m�����F6Y�wF4~Ok0�/c����� �৭c�]�Q
N8p9����6��σi(���ʘLN����[�_>W���3���^/o��Ny��W�w����o��+����/˿���������۫���i�)����W*�e�~`����,ԑ�D ̈3��9��ĸ�Ǘ$=�埮I�/�a��>a�|��lɲ�t�Ru�Qn]S��w��$�hl��M>�h�7����C�=*EC���!�FW���gh�k��Pm�e�����reE��I�{�F�{�=�{�V۟Q֬Y]���ϗ����-�<�pY}��^.憒��3��MQ<(�t��0N�V|���A��2�V�wTף^
F��q���!��_:��(#��M���!��#�3m��t��n���z�� ��A��󑃳p){��/G�yB�J��E=P��ȴo.��ي�'ڡ�/��D�^`�,Y��,[���f9lC@��V��e>($e�{ŗ,[X��X\f�,���2E�Ld*�,[P��s�G|w��ӡC��))����������@7j��'O�Œo�(�����r"����+��3(ؠ'�IٿN
�x����?�ak���G���^��Jol3�k͇MP��`�ʅ��Ǡ�їX�U��u�z�^���>NuT:��0�9dZe
nwQ�a51&Jf��W�Z��b����5��ڜ²�8{�x��;W����ˍ�_��i����J�y��i�wE�������w��?�����߻�Qݠ{ۑ�r���j~��/�@����I�:H_Ox�<�^�P���q�Ӹ�L�E6\W��F�1�N&��� �=��l�lS��T�Y�e:�p��,S�a��b��|��SB��;������J�I�����D>X��o��X�7��e��]��L߼��X�s!��_#��LW��W��d%�m|+ ���tTJ�$�?�䳉�p� �e�`(���_4f���qq='��'���(�-6l,~�Qy���ln�۾={��g#��AzvB�3�'ѧKx�qC}P���	��Oq�Q��餏��eD���(.�0R�[���8=L��N�"f����� ��T
�*v��м����C4�кu�u`(�A������M���6�|�=�Z-c;�6t�u<�Ѹr��K +��1�j��媾[�E}����y�J
&K���}����`�|��A�G�q��T@C/��]�x�Π����ٳ�:��ﱓşÔrpF��ٳ@��J���%=ߪ ���dEM� ϑ�4��!�-�.g3<��l�}��o:�)�(�(��d߻z���?���O:s�2� _;p�g=��@~q�y��@��#� �8J�e�@��&��Ń�t4��	W�U�z�Iޠ���K�� _�c/�RQ|�ˋ���*\�|6����e?�`��+�}d-��Q�p������b�݁�?��㢮�s��4f+\���r�I��P
h�p�����#(�x3H�����ȣ��]�R= O�e�p�5��xQ�]�����(�MEe�xΫg����/�dHi� ���<.�K���#����BZ��N��m��5�GY5�\��>���B��~�)#�G�7�w��}؇��q��秷c���?��D��Ɇ?oR��R�80��iF��T�0� ���TLZ�Ȫ�3�<8F�]L���HQF��xt�Xf_@Aj@<�Df�LTp��{�;��R�a�#l�Ɉ�_��xS�{�F�Cn��Aj0&~H7�����n����w����~��0܉�E���N���)Qdf;L`���S�,"!�'F�B`�Y�
&�\��k-���+�Q|sE��6�!E]=w��oE{go-� _�,�����s�4u����{�>G�<S��:����_���ʞ��wBG�>�9�z��[۰g�x��i�s�,P�p~�/�B��"�;v���1�r�?d��.���N�p���%� d�B���WD�L<y�-Rr�FKaٯ�L%����[cY���}�ęr�$����&މ��r_/t���RpS�C>�U���t��8�˅��1x��=��ɏ�1�j9ĿktM�,��A?�A��P����� �3��,+׫��s��?��C�Ue�/�1p�x�+u�`-�)����{�K���A���1������r�w<����|����:��s��-PNj��F����~��#Pt p{� �|�Y_�y[������0��� �]ۚ���%E�3ᢑ6�$J.H�����994"c���k�2�H��q�Q�Ȁ,ؽy�OЦG׋Z��M�ԙc�����ҝ4t|μ�3���	��l��0�ʰ@���8���a�+�'Uv����)	�����@[x�	���a6�!����n�XB����ЗkT�Ѱ::fV 6;]wf�޸CI��,�4��]"�fQ�>��e�h��Ϭ��o>�)�@E�1�v��Y��n�C�B���g�_�캲 |-�kc���7����9P��n�����
u��i�(�1��h1��R_��-�
$���U P��=�A�큮ae��[�\���//H���Px�t=�)E��)��33���9�c�N��B��k���'t�yp~��!o`���ò9��g����ɞXu��	����S>@��E^I�Ŕ�����Kz�8y��J�8c��h1���y�P6Pd�k��-���[o�T�o��xx�ha�5�#|`/����\��9.ä=�7��?�L|�x�@1��>����qC7�X)p������ǋ���J!�>�aK�_l���p��1nA�OP�Pz*{�C�F�����Z��SG���"}�D��ٕ�P�3Nf�)+?RP�7lX��:?���⏸)�y&�7)�wH����˗��Ry��}�2_D}��7�|`�҆�Λ�����g��ES8���A7�2ū"���{��S��N� ��'H�`L�N�_ץѵ��kat#��<�����Ѕ�B��p@Kk��Tb�,�J�I�=F����l�6��Z)�W�/3��5�@~ڌ�J���0m"\}����D����Kb��5,c4`j��/��#����i� �F0��߿��A���������^���)�o~�eɒ��o�LLTl�#fd�����i��P]�$ ���ΛSV�Z������j�]��r8�Ywt2c@GAe�^b�튫������j�I�O;#|�0wk�K0���R�<��Jhi�߀@E����V�h��V���λ�ڵ���0�=� d��2�c I��:�Z�Q�	�c/(-�%B���+���V�I뜕�e��@1b�7ol�D�w�V�PH :#��cf�-�t�J�,�y'?��Y�r%�Kh��?tv
��s��PtS�؊�B�3��V����@�޳{w���˻��c�=_J.� ~��]�6d�
���a��&/3��?�� V��Ӫ|J*{2��=�|���?�A���V�y�������_y�<��s���Yy��7˦M��Mʖ��ˮ�;5�8���G����G:�9����&e+�~p"�GZ)NT��N~�����EԳ��w��&�]M�3��;�3�RF�g� ��~����믕_|����?,?��OU������� e����(�g�r�S��K-w��n[���
��e����ۯ�����]ć��k������� q7���+��3�-�v*���_ɫ��{���X�%��[��D1	:KM��6Þ�	�:�l"�ߠ+}G����c`(�����Op�"��k:�� � �5L����#Ʊ�.@��}c4 �Pa�(+�m��Lđ��.F!A������.q%#�$\oQG����;��+�O�+�+O�<����K_��/���A)���-�8Ux���*�8F$j���޼�&_�͉i�
m���Ά��%>�|-\��3"�i���H�7B����.f@R'Qa��a�����R�@RM2�7OXy��AT�ALp^&�_'�RzͶʳ�B?'��������u r�� �!�
�6��Q�mS|����.\�@�ʭRpQri��]+xy�ޢLC�W�w:
o
z���6�َH��V�L��@��A����x��y�#~����N��)z�C��aU�����c���[�	�7���Xz&NH��o9�PŌUr%~� ~ݎ�oH��c�L�Ѓ��1�,eX
�e�L������i��U`l]`�g����L��l���;ʺ��˺u��ƍ��;7�|�y�o\�F�,!
�!��yS�!;C�Sb}�:��.��H­������p�!y�O[��x��!���v�,/��b�����ˏ����k�H�{C
ݫ��-���Oe�|��})��Ν�����r��9)�R	d��>��df$�B
�S?ċ�'�A�DY�f�"���OE9��?��u�i:݈��b�Y�W��ٻ�l۾���G}T��}L�·|P>��}�Xޑ���F�>����Wg�Yɍ6�F�����k
km[`��?���B��v:�h&L+���_�/	��O��h6��� \C�	)ڱ� �{����us�bJr}N�P�04v�=��}2LH�SyV팶���귒��XY�tx��: ��*a���~���'�d$?�8����ۯ�4�JedY!o�����%2�M��̡����6X�gΣk�g��n���r�=w{on��gO��T���q�Mb:�Q�/�&�Z�.�j*e+�)��Ip#H��V��*��G��J��U+�m��S��}�3�l��§3���f{)�̰�Eg����W�͜��Ot���E-��Y ~�.��_��g��0x\�6؂�)��!���SXĻT�y6T�"�h��0��W�o��u��/�߆���}��J1�O��&�)*�ʛz�wʙqD��x\M��h�?: 
+(~˗/-�/�߰�maѢ��o׷��4'eQ�R#>:5��O��[Q���=�ApK�� ��ֺ��./1!�E�`;�9u��IǍ2������)rE�U$��2`�p�����נ�|ٸiSټy����ñߖO�d+�V�N�9�\A˵'����pd�Ås|�(7;*��(g��P��V� ԧO�L�K9�K��5Y�r���ӑ.�(�̕�d���l߹��ܽ��ݷ_J�����������2_�ҳe�v�]�G4�;�J/�9r�X����6�r�jbM#|�}�$�]�nb����>�ꌘ�K���m�{���W]$_|�:R��������eǎ�R�6���6�-[�K��\��R�����e��e���IƟ;{B	2�"y���9]�iSToΔ����ݹ�7��PB�xֺ��Y=�Vh�3fb7;�0�B+�y̴S���B�9��
7I:�����O�=�z'$n+�j��O���D�X
.��(����ZyK���y�����M=��胲}떲��r��a�3o�Ⱦ圶N{9GW]g�ג���{�wI�~����l�$�	��j��هQع�;!W˾��Հ�֊dEh0.���wL��w��l!�m��.�X`Ǡ�w��N�n���L�����8�ik��q�O��m���A��m]�qK{zƯ�_T}��~�~��?P��EX�s��!���4��o�F�]�� }��EK����e���G��F	�اGJ}��l=)��P�Qv3��7C�8�?�s"^>v � $�|	-:$����7q���*g<=�N�!v��ȳ��b�Nuj��h�	o�%���H쩃Fzc������̝���'g��KW ~�W��ot�!8ɳ��K����9�XY1O��Vtx#��x0]N���t���|E	���Y:����6��`�����J���o\ǹ_S��Dm�z��j��Ŭc�G�ͨ��?��\��~snZ@y�.{�Vm���r��N��p��U>�}�0ؽuA��`�HmPG���l�����+�j��� ��A1��Ђ�3�I@z�M���)�7yk��h� �'���V)
,����Ȑ�C��R�s�`�%J[
�=M���l�_����\P� :ފ>RG�".ޡ�2� /���4���-6{��3�)3�B9��`d3�,i3KM��)Nd��|1�=�(e��Ġ%B��$�E�E��!��b��A��D��{��D°��O/sw3��;�=c*�����~B�q(���kA+4����8 ��+���N��+���V$A��q8�1�ՠ�#]"tc*+�]��ρ}�(槥ܒVG�4���3�f"�W�q�pɒ2�F�?K�.����+˲e+��	���.]�0Km�7WP�5�~Z?O|��-�H*�����ʛPQ�`�7m�������\��_�$��wM�'���	����ف<F^�O`�ϕb9������αi��p�-$��j�]��ë�!��C��1�rX�&���>��~���U�x�a&��a�>���Z^�.�n�����y""E�g�����#LS�e%������1��+*|(pA��U:A<���]�i4t�-:�g0���!3����t����lEꣀNe괙���=$<��h�t`�q�B�� Бq8�����A1#Ng�?�����JcV���b�����X��J�,�MB�����t�C���7�=C�M�����t��ŉ����]�C/�J��R�WѦ��B��΃\y�
9��;r塠��B��)���pq9��S�� �u�a��:����i� �/�4*�ޓ>�@Q���ʪU7�����n
�}}�lx�W�$%Wq�_�
.�/Ec�x<0�#≶�%�g�M������$��3hE��V*�kyY��߻oo|���|M�Q�	C�}��[F�;p`��1�Y�r���y�@#k�g$��L�QX�i3p��tT<���ì�1��#�~�����O�'���/�'����/�G}���C��.< �˃�?����*���@����4ȹ��~���5kˍ7�\/�������Q�wm�H��E�[����c�o�� ��A�<���!�e˖� ����k�{�1o�{ꩧ���k_�Z��7�Y���o�����_�z��7�Y��[�]����o}�[�z��o`�V�7~�|��_/���R����]ZjC_���ƀ�Y6�A�pނ��}O��~e%�|�wc���KA�yK�(�tR3�dr+�������/�+i�ז�`i��qy���w�߆��v|�����e��6zA������>!8����={�[�8���@���'��I �<���f9s��>�9_���${�@�w���[o�FdY�a�M7�/}�K�!�;��MN:������M'�}םwJx���,��iS�{ľy������[��׃��I{��N��{P�<��Lt0�YLfE)ϜŬK�s$8�xDM��g��=��ig_I�t�T�s.��fbT�brBq�@���U�`�Õ���9�gp�v�d�a�÷0��8.�R�D���1Y�<�M`�pQGW�\����Q �������i>������E�b([ �ôy�^	{��Gܧ���Vio<�T(g�3#����͛7�C���e�f�Nဟѵb�k(��FsUV(-����&�)�]Q�ت�}�v+�����/��L��:��#��mR.��X)-�2F޸���+��|�b��e���1�e6��~�-#�O�H�g))�C.�� @y̘>�aO+�P��yf��>,�<��e*3�(�(������ ��a��r� ��Xq����z.Y����g��@��� �믽j9ǌo��^�U�U _<(_5L�5=�I�ӖHrm�mk�J9�bz�-Rp�(_~�+�+_�jy�ɧ����ԓ_)�>�X����m>��c��>����J~܊1J1e��̇zD���e��[�{�@���%�=���Ӣ��/ez�' @@��⢏���w��}�ܛ���(_��˷~뷬�>�ԗ�#L��/=i�駿Z���o�������/~���r������T�򗿢��}���>t۶�S���=��G=���7�؝Eח�ҵ�^�G�cF�����'�}�6t<�쪃z���L~�[@�6�>ѭK�w2�̖�ղS��N�Ơ7Y�|�'��6�n0M��MG@�O�*�,�3q�����S���RL���	r�xpG^���}e�-�%�D�E8�`�7iI�@�EK,+"��/t*q�{��oXW6n��4!�I j�tg��g��#?r� ȗ�o ����/|���78:���t�����N2}2�G$�1�R�r�d~���`p��ɡH�!�9��{1�UR3�˃H�Ǆ�Ý���;[fIY�Cg��f?#_��Z.��=�Fѽ��,e�D��ҟ�X� 
3cT���Eel�G.q2�F���8��P#��n4C�ِ\�2Q4��Lw���.���� ʃ>��3[�\m�"���[n��7�,_���t����QOK��YW1�-��Yb�Y���~���<�K����|����]�|������0�|��Qu�[]�����C�"dQ�# ������s4��6u��t�n;>	
1c��/]�v��B�Ey�d����v���N�A�eBb69���e�����w��$:(f����=�����3�R̶d23��?ˌ6�%�RkV�q}�z9&5"��t�����жo��� d���tc ����K����ٳ�{G�P)7�c�#�w�3�ڵWJ�Q�o��`A��`g.��'�R�Ѳw��خ���QX��%�$�j�C�| ۶�R�[�P��د����_*�?�l��/~^~�������G2�}�9�J�������_(/��by�z|�[,��i|�w�w6lR��)����	�ĕA֫ah��`�g�ע��,�>�Z!�^�.�6�}/ؽ� �Ͳ@V�����s�.�i���!������Px%��,�Ҽ�}��.�~��?�m۶ͳ����ި�
"�D�$�b�
����Ft���M�K����}e{ B���_҈�C�E��A"����W^|�E��r
@ .Z��<���e�ڵ���@aE��ر��+!@�"����5�U��X�Y�d����͙����[:�[o��J 3f,%�9�&��7\/a4��ٷw� (AϢ� �%��wN8^WДP8�.9Ĉ0��������>GB׀�2\��7�3>���c���ޭ���0*\�U��I���<�L$ ��˗-����.U:J���yn�q���O>�}}���Νm�4�O��m$�ϲ��a�3��N����Rd
��}�~�A��݃�O�5uB��C�"���ՌН�����~���r�I�0�'��=�3R~Qҥ��aԕ+Wy�/��hP��8s35|��B9%e�w((�fiQP�ĭ�T�z�u ��3f2C-����7H�Q��Bv�۶������c'�s���ʜYzl�`֝��7W����Z�t�97j����Sf����ˆ��#���*e��1%A��%O&t�Q���6����Ɓ<|m�� �MeㆍeӦ���Me~�Y�j��+f#�mݦ�n��}�\öEϛ���Xoٲ��v��e������	n� oô��uh�@��}}4D�e��B�_ʅ~���]���J����K�{�׫�7��䛛9>��#�6��G��\��n]Y'$�{�ss�:��:������#����3�� �A��7����<�q�1�a��ag�ֆ�!���qT��O��y�3��$VL��C}����άc��2�Đxc��k�Uπ׸��2�;T��v�3�Y&�U.*an�@b���:�+Z���E���'��M��-c%��j#�y0�_�l��'��Ӧh����lR�]�a��(|��.g<�< �y�s�%��|B_d�,��~���GU�;�]�� �������(�G��V�1�e$�J4X� 
�=^+�>!ew��^:>�R�4T��^���v��b�#KU�;BADaͥs�U�ҋ/�T���FwVB����B`���l��Sa��[o����Êo`"�5ˎ��0���cO��`_a�2�Ls��p�o���yC����c���1�y��2�:�8G�={��X��0��Q�U���/nl$"`&�0 ��R���"�۬���0*m\�&i��aL�F��@�&+|9��ɭ"(���={v�3�̾�u��s�>�YYd���(�樓E)q��p�9*��Ho��L�`�� ��wߖ�E��px��:!��a�9\�y����m(��.m�pGbA�;���1=}���]��0B7xD��=fQ08صL�`ي��DΜWq�d$��qH��tQi��#ҡS@n0�͵g�]۳�� g̚&���(�;����R:+�B�W��bƌ�3�<S�I99*���A&�
E�t��ٍ΋� ��k_��gu��|��U*f���E[Q�{���[oz�!:D�N�%o��Ѽ��rPM�IȬx�\�b�]��e��3�>~��}��<���hyGyf;���Z�ޫ(���J��e���dbD�����%Տ7l�x����C*��'��M�a�߅=��O��J��N�?�;Q�����g�^�{��c���J���-|�J2L�����?(��(��Y%�$(���(cQ�1 �N�FO?��x�>.��z�(!���7z�w�:J��>O!��&��4�1�#�Pv]�rOӊ��9-�tY=�7�ND%��O��g�8��;<_���rHGAOE��G:���ńu�(x�^���W	oР���J'�8��"��˲�M��Jv��m�UR�Vv�s݂��kМ|"}0V��<����Di��1������8P �	&TF�B 2~� `#C-�����Ǟ��		sh�����Ğ8T*�$z��P�w���F1�������_�s ~fDXZ�[�3�e}
z��Ce���Vt���#/�7¶˭�'���=~���޿��~U�*�� ����g��E��zr��UZzP�w[sU����h��Y@�e�ŏ���U��<(S�
u�qɂ_%P�[	�{��n���X����=�z����=�t�\o��β`ђr�Wu
ܲe���~N�K�;~��	��ڑ�D&-���3S�C���Q�w�����J���$&i���◿,����������;V����|�<��ު�n�b�
_S���u�>�6):B�o��Ff�4�QJ
!h&��r%P��@�E�Yw:�j��)�s��~0��������$�-��������?�9�ykC��W�# dR`֩0#]��_0޵��ֿz���a��uD^:�5\>{�f-�&����i���P^V�Qp�7$�%$7��%}
���J~�>�~+Z�I��+��@���-�od'�"�"����� ���Z�B ��aD�A��8Ȅc3q�Pf�M��0��9e~��N��8��S�K�EK{��&�v���gL�@�w���R�I�s�"���K���K���̝S�-�W��6׳�s��u!1��}��)��<%��O�=M��+��+:s��������>�>�@	%�۪��8��t�Tƪ�3�	�e8�z��t��u�+aK��W�8������Й������U���x��*8q7�0^!t��d��wҳ,ԶY�a�M�P����-J��,�ue7�x��9��,'3 ���!��y��4s���l�fl����j�Sgp��e��އ{��a)�����Tg�M5��nݺ�������Ey����6f���z���u�]>�Ȫ֫��Z��y/g�BŕSl[a�B\,�3��N:%ӫ�◙�=�w�#��v$V�{��.�^>�@�~{u� �Hy��HK(��.�T��AT���<'�sm����[ĝ�;��r�>'�[��C�'��a�;�Ob��;{`˯�Vj[w�>\��ҽҾ���j=����8W��'�L��6b7�n��	��k��Oo�&�	Y�L0��u�����]
c�F�C����#\*@���,��Zȶ-V��/� ����x�r�O�i&�(�^钂�+���C`�w�'��f��]�\	��(�l&z���\%��X����"�c҉0E~��[�w�i\{�m����+w�y�P��oz_����SE �.x1�#fV�{2�'��Ukf^�k83g�<u�R�� �Rz��Ι;�'��/_�.��J&� yN�X+D�6���{�h/��	(/i��k]n�)f��v?���GfOR�M<'!D���a`����L!�J�$�a�\��E���+W����P��^ϣ!*�_jW���f9[�o��h��\���Hzh�����Ҁ����مr��1�@ǧs�)�]��%�B��_��W���ܲ����2(�'N����q��G��a�>�+����'��Ξ�Μ�#P��l���#RF=�s�;w����Rp���g~�K_5�R����7�d%��{��.r�)����w�_��_��������eٲe^�c�*����j��p��tu0�����D�;'s���0�4����g�>���k<R�P�HE�A���
�S�N&ȳ�g;�z��ք�lP�k�q
e*���Y�Mo�k�'/2m�
̰ط�����,Լ���o�.�WRm����3�a3���dE�և��;��W�$:H����KA(]��E�h�(���"S����Rm"^��!w���8���1�Klߢ-V3b%��#�+��ǖ0��=zܷrp6`�v����`x��4��>yr�<7O�q!n�b;Cl� H˳�`˫$A�,��+\������P��'[d�<2���ީ	NJ�\�*X)��#q��~�@|�u�Lqͷ�|��}7���������?�?������?��?��4���<6S3�Kg�~��أ��:��>*#�8LrN#�3��A.!?R�VG}J��OwGe�dFxN���<�7(�ŌI������S�đ�8h01�01]����Ձ���W�@}u�%N6���:;0���
0��Y�x~Y�hA|�`��L/j���I	�3\�O�U�ংR�Xz'<��(�A48���-�f0!:	��'��]���7�T,X�6�)��b��)�yVt���¬)3��$\'���8t�xٽ�`9��X9y��h��>��aʦdδ��e�	qfǧ��+���iP>�J2_�:z�D9r�P�?s'�y����g�)�WU����O��,?��-;���w�Q��.�Y`�����T�ݳ��ܾ��D�<��?x_՞�l�2�K_����K<�
�|�왒W|�DB>�����W`\Y��`*k���
Y����7�{��5?�0�����6h��y�3&ϕ?���&L�V�\	t2�ʣ�Ҋ�2�AZ.��D���v����[��hȨ�4�qy��R4^IRm<�U�����%y�#����;v�W^~�|���W�������_�u���Z^z�e����)�W�7��3P?x��;�Y�lTU"Ξ&I2f=�4Q��5��M������C8]R����ӽ��hرq��4NL4����ǗѮs�r$#(`H\� ?dD�������9o%�Z��Ο[n^ss�����w�Q��~��|[�by�>e�
S5Vf5P�����FW�l��㳝�&��*���|.��{j9q�l9,e��*贸���*ހ�A��Qp/3#(��Sxv����*[�{�ǈB�'���0�B��B
�/�>�}�3�t�1CC�p�g�H=5{�D9v�p9~⨅����릪^J9�O{O�r��Y|�6�>w�20<z�D9���	<��h�v�X<X�n���7��Jc���jx�ӵ�t$��{��/��|+!����={�xW��˖��|�l���M�fϱ�t�2��@_*��c���C|��>�l�v�������;���p�����q��D9uF�L-��rBY�������س���>z\�洷/�����x����?)?��˛o�]vIy=���-�n�r˾\>��a4�ܟ�}�voSȏJp�7�h?ܗ����=&y�Y�E�����c9��yw��!�p�lUxRQ2_�\����: |��p"���BVJ&#/�T��gd���Ⱦr� ?�7�3``��{�{�̤L��9>�{��W���[�Vm�}���Y���|��11?�V4�E;`V�g�2OB��N|=�V��0��߇��9�?#�����/������ �t���Z���]��<E6�x�J����<�K}�Ɵh���}�[�
rf.��]w�%?�4��� :@}�M��(����s�[�w4(����IK��g��m+�4����&Հ(�_W?�tI]�(g�ύ4P@]
}�u���Rp_)�?�Ry]���G�!.t��^�/�q }�:�q�]���4���Fza���|����}�h�yT��UՇ���M�w�	�S�IhN�g��"%�ƚ���C��	��*��og�I�8U r�����S�:���c�-�E�%�Y6`0:;��e4z�O�I�*@�.^��ޡ���1��Qg��I�uDrg��9
��<HX�as���C��I���~�e���`g"�fB�>
��O�2���2��{`\�ȵV����}�69��^Ξ�������|Bu�ځr�x\��1EJ�Hw�ND�<�-z��))�'N����+��Y	@�/�޳�lٺU��Q�Ii6Ak@v�0�ǻa��O�|�'0�1��@nΩ}ry�^����Ce��eRjWH�,*�I��=��I궥�!G����C�ϕ]|b��	b�H\�S�����=RtY��]�l�S�n�+��P9xXJ�p��CR����G��c���C�D�a�9���4h�"}���}���o�[�}����- �f���˭kזx���Tsk��o���Z��9�̧`9��uiG��3sJ�ć~@w&*��!��i��GiFvC���n y��t(s�P��<1C�L�;1�%��$�l�R'�-�5b��^�[I�"J��+�X2/^f�i9�_ŀ���W���>Z4�6s��"nt�~�]�e?�	_���c��8ot��]��HW���e��ə��M�U�f�����*�L���+�~݄���O�1���7y�a�L;���T_���A��R��<�7; /]��-"���vp�D�п�s8m�)�L��e����-$P��t"	�"�:A8�u��I�3g�V�)RbO�ݻ��]�v����I�C�X�)����;�m�ԿH�;�D�*��`	�CT�G��	Ԡ;1�	�ׁ�4�;t��L:~�}�'��Y"k��%0bC�4+�� F�4�sV�8�Rgl��{ �E}����k��7So��������3N&ԳN��O�hԉ~K��3+,Jꮝ������y�Ip�#�r۽{�:�����GeV$(��f������A��c4�Bx���~� \���	/��@��������I�֭����;�N�{���ݻ�1;W��K�DU�r�LѻR�NxT�Z��1�.p�����V=�1�+���¥!Z˵�ځ��@�$Iy:t�Hٽw�����˖�:1dUF�g��{����``��o���Wr]����<ɨJ�Y�Y�y!t���G���{˦���w�]_�z��Ѻ�e���R*�J�=�r8SN�?�O{�W�2W������-�s��r�,����۟�������Ͻ偻�_{�5_/5k�r׽��{�Geq�n���g�:�Y��8��~�3V�"��4��J6Eiﺒ��b�p��2!��-��}�'B�C[�Hҏ.��[�rv�Y�-7��Z������3g���+K�f3[4]��^��PB�� ���G���#��?�/�����,�G�zՏ�劰�r���;���k6�'�SɇM�+1�C�<ƞ�g��}�(��E��J;FVp�*_�<'�k�A��P,>Y���]�l�Z%/�J�}���T6�7���zH�Ğu�{;�h0}u0a N~#y6.�5�˟Lr��Pyq��/h|B�6�V�?��N-]��zѪU�K��Y V���\k�.������T~h��vM^*�Kv�vҐ���d�sc�a�d�8g��h\��u�������.@kו��e�N���.�]��%t3�0�+�{�yU�M�@8���=�(�̘�·�{8= /�	�sb�(���G�03��w{>����䵅�`�Iœ�*� Ln�yMYs�-��%\��������S�$��:zfm	�&���ۡ�����|�77fO�1f�r�]a��ۊyG�kcX/����S��n���m,�ݨ�`mW��_K��dy�������%K}/,�'nO�c�So���:I>20�,_�R��h9v�+��>-����Uf�jPy�l9q���k�Ω�����m��u���D��8���[�l7�12[�R���	�w�?�����y���' ���0�[�(`"�=8�3�LE
�*g�v�r�
����E��
�]��ů#�W�qx��0hFi�ޓ��,��)��0K<�%�"N-�%�9���I#��>��U�,!#J���{��;x��K/z)��j����Y�f�;%�7n�P�o�&�ɲ�������\��*,��Ǜ6��^�<��s*�cvCٌ�@W`C�l���u3k)�!��T��s�b:͘MbҢ�j���8PR���&��u�į�@�K��
.�ꤢkew�L�Uf[��`�q�~�>w�Ϟ5[mga��W1+N9�f����>�w8�.d�;���=cQ�{�d�P0��M�J�Gؗ�pt�Jo��΀�;�tؕ��>���r�]�L�2�,рO�r��xொ�e�P��2a�
=m�������<�O�#<�u9�$��'�S��%�'�{?�>��r�<ö�&��ÀaH��$��n*�뱞����"���u�隷������2Ӆ�}��2��`��y�w�E��t�Ӌ�.�X�ց�~�l�ue��5j#ӭ�r';�p!��Ug�-��.���̙Ö��։$CG~t�A��p�5�@�Ao�IK�'�68Oa���|pg�A������o��$��1Xb�I��/36;w�-�>󬯮��ϜNO�&���$�z��O��?)wK0s]���	1������g%�8|�K�z��G�����\d�,p�7Ȝ3�q ��*�p�L����}�{e����ҙ�T<��`�94H�S)�����o~�˷�w�|F'�s2��
�=}qj{֬Rf)���gO�.'T��ĳ��f�U)�D���|�E�2�a��A�ǘ5�|B@�͜w���.~�ǈҵ�&�	Y~�`��O&���Q4��[�o��:�i��Qy��P�Dko�ͷ�0p���<��o�������j����y6����]�˅Ӥ$�)35��&�ٲs� �YQ�i�(Q��D�!Py�ˈ�5�cv����Uz��u�?*ǏR;Fh	Yz�
R4��r�4A�F�r�� �P��Q�����{�ycfn�hf���O��Sg��W_-�v�B���EE��ek�B)'�W��so��b�>��� ��U7ܰJ<�`�q+�\Ih�]� �q�A�9 /8�|��Q��̸3|�x�����+套_,}��i��r��ַ�^n��F�_x�o7�i����p�c	���!��72<���呇.+V����GqfI�*�����O�#������⋳�kȧ,�,�:�p�m�f��em E���A�EIƪ\�oL���3ѯԺBib:	��sw��ثB&=��1q7�U��8��G����R��=�pl5���Ӄ�6h��Ǜ��

:�݀ӫq�9�
tF�/��s�S{�hzx~�/��>tX�	�r6��}(�����k�@~b����Po��,�6��A��``-�
����3��C`���ÏCaF�#U�_m#����!󄙈�|�8I_1Y'?�s�����eA�^�1c V/PHY�w�r'�Y�vǳйb����b.�R>�1�����E�)��B�'
�#���"ʞ}�;�^�{NIye2`�t&�� ��/ȼ�l�R[f�}���A|��� �Yk>��Y�֓穔��n ~�eI�¡ ҟ�կ������O��?aĈ>�Pv?x�C4ٱkOy������=_6K�%R3J�Tva>�0_��G��yowq�1�p������_���c�Ł0�P�ΘVn������������h��P��f�X�����'��c��U���z�_��]�f�P%w�R�Y�}�GʓO~�<�������{t^c:�,��ǎ�s�h�t8��l���ˬ�9u���{���y�x�O|�Y�����Lq �m��_X;py��*�q�0�*F���`2:ZEӸ����_C0�c�6�!)<;�L.�PtWK��ᆛ��.���wj3'���n,_���,12���^�� ��v�0)�(�5�?��W�I�e,�1���ܵ{WٰiSy旿�pۢ��a���@]�F�^K+�tz*���<����	�%d�av���iq�';�P�Yn���l��[|��'� ���K/J��t�
�6%f�.ZZ�.��H�j�=C|P;�P��!�6~F�/t0�@Q�%��~p��&��Kᝢ��XƧ��Q����\�/��+�888C2rɒ��'��/<�ڹ��b�Q��,˖.�Ud�O�����1�
����|��s�{Ty��:�}`����������?V%yv�e,[��%�1"CQ��-8�p��,'�;wΜ�r��r�v�J���P�X�ә��N�<r�,�]��i�tL\$"�Ca%��)�/�F?�W���K�,���I��$�\�Ȍ^��f��G|9�˾ԯ����1����D�Q����j�R�^�M���̪����C�W�~򓟸�۷�4��2���G��;��LZW��V�E�#M� yT��.!�J��q�4�x��p��-�r�`�ήL���#0_ez���gt��P��{�)���a��A�D�������1�" �'�.�:"�y �g��슧�g�I�)��-+2V�?e1���U��'Vܙ�cf����'�$��Wq���Q|�yad7���7�$Os�Q�~���W^}��L� �$�%�e���$����)����#��!�O�e��X}A.�a@�}��}*x箽��>�Bٲy�#>24��BV�,�02X�j���;
�|Z�ƃꆧwܥ���[n��\��'�Q��2@t�(�|���'xQXS�<z8>yG�i�gG�<�&��
��Dft�����S_���S�(h:~1�@���/ً|�9z����p���3��H��S�]�JK^����˺��?6.��\�r2.@9��8[h��(��LFG�h�����R�l�i�����������^��zK�a�r��� ���N^P�d��;�2ˬ(|t�U�O��#,q_�Q:�At�B��_�	3̊�߰��/Y���-�d\�T>,��ot��)��:@������p	�Е��ь��tfh+�� ����._��|�������[>���^�,C��!���z�yR����sP�Y���)^�G���7���4p�򢇢�C��k�O�R��|��F9��l#� �mذN�KNQ��4�Yk��g���Mĵt�z��V�QT���`" �H3 ��7���m�������g�����~Y~���m�U�(����$��J��Ix�,�>���<љ���'K�w�uWY�<�Y� ��1c�ם>�
B̼E�}��j/So�Ó���Ŋ'�C��5$�R껐p��s��䥫q��Cz~ �|F�}خ����)ܺ��4��F� [�):���V��[*>Λ�u���w1ǻ�;��%�T�=�L��\P�)�T��w�y������W^v�� �ʮʕ:��$��s����qUo�v�3���z�=�V����rd���O��ոg8ހ({�B)t�zEz<����]�o;aC��^�N�	�ɖ(d����.��f9����ɿ�u� 7fSQ|�Q�����l-z�2���rmzhg��K��
oє\�,�K��-�֬�y���Ϝ.�f�t8d8���8,Z@��}��ҥK,���������e��K\�
�!�X�'m�?Bٍ�i�I�QO(�(�+���L������'�x��]R�=x�hٵ{_y����}tfv�D��CfU��M%�Ŏ7�J�OB\8"��չ!�\^'�������N��!ݓ'���rw-�f�%B�f��� �C ��8 d*/���6w�>��C̷�Z"FD���,�a����Μ��N4�"1s�o�^�z]�*��*��]<.E�JK�"Y���^CI(o��;�Úq���+��q�0.,0�������(��孅�-3���D����7�o��_�U�*�����3;WV�\�����%��NX�_;w�,8,.�=�.�%А7��I��!l�r�*���mf٢�e��r��~���8�ĩ$D!�j`��
��Ӡpx����*z=G�=�����O��,����s���r�wze���kw��4h��KV�#�9W�%��>KJ�lɇ�]��2�2��p�Fy�E����ȴӢ%z��Г������X�-R�������sq;[ZΞ�W����F�d2���<I��[��2E�0i��[֬-���o�;n�M���AD�T�ٟ�i���w�&������&@��aǰ[A�/��At��Q����d��Q�L�C<^�zƇ:�qJ�FXb��#���+��Y'b����"�a�{�l4�*���K����Ė1�.��!��w8#�Q�����@����[2\����(>��?�Vz�x�f�U��WS�������A(��Or���ܾcGy����~�}+��Y��'Ȋx,c�G:��������顯NI&�ve9 Ԡ���Pv�*L�	ZI�9�>4 w�;<�8�9X�����gndV5� �]�rp{�C�$ݠ�D"I����@t+��{�	=��^%�r=�i��(eTB�4 r��8�H?����;�f�_�;�)�I�z;�t6&8!��SO���K�!��@�8}Q@яP��h˿iO�#���K�?˾hG�Rψ�A��������?!:��qԸ2k�}
_�`S�V	{��,tL��bw�� �� ��p�ر��U���SP&#��3�s�fV途C� �L-���4;��9¬K.d�=��>���0�i�C� �䫉��1C�q�Ca	�Fz��I�c�>�v��)x��E�=���&w*�)�?������5_)�  89L|�X���K���b�$p��0��qT�~錢�� ������0/�Oњb`�l+�����P"����VOX9c?�?u�Q;K�|�e�UVa�f�����k���V�]���{���i���޻�z�%�C�(�(_j�(���t�A�8H��Ot0���T�r��"�"�,�Oݠ}(Gi\hr{�t�Z�3(|$F������.h  OΞ����(��?j����Þ�=y��]�L8&9s�~Ν�덒��>|Hv�Hn�>)�v�
1ݡC�[f��iY�re���ˢ�U�G��s8y�l�fʉ-?�H���{<�;[���j�^���n��O~b�3����䣵x�9��a��G6�|�h�A�Z�p��@@�rAE�����+�#r��6�!�^�fu��;�Þq$ڏÅ����ϒ���QP��0���U)�0��̠#�>���qx�:*��i����W�^�!0�#o~���X顬\qÞ�qΪ�LT��D�%ۏ�?��p��Ѳe��_1����i#m��Q�"�&�����7a�aH7���I ��`J���q`籺���$؞����q��&1�}�Gu��M?��	;�D�Z�eO�g(��ag�����w2�,{���AY8~Ғ[@���e�$.h�/%��©ݲ�t�Ҳp�B�)�E��/j�P�B��y���_�����k�ِG����J�0�/����H�i�p�U�$��2����{��I�]��r'����˶�۬�2�M���U���|(Kf(��D�sJE0���hO/����nQ�` �Iۗ�Kpfc#���6�&{���0��Q@Ł&�L���V>81-�e9s�|9~��˹�_��y�5�K|����Pv�k\���T�]�@e�yQ���r����A���~��\��K���;Fє.�%<��ІOz��3c�ŋ�׀q%�y�X٥������R�Ny�j���4͓���,[�Duv����I�s(v\��^s������;:�R�7K�ڸa}ٴq�u��Ȩ���p���8���0�='�=�*�u>�л���4Ν��*%潕l?`&�m���f�D0�p8������Y���I�3��v�PT���y)��Ok�p�͓'�o���b�.�3���	\d�w�6jf	ɉ�u�E�����pҞ�7�`.g!�)32�M&+�A�]nph�33�;���W�������8-d��+3���)�V���W.�a"<��(�|j�&)ܕ>�u��'��2���b��{���S\�� c�5��1�o��yُ������aO�������D	�.i��	ZbY�)������(���N㊰�G(��Ͱ�1z�L����<zD�%�Gy�[�!/��7�R�G�IK�s7ԛ�]��F1�`#{�w�ڭ88X�?&�hYG��R����zF�R�	�� �u�:ҭ>5Ͻ�TA�?=�qi�LD�{����5��#?�c{����a���jG���ϊ(y��U�xz���T"[pzMZNO�[�R�2I�tˌ:H\�&�>b��ee�d3���C\�qI~ϟ?�zv�׏��֛�/��/���	J&<L��N<f����%t�:��)���`��-(�肓*�܉yR��W�I�e�e��43���	��y�*;J.�h�"/��w�l�z˭�5�b�!�U�__֮][֬����e�\�RLa*�F��� 4�Q���TEҹo��A��@6X��v�S�]���iv����~B3[
._���b1��� Ƴ%�Bd�a�걤1
�<���%lb�W����������o��0dW��(ǸXC�Է"��s~�`I���[q�3��=�Ƭ����k���=y�ܰE!�{�.)��%NXYe�3�+  ��IDATKn���$��R��Eܵkg��Ï�j��ۤH��"���J$f`P�?��?�nm^���l��;��_[�m\pXc�-��VQjQ c%'���ˮS��/|]j�u�%�(�(4�|û؟�o xs=W���)0X`������'%��(i`��gnq@��,��X���\�l�gi���C�� �]>��(� ���;��g�9�V1ʔ��������/n���lr|=T�	� ���Se��������{���<��v������ �!.+�UID��\��w�1��D�U��~��v���5w�4���/��?~�~��v�����t�=��ᇎ�C�O���1(>۞�fE�\�B��X��6�;�[�F9gP���ZH���l��nW�&}���B�׀�;�ν��~��BR3}�`+����%6�s*g��	+I�b?կgr�L������[k��M�
=�F�`F�L�2Z�'h���=�J�:��3�1�ǖ8��� ������Y�⠭?l��[��W_���?����I��.��,�~�ϧim�{�J���^�e�e��>/�Vv5�C�e���Z�  !F4�p0�Q8MlC��imF���{��~<����~�{�ϧ��u@�*����;��o��&�0fy��T
1��I������` ��64'����n�z��O%*?�yL�f6X���(�ޔ>%f�ċ¾b��0��1����bf�%ɨ Ag�i��]W���]��31{�:�+�K�o�d�J�r)G�4��ޭ
�q��Kߧc�|��������ƀ�ƞT�l㯽��b�a���������a���v����|<M�{�b���ڹ�|�y��|h�7���X��#��X��Γk�P��t�w���>F�h��}( �?��	aωjܹO��P�ؘ+Jz��!Fr�̜5]~�)�q3���(�����Zٕ�̬/3��֞<����)��N��.��'$?�>n��X� 2@Ϳ�'��$ +H�72lC6I!A9G��?��Z�!c6��3Q���g�}����;�c��9:L�ޱK�90�F�4�d��Ϊ{v��;h_���a��3{�D{����ՇtiJ��?ϧf��<E�E�g3��}-�/�<؟�<�?��([<����0&M�2w����_}�＿2���i��w��<�/��>0��`�{��Qx�cf5de�FI���\8�6��l�.pȳ��u�a��NC�Yd�&[�����@�4�ޞ��i��4&���7�F8��c���'��� /��>
[��?�0��*�=&o[{`�fϷ�:f�%13&;�����U.��y���]�U�̎rK
���A��v�� C8S�y��n�����{�̍[�.��W�ME�|P@~]�fg�І��K`�{E�v��?�?�3�ʯ	���;o�S>Z�m�U~����W_{�WG����历�D�2�3�-�pṚ������?���HB�>�fTO&���A��SҊ����^�aIj玝�G?�ayY#�2z���v0z�8�!�q	���Rf�W�0���r�Mht�f36�c�:�Y��O�:/�)Ο7��\�\#��|�ږ�7�c�l��N�N�����W�J h �*Kj��Ё!�ď��<'<�Z�e�T�(�-L6���O�)hi���]��_
�Q�>��aG�� w��>�����3J�����-���(��o�ي��j�����{+�d�K����C{�mOG�R��d?����o,{w�u����k��rbR,L%`�N�[@h���P�H��ƌi�5;A�=ٻ@b�m��=��-[nH�#���K�t� A_֏�٠�e�u�p����`&��8�pN�ĩ����ŋ|]
�F>}�3
���R�9t"�)B���XK��&_(F�!J�d���r�<���?w�Γ����r`2��ޠ�Ӝ�e�5�@\/���\+�9���x��C�Tf�Y�d s^JL|�~�$��e�	�x��F�e"l��}�������vG���;���}�a�\��J����q��v�/�-�ÿJ��$d'���'@ �Jw��5�"][ǂ��3��.|>c��W������s�����϶�O���?i�wA�@~��`��<Ο0 9x�@�����/~�3����0��N��tKR����Z���{��v�;��姧���z����z;z�D�EgXA�r��=�m�x��vi��1c PW�u�é��[�bK����]�p�*Y�ƀ�!s�tm�p�g9X�D���W��[d��{���d�6d�Ӗ=D�Qz��t�)|������9�ol���a�FJ/�]�����Iǘ���\9�R-s�:��7y��:ɯ9�	��ڮx��͞���f�=�B��o��?hF<������#G�Y�D�"���'�B8G���M!��QD� ���)�o}����=��t���F� |� qP��$(3Un�`�X���%�JF(�f`��L��
C��s��'ۇ=�����5�sp��_��M�FN,B��󢃡rr��N�mT��N���1��'�%`��#��Qо���f�t�j�n4���(�/'�c�Q�	�;�����]֡��w��̣���P��`Cae�o���W�����ݻ����=�::%�Ψ��=cF�=�|a��=�|-V-N�!�*:\�H*IK+��Em� Heoh ��L�꽡�#n�A}q��lr����#t:цy�-1��hG9Gǂ��J3
;�uW����:(d&>��O�9kœN���6_4B'�=�C�>й1#�lIlI��[���<�+Dl�"__&g�Bq��m[�Ow���Ŵ%K�5����<о�5�5k��V�pw-sR�N9#�~�����Dv�HP>�}@��
/��l5��ERؗJ>2K�,E�G� �G�a�Ù|G���v{@����{�e�0��⤾:���m�E���O�ֳ��4�C�av�ĩg�@~��[z0��8Z
;^v}{(C��v�Uf�8���Ǜd���ct��ᡅҤ�������NE,�j�N���뱇�9�A�{�����݃�j�[���_5<y���q!���&?��F�e"�dL{(�V�����b�i��&k��,;x��"ҷR/D	6}�K�I�~�=d>+K�;����ú���2|L�![2}���2&���1��4M]�"�9���<F 3� ����*&S��a�礐m��j����'�>�K��"�$&Ď���� n���ʗ�e?�կ�Rb�yS>���X4w��{E|��(��N�ȝm|���������`$�->����5����;#�-��p���.S�tB��#�%���/i�899KG�p~�&!�;ܨ<{���Fd�WH�x��פqG�8�_G �͘�B<�?0��Ը�
%��%���2Ã��>�?��l��w�=����v�O(g̔"��+��M,� �6���4P&V2���1k���ޚ�}�qZ<��2�r[��^u��#�����m۶�w�y��r� ��%xf%�7�����<+��7׸q%�dO4wP.^��(��Y���F��La\��'nc�����R������]�H�BČ-7�tSܛ��������ffh������k��R>x�}��YRf�a�`oԥN*�L�8�������٨���ԙ����wn	�#Ts��w*N+ ;��$�~('��ލD��4	��]�-2�8��B�/�xkܓ"��5�,�h�І�	~G�$���e�ϵLF�h�k�>��2��ʦ�3�v��0��$2hL���Ҫ��Q�`m���w����2ȁE� �P�c�x�	�1f��<���4����P�IO��fܣ ]ym�/�K*���P=q@k�t��P�ϑ�s��o��3Kd��cfB-2Z`T@Z�� �9�O��F�4Ah�9s����^���q�������h�=S�C��>G�D��`&{t~�P�)�!����Cfh$����|��p&&|��K'#U�Gb�
3f�ڪ6LQb�]��~����zT]S�~%����ˣopyp����x�ʏK���7�(��P����OHx�͔�t�W���\�uF
L\hnAia�B��:$x�i�irHzP�P$��%�2�E��`��|pMPD,�q���|PvK�&��|����U`���W��B� ����e��l��T:V̐�s��Ox��;��;�-
2y��'nSEW.׺u�����Ν�-��O��V�n���,�7��mc(���WJ$��"�����������Q�r$��r�r��!W�^�@��DN %ʌ�0Qx��\�4:�P~Q�P���@�Ʉī��4!�2����s������Q~GB�����xv�n��ۆA9ak����	�Is��#�N��?E��	�W((�D���U�(::�N|��-�:��[�FF�B�0Z~�9��@�ҍ�� {=(�s�'J���O�"Q�leS��� �����hc����`�����}�Ȥ��'�O�2��z���z��({�c:�o�ϛ7�3|~�����˿�7������˟��?����#�������D�_���R�������=sև?�B7=&#�1�֠�g�d�WC�?!�8��(qP���B9��:�#��è&PDX�mg��+�H/H�G�!���8Wɣ�3:�%�z���2����B,�L�yM���A�{Ih��B��qV�|9��Nj���'�.�&=��σ�u�͋�E����R��Qv�G���s-%�U
VS�1��p".��r[�ɓ\��FQr���ճ0*P4YQ�uzmm�����xY���±㦏��^�\a��3��G�]��2]Ֆi�3�|�M,�|#�Rx��}+���߂����.�.���t	���U�(�la� �`F�C�|��3p��b���v� �^fgʅ���_��;0�捅��e�
g	��(_����O����M>�1��ԁ�\R~"P@��D�=�/�˶�&��;�R�t������O���?�I�*�0����T7���d��(���r��7�!�I��ڶ�@�w��s��0c�� �L[_�a|,N�/�P0H��2B	��`L~*O���_�zrCX�0Lھ+(���C򣵷�-PK2i��� ;�� ����/&�PS��6�������^ډ���oD�	g���*�ؑ��Ȑ�r��@����H�6m3iK$|ƛ�sN2�{dV���}P�I��'!7�~N��*���:�Ʉ=)��ϑ�P��L�g��l&Kqq����w�{����?/?��}��g?�Yy����90+H�K�§F����їY����t9�2i:ە�A��Yء�E���q�9P�&-C�%~�q�
��iߵx�{v��gd�,^"�~��=�����;��<�/q�k�<�]��(8f�x�b��~�~(X+�� ��w��Ap%��(h�����pgo5�:X҆�'�� �i�5( [�<������D6 ��4���i��Kcd�2𯇴������L�Pft <c�o�+x�����r��ܨ�Ξ��
�S���H>���;i��OZb����&�P�|k�c�?^��N�3���w�2㊙�n�"�Ӧނ��n�!O�'�l'W�z���&~�;i���e��G,o%^�[��v���?�r�=rX
�ֲa�:)�;�����3���J��טm�Q�Y�ڷw����q�>���"�R�ŝ�C~(�ki���!cx0��>]��]��rl��v�8��~I:"n���[�?��=�Έ:ˏj��f�N9vm�$F�Vw�ao ��2�g�T������$3B��.�7qM�}=L���g�u���f{�~e0 ���h7n;Wջ���@+dUG���qо"�aZ�b�"N�>M �]�q��D�y��i�5�bV׼5�,d2���@C������"!�����zeUv�#d����U��!��G=d�qg�����H�b�s��ں@��;��z#��P�Ơ���?}�Xe���4�(b�@f�����4��!T}eNŸ>縗H�䛯�q�5Bwr����oڸɗ��eAǶ	�=���W^y�l��q9r�����l���2��h�tt�b���ٙI�P��)��fE�ԦrT�/�3�9��`�.K�\����rkY{�e��e�Ը�c(
a�o$��?~�Y6��<6@ܸy�X����{19�Mŉ�~ܟ�{�x��v�7�GG�O��a8��	q:{�����4t➁WY���OC�J ���xpE��7x����4*x�"�a*|��+N��yZ���+��c���t��#�7S�>�/�D*+��3��Q�<7�{�S(K�����L�㓗8���Ha���-*w�uwy�����nS��U��KK(I1+��>��I��?�U��j�8�vhz��DkFH�7%��3Z �τ8�(G�B'�G��7�ǻ)>��ӧ�����cG���˶-��f�9hE�F��֊U+Wy�,��p��;��p�<�Q����_ȃ� v�E�(%���kl?#�(�:v�3��}��[����:dϒ�=Gm&��];w�W^zѸ~�GަB�"��E��y)D���V0;�o��_�,�MAD��H�����+�+^Wt'h�@i3펠��h�D?'�3N�[ҫ���b��0N�-a��^Shi����s�m �W�ȃ9��Z���92}33���Qe<�a�^h{��s`|�$q"d\=D��J��K�m�t����?���7�Ze���pV�dGw��q����%u��,���}~�8e��_|�y�Ǜ��n��6���>l�0%昤���`n�B��F��(O�H6&f>�F�+L�0d�/&�3���&�r@<�f:-P_�7�ܤ0"�U���Y�g���Y�t}��t"�r�&�B�n�y�t�~׀���#��\=O[i��-^�]�s<���*
U
��T;����sD���x�`3( K?�)@gI��P��i��%~FQ�+i�ό �A��,��<R ~f���BA�`�)�$(����x(jQk*� e��}R�N�>m���,E3���!-&����E�$Z�x��k�ƞ�S�Z�'�"(�a�؟ @y��)�I3����c"-I'`?�m��O�ic�2)�yH̧J�y�[8���ox; ���ꘘ�e���+W�57��>�s����n][n��7)��LöTx�����[���3�j'�Eif�-������4���SO��~�������a��l� ��S5h:Z6lX������Mo�`��<L,��y��At��Ì���x�����	F��{J�g ��	X���݃��0�w�Y0��o��s���r��By�ޏ�etA�����$��?!}�cr�����|�!�:���d��~"�&�6,���j��2 �D� v�B�Ǩ�o��]��ȸ�?��X�C/�9��<��K�A�I��a&����L��2q�qO�Au z{��6�9�z�iBdR��A��m �L��K���7��� O(��s�P3g(�ݒ`-�TlQ�Ӯ��ⷉ#>��h��8p�e���aF��V��Q�0ilUa��k����(����x6w��A�A�Hk�2��KA^U�Ѯ��a���V�y����>D�y�9�ٗm�+K� �q��_o5Gʥ/؟3�J(i3CE�#��W��@<� ���{��vv�%� n��W��)�Yfn���� ��u��q�d=�j�K;�
�_���� =��":�O r�ʍCk�����5>��17T��UN;f�:W�|�|�ջ5�W�;o���u�]�����y�>�+W�M/_���\�"ܛn�#����r��^�FJ�塇)�>�9 ��l��mQ^�+��2�޻ޟ���;�e��7J�'~=�(0��i��o��4��y��x#�PT;;�0�1��Q�\���w}�D����(�Zp^��q��W��Bx3�� А��$29P��Iw��}�O"w��j>:l�I���}��`��Ą���o���s�@���V�k�֟E��ӿ��Y�� ��;�*8|�b2�qk޵@ܖ��)RhS7��I!���߬}B�8̃|n߅=H{�%fƇ)�i�5�&:yv�0���<�5B��a8b�,p�8FM$���4����p#��N�������7�d�}n���P�l�SyN� {}��x'�
@c\��bB~)@�	�S��1
��=�MBЄ2�B��`�b��"C!�B1�^��P�-^./�4*a�;�S/q_�z�&o?s���7�&��y�A��:V�\�����2�/0����K��颉z寑��� �WR��0i�����@Ad�)��чeRvf�?�U%�w8�w�A���T�(L;|M��0��z+vLa���w���@t� �AXOk��7�r�F���%0��,i:�Yh?��ޖ���*O�!	a�7��ʲ[�c�ٹrN�����e����Ï>(�I�d����y�ɇ�IY�I���ko+��uw���;��.�
�꛹U�N������Ï�{��3Ë-Q����E��n����#�<�m%(��3����O(�|���W^)�����_��ݻ�e5�r�<��; ��jK�)G��x���c�YA<�����>�e�k��#�?����G�_��wB+�����!�5��4��$������ʨs���q��y��}��p �p��;
�x���oҐ8zZӎ�_5����=�bO�}(�^���b���ƿ����BG��ϧ�_�,�Z��4U2*`*:��?	����	�+eڟ��w�C5��U��~�[�B>F��jtkl�-ݝ,��2���L�s�"m���C��[b�ac���:��`�!Ȅ���b/F�ri`6�/3�g�O>���ci�nQ��y������	�J��� �F�3��@/�x���{�svlp�J���َ�uê�#^����~�.!�HLp>����ՀӐI]@��^ʕ�����p��)e欙>����-W���Há����|sh��t���2�^V�n�'�����0OGa��ޤ�m�zv�Yg|�5��Y���3�]���7������g�L��=cQ6�rh��9��6���������tW�̦+��g�y�s/�cp�  ����#�-�e=����{�����e�G�|��՘�E��1{nY0��Ŗ�˯/7��V�(v���G�}�=T���/]�\rd��A�9�{�g:N�ہ0��_������i��g�)��n9�2����e�+�P>g^1�Y�����̧z3�Apݡ�\mꉃ&޴u):��$�.��<1�ꖯ�_����e���`��i�1�0.3cx�0i�l�<�c ��W@��Kl�1���Z����Հ�(R(�@\{�pC.�	m]���O�R)m��v�@+�M� �F�a��?� y��AJ-y�ؔdȜa _��eQ~����.�n�����x�!�CY�4�v=�݄JC�)}q�,�IN���2���
�,f�j�t>��g
��G����PN*γδﲝ3C�_zR��X�JzL[�9��#j�Z��6t����P�0X	Ə
B�PŎG��3�
e&Fd(aV`鼬��`��}`���"k��ŗ�����,)���|��z�b�j�}�X���r���Qj��cOE	��`�,{���DH�����0�:x�*�	�}�)xrR�:���!�`���'�4ƥ=5��DB��/%���(�l1�f�.s��s���(�G�2}��Y(�j�.��zg��Ɇ	<�>�CpR���c �v
���ל�8@=ˁ�0y��kt��1�F1Y���Ѷ��8�j!Z�*x�=�'��+~����0g,�ط�w�޲u�q���^
ﺏ>,[6���\�xN���8��6�̙��,���,]��,]�J��V��_Z��Y�v2_m����gW)�z��nܸ��������-/��Ry��6���/ ��zݴ,;x�{*�q%�ݖC�\Կ�����]��#��	X�\��:c���(��`���~L���m�_mJ����w��A�	��M��&B�����-�2*,ic�'�?a�6�$0��7��7�'6��`M7��G��+��]\�[<g�Qց��߇	
�[H��H�,����{����{n▋M��Mn#��a�-^	���3��}(�+��%����
�4So�S��e" A(��0�{^k>��S�ţ6ε���	�d�}6��l�0��4u�W��f�1��8�Ǡ�~��uz� b�}���ط��<9ͤ#�|����Hp�VtA�\�[��_�S��(f� :o���c�;'&���A�r��YѸ���>�;��H�lP������`0�-:*�`�r
��|��#�t�3t����< Y ������5�&�������NSAv�oM:��3gs��
�Q��B����Z �Zw�:��A���]Y�v+iRv�<I��:}�Ry�n�τ6��sB���Q�}?��m|�:�O�z ��K}�
͍�]4{o*@�B�1���c�-ȥ���>�Y�,)��	���1H�;�+��x�	n(�;��=*����mz�3�Q�O�9.�Mz\��ҍb����Q�xE1#�ȃ�c�@�*���O�G��P�o��`�'���#�v)���P�v7��B���"h(�S,�xG�dV����e���R:7�7^{����k���/����ؾ�
�ˡG���RFϪ�O���l��/\���7��/G��,<�Ap��vŽ~�z��zy�g�������| �-��"�G8���0P�0�]H�e$F~C�%���Q��ͻ���61��'POa��u��Յ�gD[e���{�������-_��m�M? ���׵��Az�������꼈��j8-����H� �D噲�_�|���d����ГeB�A_�hxU���a�M��VZ@�@��FA���]�Kp?Z�=�p�Q!��=�t��[p���s���DZ]z��z�ą3>����q�7��$F{܁r
��YX#�ʾ�XG_��s%|`��_������L��o*�0)� z}'�&�����0�W�tz	��.-?}4�>�������t�w��=�L2Q�b�c��UH��I�] ^�����j�/p&3h��(�"ѩr ���(< ��cr+�Xn�X>�p����g�~q'F���n��� �<�E��X�3w�n5O�^#���� ��%�S �	0>�3j�\�E1?�43t�7��'$��#~_���95��mT�a�%xžC���D�l*�� D
7��X����5I{ �8V��������W�'���LlyE������@�k��
t���9�B��e��0D'�/���a�-��)Xi�\oE��̠��u.�u���kǲO d2�J@�Xn�<�p{����g]���VY �KVm��co'`�~���������?����JA}�7˦M[��5|~��e�޽�lܴ���޻�_,?�ɏ���_�_������������&%�������y��L�a�d���rj��p)t��<�n�㮃z�1�}|�X����G+���§]ɯ����w��i�
�M<v����{|e_�U�	i��A������Y�m�=� ��HG~f
3tؒ����K�O��y���{B�58
T�w���ɲ_}A����'����O�ߖ{��L��������8HZ3-���A��p}>�_8���L����u��Ϻ�K|,;w���7;w�,G	&�S� 3t|Q������^/ǎ+Ӥ�e��~���?�~y��T�zYN4Z٩�3��B!�hb��a���p7^&�X
D`���&@��T`��?y�f���c������CY���������D@�J�ُMy����)O�>��'c�'ە�h���K�4P[�=�
č�b�JIg�H%Rc
W&W��sg;mΛ�{m�kƬ��ݵE<s������(1kK���X@���3+]& ��`���PMr
ċ0LA�1��/-a/U�W
��oR \��}|�0(��'F-��b��Hư�ل̔�u�ؑ�e�=e���e�έ��e���w�}�<����O~����')�������-?��ʳ������/�{�Y6o�X>�xcټ��m� ީ���
� �=�1�)B �d��x�G^ȧm�.�B�7�9�#���A���'�h�Pq���n�S�Pw��;�G��ѻ������6҆ǎ��V��C����+���i��&{�#��{m�k�ٻ�v�f���Tl�����[��]P��e�P�6]a�!�2�\�ӗ�#��m�k���_�G�LrHj��t>��<ʢ�S�#��MV�?��>�NF�I�~��a�JH�>�5_ w���@�-7G� �n|�̙�0�3m~��vO��U6�(B�6
t>��xH���� �%d<� &�G��w�-���/�O~��ʫ��j�{������k����f/�����41u���V~�������G?,/��bٴiS�3��䅢ʎ	睘dE�����"���}(�0'���q�,y�Y�q1AC�U?���<o�3�����Ә=��3�����aZN�Z �_f�G�Rx�N�=�l��M�����Q���å E:���/l����~@[EM�<�Pa,�k��L�`��F���s���41�U<i��k<��E:�'�2�����ð~C��7�!0�%�����O�O/D��.���hZ�yاs�tG=hq"��{��11ݶ��(E=�XA���@BdQVl�~c��
R��?�!dp~�8+S�����˶��ˇ��*o��Ry���4�F2�=�Rޗ��n�;e��&�r��>|�;vD����ܳJ��܆V+2-4��zkY�q"����I��~Y@�>~Ǫ�}Y#3��ـ����O B�կ�3�=IS����/f qwX�t8���	 k�n���I��-�9J6֕�p�p2��zJ3�=�{��K�*o�x9쮰�Q1ٍ8�W�E�s����k�q,�����z���5��7	���EKWB[�F�_vBN���%VH�ۨ�ۚF�:��נ��w��)�t��$^�簘�U�g p���B�]��[Ӛq���>3Z�.�t�%8/Jn�a��θ��M�P����c!��2��Y�������R��0�/��/������˿�����_���_f|Q����^7��P��3�1k�epu��{�?/����O�g�{p1T�!Y�p5������~�p��*�*�?q<Y&AW`�Z��JQBP:PQ*A�r߀�1y��Pv}��3��Q�P�X��Ff
i�p�p�7��h��n�#{(n9@ȃj�,@��Jf/�������A|�+���?�,�3y�R����r�\��Q2������Pa�%�d)+������I<5�_�<�����HB9c�@8$�&�DB�{n1�U�f��]p������y+gϟP^%��/�RGp��9˻�ƳgOJI�`��r��q���L(���j]���҄�2�v��J��� �F}��C��v��Ν��Q�e�/\I{� �$�'+W��p����钼�h��,;���M�\�4ud|u�"�|_;��o���Q�l�)M|�s��3B���T[1J�CcУ�m�ƪm^,�D�W����j��_�Գ����(�D�Aq��آק3� m��.�t*�-D^"���Xn�&�M���w��:7[�@1�Q�K�x��&��F�b(E,s0%�g�YQ҃t��Ce6���{�[$<�9�6�\Z���0��M0A`چ��	�#�A�:O�<���:8��:��_S�^�)�ua���ɀΖ� ��q����3�_��.&�%�]���`��<I~��>s��:rgF�:����H�`�P�&��*��u>�K};y�d9&������l��+N�(�s�>�+����ɏ����Q���NpaH����̙�tI���^�9s抮�.ϩr���>�t&K�E�� O&�0�g?{��3g�H�1`;�*w)Ҕ��,�(O�PUƞ՝ sȼ��]_ ��v�>M��e�Y!X؂�fAzqM�NFZu-s�:�z"9�v�,W.��@0f2��N��ep��5�Og^���_�'�ϔ�<�ث�ŋ�wyTYR���bf@Ww���A" 'A��b�	,���H��*L�ω�\�"�zlT�cUk������ߊ��y:^"� ��Ο�#�8��ա8��\#$�"O���Oą�X@� �[����dqdy���%���e��Т]��?�����mE���d"��0��pI�PU��&يyv�<m����Ox�:�}�w~�#i���t�?��4�Q 1�Asm'�5���r�>��e�(�N 3Cq�*�L��;d,��_"e�rp-@du�+�0�2�sh@y6b�Ŧ��-��6oX�>�vA}eKm"&�B����4҆�K�r��K�;}&Hg[�%t/��P�4��y�������S�Y�N
�sS"jj@<�&�x�$ �0���3`�j�EV��&_ⓘ��zK��;�9ͻ�y����m�;ﺫ�uϽ���o(,S�c6BbB2�B:!R�G��bJ��=�zY�W Yw!Jы�8��	�hP}Z�p4@w�A*�X1��պ�j�8����4�xRi��x��d�:�l.u��B�
�G�0==�W�N2rDHc�R�;~�;G\��y��y@��E"k6k���v�B����6<	�v|����̲bF9»��mq0��H�D+��ܽSY��]������=�����6�A�8&�H� �G� �a�pF�y)p�w�(�${��s5؈A�t�����R	�$�	�)�J���ʎ2��a������͊*E ޫ�����)�a'�\�Vr1�^oV^�,�;&C)����&L���y�q"�#�H�2�AM�Įa�z�S1�0�#����P ʮ�X괻�۬H!�RfR�I$�D9�HǍ출 �tVY$o�ԇ�Je9''?�`K}ί�����(�iO�
p�-�tXI2}�Qv=���H����7 ��'a����k��WW(��El�?�0P)�����M�c�����a��m3"O5 |��X���3az����؇�:�Y��:��y�L�jy�W�W�}�tE��i������g;��~k�oD_�6�K�D~E��	�mN��U����-m����޸~�w�FL�%�_��2�2�I+��)4���B�r����C�-���6� q
�U����Z�����c����~�|�������^��w�S~G�����������/����W���/��ko+�/�L�V�9=^�����d�M�y� V�j
��&��-z$ry�].VB��F�y9y�j��	��J�@�����g�ʠ'�LF���̏�x\P�H��w�ء�zk����OH�tI����4��u�|�-&�ցJ��9�	P��&jݫϠ�ٯ�Q�����<G��m�p��J#�Xl��1�}f �2�@��0%_$[�r�p��u0����N~Ǳ{,�g� �E8�OVz��Y�C��g{���H���I�*ZWR�Q���A ����q�sy��N^�!�f�W�k�E�2�=[���gx�Aep&7�y�bҮ���NY�+��90�|Rޘ�6�RV�*ɀ4��K�(�m��~N��rNu��>�)'���ò~+�8R�&4��`W:S��܀�����G�UH~�-�%,]�U!į�U\3F�N��J��i֣O�0�Ή�
��1!�[��x��n��.Ka�lBF�G�5�E���;h��ڶ�d[����Ǧ[aA��Z�|��s���������	�l��Wc�ƙ�v8����/�x����K_*�GT���럖���Y���'������������s�;�����A���������
e��w~G�������S����S��~e��c����L(6zEct���2m���Aa<§���(�e/�.t~b�Q1z�0;gy�G�Ud�r�g}!Mh��Κ��������ۘ�5�><��<����?u���q�w�us�� .2p���sN̤$�I���%��v��v[vk�z-{��s���f<v�jK�bs&����ܜs�y�߳k�s��{�� К�~��:w��U�+�:zW48�2���w@C#�ąu�Dݐ?yѠc��:d�M�'�N�سC�����I��%Ơ�7Ǉx9nҤ�@�d(^ۑ�Ϡ8Mby���}��ػo���ڻwo��P=����=�װ��dŭ�.�zF��+��F	m�=էQ~����)�n{�r$���܆�yCiMԳ�X�ElWoQ��jn��u�xS�I6u�{���Ɏ.\pa��|V|��s�ԩ�����c���0��h+�N� ܠ�/��L�:Ո��Q��b�����}��X��3{N���˅�rb.��r�e�������p?�~�e�#:�Ĥ>w��u@�7�}ɩBO;��@Kۉ���Y�����_*��=��.�_=��{/&�4[��F��fLП�5��Z�[�%m(�cFm[�Q�/Ǯ��/��d�}/��R7���mC�I�f_Mz�a!�\�'�a�OV�����m��V���r�]w��W��^|����/(�ϛ������r�Ys�0�.]xq�����Aq�F�r{,�S�{��A]!��uO�߇�G ����g=�����t��\e���4"`���l7�A���A�T�h�j*�(�Ї3��\fp���[��v�#V��]�Q
�4ykR����
���{ë�@ʤO��
���D�d9�;��;���6�ĉ��E�]b��/�0��V��ep#�d6��}�B�> �/��$�p^��/���/�29�N��$t�i��nCPW��/�$��b*�}n>Và�_?Ӆ�qO�~�=~-���~�`�j��+I�Ce�\�[le�ը����ޕ���u'��Rr׬Y�O:/_��lڼ�� L@���(�0]�5k��ӝ;w���^T�{�9_uɧ���������_.���ry�����g�y�<���)O?�ty��O<Q�x�q����|�	�y������m�!+��0�����N�v���Br�d�21j���3 �@f;4�SO?����+�'��Æ�ֆv,å�_��U���r�����8-�3�E7�)��7��G�ⅴڶ���x��ǭ:nf����h�pY���X�T�������7,81��e�c4-�� ?ҁ��5���kˍ7�X,XPΞ=�7,XAU�d _������o��&� ��4Yy�1c�f�̾��K[1����2��<�n�z�*()/�R�#B��e���C��E`�[
[>�����Ui-t(K���
��B�Х3λ����s��00-������.���(;J��]�����q���"�]~�C�C�u��iC���#V�����Wo��$o���ӿb�C�� 7����bp�+=Ђ��v�a+Rw�����o�� ��:���#�ȋiL��PrY�ݻ����NX3�P�i�����	Bs� BE
���0]��AK��Q��>�O��4m��@�s}h�
�)/�qdk�ga(���"��ȳ��0����ي�=�[�m�8^���֢���ի��*��1�8r0�L����e�ʕ�q)������_��_���k���;���B�����/�o��}��W���+_�J��W�R�
~��Ư|���z��T���/
1���/�-����[��V��OR^z�%ߣL�݇��x"��7Uvf���q�"�g��S�!�@��9�N��Ƴ� #q t�B�;�S�^Z�Лp��-���K�n�����o�%�>�1��5��B�����@M+�d��T��~�AD��ҮC�(g�0���Ÿ����%L�������%��+E�wQ}�g�'i���; ����gʃL��}H�&�N�Dw���JU2&�[{�[7�$�΄��c�}�|���*.aY5�Y���N�̹��V<�L���u�V#��cۈ�g׮�~���|ۙ�sv��s�KLF��.TC�H����@��/� *�M[!k�n\%M����g�l���~ <<��(��:f4w���x�)φA�h"���VP��|�;�$a��朳�I��]z�`޸�U^�H$�.������p�158�1�[��<P��{�0ξ��xn���kd�h�J���ۃ�A�_W�G�U�)�IȽ���xS\�]-�o���*>��Q�G	OYE>U>˗\������.��=e���J��I2�;���2ǌ�3��l��Vn�r['%�U�w�n��B�k1J+2<u��:���>��=�״��]�4�ڏꁣʁ��5��t��K�8W~2
L��Đ��F�?/v�܏�o�Pd��a�Tc�ڵ'ې��6L�Pݺ�� �Ѳ��/A�H)@[az��Vj%OȤ�Jw���z\�_�>����ރ՞�熭��W3�u�d6.�?Xvk���HƎ#��}{���;vw��㶈|������˖�5+W�իVW�M7��kW�%Ｃ�e��ur������˗��˗��K����˖-)+W-�����v�P&a׬]#�9tٲe�~�f�S-�l=r��i��C�����Q�mBVh��W��r�B���a�WL�x��*͑rBf#.�f �6R��#%o���r�i]�rP崞�\u��$)��?���4�O�m�m(�2���UL����d�_�w�������ѧur���
�:�ӂp&����d�]h�]GX�"Qe�_�X�=v�%�G�>���8|��=�g�(�g�(�wnYp���[o)w�uW����ˣx�|��)���O�?�[�/����s�<yD��߻���d�B�{��N��{Ƞ?́�z�
�AqT�m"������^}����+套�z�������Kj?�яʏ�����j���w�Yl%�o���-3z+7NVd��K�B�a2|�#t�r�Aa�M�Ӄ�|�2���k��S�'iQ��WϜDf�
�1ˏ�Q�����T��1��ո���|��w�thU�:��'���] |?�.�#}�1�8:���3-Љ�>��
���C�}��S�� 0doʣu�
欹�3�Pp�&�$m�ە�C?�蘎Hɍk�b2e���>�v���kݥ\��ʬ<_�0==4��}xj��-����� �c?�[t�S��(�gMy#L���WP��Fx����V�D��4���+����*+z���2��4&��pI��	������������~�� �&L�?8��<�brɏ�ί�8-���d��R?8_hy�Ϲ�_>��Є�{Cq#,Wϡ��y��>s�� ���l� m�7�H�fq&�Ҍ���-8,w�$2�l�=(r9����vo����v,E�����Xm��n8�ʦ����ɳ�G�������WH�\U�^�f܆�š0��%�߃�UĐ[�չz���*!x��_u#,�B�������@<w�o�ɣ'N�W��%�_7\?�_7L�IH�>MV�[p�[f�T;��c��]w]�Ї>\~�����c}��?W>�{�W>�9����������[��[�㝬��?�񏕏|���;�,����n��0�Ԃ��'k)8>,d��$}��[��42X�,]����W������|���?(��~��������~��Vlq���v��׿�l���?�y*^(�JS(���8u���R�N%��A�!; �uV�/���[�9���8*ω�"�٩�5���We�/Q=fy�-��m�C�v��e����#a)k�%���ic�o�D�;���w�TQ��]5��Y��ޞ�85-�?Ҁ�V�d^���2�Teu:�r�#��W֐3��@M�M��o�i?9��2u��^�b�~�aL���qy$��~��h�9��f����~���]F<~�#m3d���?�'v�XV�|�A�rQ�ׂq�KvVL�zϼ"o���3�G�="3n{��*�u�ܧO�V�=��r����<|��
���#f���'2��<3�d׋���2�s��c��^�\�A����x:��fTˠ-°G{�-�:44ռ�<�f��R4�v󨢟c<Fg�.��e��>���~�	�x���d7�EB5i��T�\��V��n��|�-���g���~���?Q}������ﾻ�z�m���/W]u�o����>����W�262��W�CSXA�0��k��)N2�t��%��tH׮][�z�)�g��_��˷��m)�a�9��^{�,Z�Fy�E·�믿V^}������e��e>ހ�8�lg�S�m`v&�:�K�w2�:�^�����T�� ��C�AS�OG�/���d'j�B	qgV�C9ϚB�B�7�L�B�=��]?$�r�	r��B}* ����?^�D��!�I�c+[I�Lh��$E{����, $y��@�W�3�:a����}/1�ŮW�D0��d]�������S��%�.�_�˳�N��O5λ+�&��>��-�n�Mp�n9�]����B
o�i�k` ���.壺�r�wt�2e�TZ�$��ǁ�Md#��ﾫ|��y��(�Mğ>�A��Օ'�b`�vϞ=^Afq��X��GhVr9~+�U�V|ʞi3Ź���@�{�7�^������
��C֛�U��$��� 0*��e���G�BG�E�::���~B�civ�]�6MhK�N������<�����b3��zO�V�� �}q�ɼy�ʌ�3���زeKY�jUY�b�����[o�%]nyٶ}�Ǿٚ4^r�%��`�ƚ��.Np�!�����>PH��,�A ���N|$�"+�{v�)7m��\�+a�ݻ����&6�M��5���:��q�w6�]���$t�)����-�ς�Ӡ���n`�[n�	��?�2y��weģ��4�@���Tk��(�_��8��Y��p�@��i�.���� �,
c����r8g��m:�ѝsE�)��ͱɍ4�)�r���T�?�����=�
���%a��U^�D\L�7��P)�x5>�d(��^y�τ����)uǙl��7�A>�t����x���1̲�3u�a��5B&�<�aI�Xe��?L���Ӡ�FB��W���M2��vY�Z���"���!�!�q�<�B�?�MO/���:��'���&��c��䒋�=�������c���~��t�M�ʅ��	�:������7삐�0@J̅ޭ�6�q�<׈]u�U�k�.w�q{���{����A���P��.��ѮX���xN�:]0�B�0xO�'�L3�� �m/����;�m	BG�6�*����s(}���E��G�	N�#�2�S�hcN�;I����5V�K8b��}�K��^�����(�Q����?���P�����?���T����?{ѢE�Df|v9X\�,_���\5��}��������G���fw�������Ne�T�a~���$ȋ#q�mˍ)�K�a���CҔ
'c٢��ʙ��)�˅^��Xj���k}�!����'��^��I��QX0-����,��V��B�����)�Ua����v�۫����E���ͧ�]�>����hdA���a��@�!4^Оe�ك�x�܅t�ڻ8ȟ'����a�b|�;��E���� �_���a0������\O�v�!�v	�v�s�Cu�=���e3����vG��L�23�@	��v*u�ʒ�g~3Ж��(�@�����ظU��OؓO����՟w��^�r���>�
Ol�t�x2�	{������xП�e��yS7�=륭����1�eo����s4��7�(`ޅ�E�~&�����CG����'>�[��Dy�(>�@�����.ʜ�s|�&J0�yū�Z(D���c�u�__�����q�V�|�����>������}�C�C������^i��BxN�C;!\�t��>|=�'�DmbY'� ��$��9L�3��oP��n<944��CR��&c����S�����Θ���%��������
�r�Ő��VO~-�?�CO7y�;	�'�;�F��Il'�Y>;p�?�L�zsQy�W������{����~�?�����ޫ���yz���Lb��id|
R�0Q�E 4�L�T��l]>�kk=@�A�vR�Q �D��ʅ��Vj��N�2����Ѽ̆���C\;���ۿGm��5H��]��B��Ng��
>x��w3�1{f���������?�|ur-�����?�O�������͇�ٶ���(k�GGԡr&���U�C�yU�?B�*V'�����,�R��0A�\E������+A�"K��Z���$��@6V]����� �H��f�:ϸt�ܳ�k�.+NX�+�,��'�n��/2�s;H\�>j_uce'��qcǗ������#?S�t� Ux9m޼�$'�4Ba8��ԓ;K��V��/H7�v���b��_(A<���h����-�$ހ<a�i{�W��7�G��>k�)�u�:�[��{`�uǩ��;A(����P��	 �Ƃj�L��s���ka�[�ꉱ��-�w*�T��o8p[� �x��S��T�G��4)=�vs�u�E7.�6��6�)��#;&71�[j0ݱm{ٲi�̭��+���f��.�.��BOx衇����я~�|�3��^���?Z�����@J�m��V�������V��O���?)�����?��X����O�I�g���R��?���_��Y�տ�W�O��O�?��?)���������`���?�(���rES�t��(��p�	�p��?�!{�y��~-�%��t��D���������q���0g��R�Zt+�ūzf���m�ň��>P����@MQ�Wý���TZ����MZ�x	]:0�!�G��B��;?�/�N����2`�U�@��dAD���|��O���x��{מ��/��_{��Y��8pH:}��8̋����=��v�K�a�M�x�H�7�+Z�%�^�o ��y@�;h���$@d�	����i�4����`"�+��F(�6r��
h��-�vv��!	�T�X�ܹ�9���U3�6}��𩚱�_�����-��S�ٍh�⡬R*��3{��l����Җ0�� �9���^}>p<�%��F��U�BKn�'�:G�Џk�ۿj܅An�`�j�n��;;ufj��+��1�'��TCf��8_xS���"	��A7VJ�_�'3��ʼ&*�ܬ��g {����z�������`8��� ��|A-�B��x��k�ȣ� ���?����'Ä��v�1�/^i�_Vd��	���w29��Bt��4{��Y8�.��r�邨t�C���3���ݰM�Lɩ��,�16!�V���*S�Y����!)
��B�9����� ->�j�m�~��Z���:�=:M��z�����M�}����-�ii<�7�|��p��X�Q;��iS�ɔ�q
>���./W^yEYx����]�Z�&�,��j�_�g���2�xt��e>���gx�5/@6��������Y�a�Kg�zȓC����֡��x�e\ �2�A��#�����/<�~%�b�
ų.S�&�2�~��o�w���E}�B�W��0)K@�J��xL�GM���+m�Z�4>�>}�������
�'N�X�N�j���7:�+Lz	����S>A��0@R��a�&s�Q��Nf[�|���i@M�	��Ѓ
�~]N������A
�����+\�,*.o�����+���<�TI1����[���
��wKG�"�'��b׾��-h�׃�:p%d!v���aʊ{�/���3>�$McV��+�ä=$��])H��B)��퀖4�;a���\D�Ӯ<�|����Vv-��V��t\ �S���lB�ʐ�`����`�ߤ���*�]L�.���<���{��<��9�=�Ӄ�e�L��Y�2���9�#NAo`�=�2�ٽ��r���t�Du�����N��1�vQ�j�^H�Tꉏ/q?��2c�tߢ�J�b����[/���b,A�Xq�4y�w
�:�,)���V9��3g�W�䇒c�ܤWt��|��LhN�r��H�Q1?�!!�wH{���C�q��!$�xy�P�MФ@h�4e�4����i�~BO
���>�~vd}M�KǑ�h�0�Ხq��[h�H'��Fo����R��$�/�i��;�s�M�~Cv�^��^v֋/��,��u�����z�����nc`%7��>�#�?��`>�'H��i Dy��&��`et�+l���ͮyN����8!FAl�O[W���J��t4,�O�`x�M7�����j��bq�U\�~}ٰa���Nߟ��'���7��H�!��4<�|����'���"w0�A"3<:��cםw��D��Iz��0G��ˌ������v����lpxt�I��aAq�7E�a�@ֈ��#n�<A�U�S)��|�60nO��!����=;0�f�n���/?4�tz�\?���4 y�E��Y9���c�����8����w��p�:���v�s�r{T��Tj��PXO��B��ئ)I�m���x�z)c|:h/���n?��U�TzO�`���e�����0��x8���/��Ǫ.�"�c(�|Lb������k���V)�g�N[���:8�|j�I�޵2�-���8�c���m�b�k��*a}��1BF�|���>���
�,N7��!�_=�p�b|�B�o�?��"b
�V����4+��_�'�����9�L����sB�]��{�aUJ�E�xf��x�1�T&*NѼm�: ��qA�*]��t�s�
����5��E��G����~�g���������#�<b�#;\T����j1	N^Tte�~B䆅d�邪Eq�,zB ҥ�?��g�ϙ�q�
9�ʑ�M7�m@�À��b���+�7�Sa[6ovGɀ�/����j�]f6=���i�g�~a�>w+�~�@e����a��2,�,+��~th���%�|3o������Ocn�&���@}[�V�	q�0��=��|5<SE�LO����L&�G�-�L��Wq��v���Ӧ�CV��<����A���P���ae冕�9sf��s�4��p^��>ߙz�ye���=�["[դG �g/'N�2-Eņz�װݬOX9������W��)OL$��t _Ђ|�̧p���E������29���o�m���eBۆ��xn���7��U�=�s�چ_����cS���1 ?P����(���N{ N�\�v]��0��cG�&,m��YD>V��G�kũ�i�{�}�8װ�&��3�*�����̲�2���n����©�?��&o��]�P��<���,�(��4m���}a,1>���-����_:�=%�^���￿<�Ѓ����9�D.�-�e��_x�/��؈�ub��A�/A�Y-���>h����ո�
 R>��2�kk׬��'{�����q��E�A�� q� �>#��K{4��' 0� u�T�;=�
�t��9�h�ԽR�ptV(�lC��U^-��刼����!�n��o-���G��[��k9��A��
˩�2c*m��0k^M8c��n�����|�9Z<�8�*� �0I��v,^p̳vɟvfJA4Z��f|L�q�z�S�ע�A�Pg��M��1�&�gC�I: 2h���yl���WjI#�E��G׸�6+e������<�^G�ycii��HA /�� �؋ì�����(5y��r[E�6�]���c��s�-�	��}��1�=Ĥ�E�W�X9$�8[ږ9Wa�*���&!9ڕH~�m�d����8s^�� ��(?2�Eh�K^����/�K_�r�)v^"�ߍAX�Z���$ d
�[{��{�֮���ن��c8��5���Ä��b�����j��1�޸q������K��ē����/�
m�4�'He��#T���F_�4Ʌy����/=2���[/"ȥp#���2�8�l���d��;��?VoӄD�"���H�r�s
kǞ2�ʚ�kO��z��}�0��lK��I�Yt����a�Pf�QB�p�]Σ+l�K�d�N(��Lt�x��|�?�Tah�H3ꕧ��OBD�d���cR�#�삿���ߴi��0ލ��g�f�e%�	�ҥ�ʓO>U~��_��{�m�c1&�$>i	P�JP�!t���Y�c}����zr�V��{������?&��k��m۶Jy/�DF]���V#�f	��F���z!�XQ�����cOsp�C��v.��>cz9o�y^�a�?a��2M���v`�<�W�X��Mלnl��<U���.�
$�yg��X�&�����
��T4aO���Ғc�5}��~�&�>ǤA��wS�����H�!�w�d7 �,�N�x�K��K���l_(��q��3x�˒�a�w+0��@C� �᳡tjT :,dY�,(-d-o �H#��H���.�KG�J��v7z�y���;�_��.�j�rZTw��p�h��%�O�-�~����V�m4�3~L��H9��m�6�f��-VtxQ��Mƍ7�6zm��~\o�bt��v�d�n��@��bnAA�0��+��E���N�A�SvܬnUw���P}��#nUi�ɚ"���>������~�g���;v��`��ݻ_��!��Q��m�Bư%��4��� &�P���to��L���+�	��d�A8h�H_�71xU�eR��;q�=w��1SLW-[()�;���"t�]�Gهத��s�/0�/�]z�]�D���U�d��w�vdOeP=����lQ�r;�t��=� B�`��1���AK���Vp�#�tG�8'�����r��3�Y�+2���tw��ʳ6N`����~��z��{�~���˲�ݶ�+�ƨPv�#1��,@ε�l<oh�N��z��j�6�6����~���3�3��$=����_?�����^���[��,]�L���L���%Kʒ�K���Y~��3�r�O<iE�U^x���(2v���!K�F?0β;�"��b�>�.�����/|��������5k�j��c� l�de��q鄉���)����SE<�B?�&�q*��
0���@m߱��k�����������^/��w�|3�U����٭�b��ߖK���rbu�.**f'U(Dx�qg|Z�>/*?D�}���G&.�ܓ�.P��=V9r���>C֕yU�A�N�v|��R��h��d�Q*"�0�y��b��u�F�L���+&"4h�y�pڂ~^���e�'�X1Ҥ�E]eٙ�x�-:P� ܳ}����]�o(B ��"ϸY������+k�c˖T+��`0�����E�c5�`�3�c��f�5��=gn9���eҤ)�"o��8�
��;Z&T�6ȋ8�fЃ������Lk�@D���݂
�`��RFp��wF;��+�Y�	n�2Y<�~t�g�[������'�,��~��ը��H�^�󽀐��JI_�f���_�u���
=��n��eL<9$Kȡ��o��/x�r�߾�B�2�k*����jG^Y�G�M
%p(]�U��	�c
�IA��H�=��w0YH@qe!a��%套^����>�\y��/x���//��rY�rEٺu�wֹ��t܆��Z�*����p�v�������>aS�j�I��FǊ+#+W�@۶y0� T(�+�Q"�����ܲ
���.+�a�
�(Fo^'o�IX87�����{�=��裏���o��ͫV�.�7o-k�I���Վd>Yg�*�80�`8���������Ӂ6�|
��(9��m��%
"�8
O�`���(I�9g�V����@Z��#��¬J�6�&Mbx�J�Wc<��D�Sل1����ܓ��X
�V:r����@^�������K=7�|�r+]:" 7���m���O�H�I�X!:�EY��ѓ������ ��󉘁�g'x�E2t��|����N]<�Q�TE���\ˎ����Q��N��L)S��V��r޹�k���<p�����D��O}�|_>��ϕO���o��o��#��>X|��r�m���._ %x���u�UB3}a��Aq@����Duy:�r*����$vÈ�.P���0�4 ��8.t��Z��|�{�-?�я<�xd�fy0H�N,�͏�j��i��	2J:�Y��Mf�TR�WBD���Q�~첷�/�����ҋUb�M�v��8�b!��-�V�˙ ���.遠'hJ�Bu�g^S�L�U�bE��@�:��6�o�d%A���N�?V >F�18%��BhE�>Ru��=�6na��[}���]z�e媅W������
���x�M�����܎�ǖ����ZfS�<�h��/�Jl��@9�5�C6��'DB$]��a�Lү	#@1bC!��/{�E��+������+�\� �1��v��s���3˄	�d�����_�.�M���`�y�7������+���m<�X3s�L����o��:��e۶�e���e�;��Nu.� �@%�_�![�:)��t���}и�2�s[ޮ�_ӏ]�)Ƚƫ�aJ�v�D)���貊Y#ٲw\�axQ���ių�7O�x�Ϝ��@�Q~z�.�0�`�$2��Q@<��vUҁieW�n��G���w�&��j�OH���N���6�� ��*���V8n\�q�9��ji�=i� �߁n��aC�P�Z{�ބ����}B�L���Qp�r�c2��"<z�2u�����W,��{]�|���*)�7�tk�����?j���G?Xz�r����{�&�?�hyPa���r�uו.��̚=�L�:��S�8B��%��� D�]^����T �:5H�U$�^ {5���8�G~-t��f��=a�~��%ls��g~]�|�護|�%v�b�����(Z�w��Ga��Z�^��0OX�f)W�@���p��pqҭS�����ה�4V�-0S� ��o��<BVá��!�9�-t�����q��I�p�}3��},~��<^��E�^��\�s�i�*d�xP�p񣫜���We hd����P�5����g����v�5�I��R������������{�_*dG�`7ؓTeg*Eb���us���.@��MP�{�Y������={���G��D?�.�? �x<�DCf���;�p�>�ϔ���Ϸ�r�W\/_p�]Γ�r�=փ2����T�/Z��ʆz��k�ֲaㆲd�����{�Y/�/]�TJ�N���\ޚ5k���2[VD��䉓�,�Uf̜�7�w��Q��۫�|���(�s�l]#����٥9�2�����x6V����3� u�/�)/�$~��Ho8�;���F��Zț�$V�4�cՒs��D��r֘+I�"��NB��Ӗ��I@'3Ƌ/�ą�3�tAgi	:[�P젓zvg#�d�'�?냳z���|㺻�%�L�hYY"�<�ẃ�J+3��� |tB��N�H�̘9#dg�d�#d��L�t�]q�^-�=p�*W��� �3ƛ�l���yG�v�t���x���Y�'�*o�̾���@9P�B��&�x!�l)��_~�������ߜ��ʹ��U�����{���[�����U��LU5v,�;�\p�E�}'���	�_X1&�C�O@k��	O�Q�Z������D���/�L�X��f���̸�t�,�+z����W��OJ�~����ح`t��r����Y�cA�(M�4Q�p��R�%��-�0�Woؓ='���/R��kx����#��nH�>�v9��'�M��bW��/��ݻ�lQ�_�jUٴy������  u�]ރ�����b]Y$��>�/,~�����6��R�݉t�v�d�s׽k�w9�p+�MŐ��_�w'��]�W���8�M�w3�z�8XJ���ۉ�,ǁ�]��h�,�J7�E���t��J�.��އ��*��<Y���缩�J���N��K����]u���g���֟Ӹ�����}^P�����f�����9��4�1�4��St�v�m��+�}�weW
����=(��h��{� ,P��풅�9EULE1�r�s��-��zk��>`%�N����p�68k�,?��Kg8�Q�s�9�̛;����a�_|R�2T�~:����1>)�B޾mG٤����A�Yo,X��k:HW�fֲd"F�}��I��h�9�$���,���`F~�H��'ZH%^��$��{�����`�'�M�|�
^;-�OP�P�h �E�̺Xat�"�<jf���o!�J0:��V��9:8�鈔GL6�V��	舆8z�����_ڦM��I�7&h��L4d����s|*�I���|�P<�^������0��ɟ�t�&A܀�?�����݊����A�J��Й��k�)O���n�y�"���0�7�DW�\Y��X�I�y���pp����u\ׄ���̙*+�{w[��e?:+:�L��&���g[�� zhGt~rq�W��VEt�Ҧ�t0���N~�7��8����U=;��6���B{�+�(������S%k�_pA�����{�5ז�j�ǔ��=��	A��B�}��M�M[����g�n����,��h���e��e���'��S]͞3W��� ϙ{�H�CN�0�B�_�u��s-o�'��_b�#0��r �t���P�Ż\y�$`<_����*^�5-E!)�d��t�_�g7�1�nR� �f����������);�ۭl�ҷf?�����ݲu!��?yg�Y�#D��5�rך��F��@���.픱��ȼ'�&�S\x��m��]B'ÊI+��n�"!�./w�Z��&�8Q�}i(}�����DX��^�|"��c��]��Yv@�o�usM}Hٳ\�^�m�&���=�� ���Oyc����L�����0������x7X���ߠ/ye�D=���Q�kqS�_���1��I�aүy�RyY��<�Q�oj��سo�^�AT-��V�ڱc{9ʮ��!iDc!��C�#o%z��r�uחIR`_{���������?���xy�gʳ�>[��9�>C\�Ќ3=ƠGqs��c��]Y�b���MGUvY@�ca(�3g�P�*�!��%��ͤ?���`<�7�����S8`����a`��A>1��;s�r��]Vx��r�����w#�F�ŕ�G[
I?@� ��(/��9ܽRlxFΞ=�\�ʺ��˭|K4��,U4v���s>f��G�!��
��Qb"Q�S�d����
���@�'�1�`+V�@v��?0#,�t���!~�����=.���l��M�����W0����c�t�*O�.�P��C[�צat=��DX��A�Sw,J��	 ��L��$�q��&'#��s�_��0����2e&}�8q�q�Y�:�\�i��=&P���&o�s�-��c��b�I�9�O۟��-ȗ���CΙw��~�|�����I��;��R_1m�t�-��{{��`E�Dw�٭��`$-L$P�!���>֊��r��ו�﻿�s�C军o-�^pa5nBٹw�(e��.�v�o��6G��L�J�g5&�A�^:�/Y������x�r+ó�:�,���r�m��{ܩ	ɍ7��s�gϙcZL�K&��.Q��
��_>��߆����)�����E��
!!�9m\j�F~�g�G�+_�l��g�c�Mf'>�#Gp�xMzΗ5]&	E����p`n�xDS<��e^G�j��^7�#^ͿMw(v!y�
���t�dO�6���e��kb�fB+�e A]@�ۚ	���>�lÁ)�����O�k̊�FO����4O�|��E�\e�_��p�)�0���Fd.�\Vh�؅(�,�d�&��_�u���Zz��Q�Mm|"J��KOX�&��`�@�b��1�E#��?��0/�2!{��g���������?(?����������HJ�Se�歞����B'��vl���%����V���0���9t#W�I�$ s��(���#��'>Q}��D!�� 
5�8�� [$�+\{4��r���Gm���"M�RХ���PL����I��EȖ�����#>Cb���^@�|���<ܨ�j���7�j��\(L ѳ�=��p$�ТC�� 
G�DV?P�PtDR����o[���������̐���7��1�$P�Vj�qX@9��~�6��V��J#����H�9=�D釘�ԇS��"U`�!;6���|NF,
CG5N���Q�[`����p�����m�ʎw*�@+; �k>�ʤw���s��]-��n,��z��&7�psʇ>���я|�<��cvgی��;ٷ�� �����i���)�c�G���<�L�q���;�G?���w~��e��sʎ�{�����;�M2F��Q�q��e�e��ko��������}�<���{?�h��˭����Q�;�,7��^ziٲ}G��O��}���Kʾ����	�y�_Pn�����|�/�^�_���E�J�.?���-��	�����%��G��U3�7Lx���rྦ�7 ����1�l�fٱq� +ɝ�^��,`˛:EA�w�P��]��p�}�㤌�ĸ�v����H3͈�I�M����0�/�GR7ܢ��vgS���(���W&�u��u0���_,�)͚�����ua[����e��eY 觽qU#�BW�\��K���V�[�r�����/�V�<�Ǯ"�Z]IfM{8�Rm��˰� Iz���wo7���Ƕ�TUP�x�S�N�W2.��B1 �0�[�����~1�7��5[#�h�����y��i�f7�@����r�7y��lH:N"|0?��I�*ҥ`x�p��4Ә���I&O��X�?u�'x|���V�ФQ"�D'�EAak�
����AH������k�y$���S�I�+��YEc�E7��	�t��!�ӯ�3�S̃`4�8_�:&���h_���[3�  T@�����$\k��޾�7pB��( �r�4e�e�Lu"�h7)��!���V�:m�wZ&jrJ�](�ȇO�8��0`�&N���ef՟s�L���:kV��K���^>��ϖ?��?,���/�����}����~�|��~�|��-���������	���Q6{h$�n���
��ZE�l�F���8��/�������o����<�؇�]Z��?T�o�X�.[^�Y����3�RLFM_FL_FO�"�Z��S6��]Vl�X�mZ_Vo�Z6��U��_�;RF�'g͙k��ʅW��}�C�Z�vy�ͷʖ��|���V��/���w���P�I}$���$],�.��tD8M�2[7Ћ_�k78r�~���*cK}�B�|14 31w8��ӕ�3�# �7n�J�KY�^�8tf Kre;����0�q���ae�����2nBZM'a:����r���~�]ZO�|�m��{�/f
���e�ǢJ,@�-Sٿ���}l2�~����à��h�hӂ>h�����;��7�͇l��X�č��'�5v�dQ���W�0�4��n��RMA�ט�AN��A`;`��'�g�fN`��4h$(C(lE�(r�{�~����~��69ñR�?窼/͞C�O=�T���~f����YY��y���/JyF�"?��BC�i�t#
P�0f���x��G^�ЊB(���9J����㆝���ЛnC� m�����8/+r�������՟p՞�m��,|Sq��'�<�n��/����}�H��O�:>�rܙY�?̔�O�bRVV��i��
�=;���L��`�KDu���b߆����3�j�l�ꞈ���<YJ.;.Ӧ��x����:>h ��D����;Ga�a�hݺ��^!_�E&	�q�^�v�m�t�,���r��W�k��\��\u��,(.�nG��;q(��X	�<e��$��r����M=���f?/=�|�m��{�/7�vg��E>�e��u���,�4���	�Գg��3���cF�mG���;6�7׮(��ZZ^Y����|qyE���%�u�+��ו�������{���*.��P_�n�Ʋn��m�β���	�ŵ�R�Q�y�B)Ȟ�J���|v�I��T'���S	y�����:2���}���?�ˁ[uO;f*��Gb�"!�K�p�UN�q8���(ܩ����6=�d1ŝ�G�Q~�j�a��~t�|n�~��}[~�σ`0�j�=�k���"^�����A?�a��ǔ��0A��E�H�>9hK�r,���~5^����
߅[��%��>:��� �K>F�����5X��w�[��`�0 ��w�9���ܩ����~����/��c��3�ca1�l��4G�mfM9�3������)0!�����%T��WV&�QXM"]� ��㏗����/��/m���(K/���A���ʼ���,Z���7��4�
��yE{�E Lx��RN����J9g�#/���#��o�Q�0,����v��ڧ���Yz���f�[�ƫv-˘�tE��+�2Q�PL��AF�Z�7 �<�*灂�+������<@6�t��@��L��nm��*}��I4��%�"᠙�PY�%|�K"+����Z��U�오�l1IC������&� !b��B�:=0j�G;Jn��c���"�!�
ί��䎯�e���|��B�g���=q(���@�z#��h�9�S���r��Ż)�4�Ǫ��jBcd7�/�I9�_���ᅣ�n����sꋺ��[$/�#me�Jr�0�)�!�5���|-��7�R&L�V9^���]6l���̜Qn���r��7��^V&̙Qv�<T�޴�<��k��/��<�����K�(�-y�<�����/�'^z������S��P^_���8��L8kz��څ�<Zf͟W�=T�l�T�o�R���U�H�ݵo���RΚ=��z��{��$�~�c5܍z��M �We����������]$��!�g"�y6�j��U���S	��;H>ORN�+HVt1wډ��%��r,?�HY�U�D{g9���l��㸴o?��r���ք���e?$�	���Z0C�{�:#P֞4vH��H|�����;��!����M����,"���j����Ow[�AGo烈S�/ҎĉJ|z�g�*U�ų�[u����y�M!<�]��6W�q$.�r��)S&�+,(��{�oB��nb׌t�>']�#���9�\$���i|ճ�i�kX��I��Ta@ˤ����	��Q�E��rЧ����|'�ۺu�?��U����m���GJ.Y���'Q�I�`F!��AK-���q�)�|H�����_��������ݿ[~��r����6Q4s���o������;�
���G!;�T�p"�H�J�_uqڰ�yi�h'+xM���L�I186B��p����G�U"�P����t��&WǪ��I�/7V���)�K�]&��&i23u�2e��2�Ɉ l��Xb�ס:��?
P��.�$\�ʛݖIϠ����2!��-������Y_���w���YW�?��.rm���\i" �<�[����=��$�N�����%����pD2�m�n��^�,�#�n�W����_��k_b0C8� x�����&��nlP��$|�I�J��_��W[��9�x[uȚ��j&��g G����r*W�qD����\6���#X��Pa��+��C�9:u��zG���.���\�EnLঊ��Y�g�>[�f�9���_&q4몫˃�<Rn���2KJ/���{���9/���K�\P\���}ѹe��SʎQ���=[�;[ו�{��G��㏕m㏖���}S�7NQ��9^��<R�;X��S���X^Z����fIY�{s)3Ɨi�-cϚZ6��^^_����xQY�jy�,�: >��� 3g�\_�~��וɚ��\RUV�u�v��7��A�S�Z�h�M)���ԃ)o`�I����a�|ǒl�<y;V�H!�#vźn-��i��s�PU�dx�,6Whr�
��p�F�}E��hw��W��Sz�HZ��l^:-<�,o�����Go��E��ϡ<4�95����Y�nA�[�z�I0F}���QWc!����ȃ�c��o���tZa @/ ��9:B���UdW�g@��������"��o82�G�k1�%��Ǩ�f�\�liٸa���q��;o�d��r���}N`�E���K�7\��;�SO=Y��ce����G�\��hDh�st$LZ^���d�2�8p��DF�t�0�F�� *�<���3^L:��C��K Y�U��K�9 F�K }|AHJ��(h,Q����B���2���b6_L�^�뮽�\r�eeƌYV����E��-A��&^*���(�ȫ
o���F	P9��Jv�����3o	/p^Bx�d ��B ״1Sڽg��8�֞Y�n=@���w�`c�I��ZA�&��9Q=7�f��]�ZHh�H�ك8�<s�w�Q��|�/�1V�d��PY�D!�n�-C&_�j
+����2�謲N@�<�����U=�A�޾m����\w�P� �M��(��4xw�M�cHAQ�jhK�)��~�g��KFx3�6�j6�ˡ�'Y�C�k�jj��t��7@:����9 ���X�@Μ�⛯*�8Qh�N���3�|VY��?�ʊB�,ȖZbW��Kק���e�r3a<,�N�2�`�军o)���c*;���o�T���.ER:�9�˘�˦C�����W�%����F
��#�1)�{�+���&X�G	G�Cc�R��)�*��ƃ�˲���k����Y�}獲v����*��d_�y}Y�veY�~MY�eS�)Z��1��1q��k�TΙ^-%I�Ege��� #gF�e~���OV�̈́�� �72X���$��!@Qp':�&}[�,�H���r�ϴ�O@�!�d��<V
)K�C�	���r���G�Ӎ�w��0�k�(�����V:+?��?M��"��2�&��Vp�q� [LG<��~����J-�<2?��nLM`�� ��Ǉ����:�h��O~-�~-Qm��+��8�U���e��VÂN�a1#]/�H�x��7�o�Q6lX_�L���2k�LR���C?��&�Og�;�駟�;Z��@�
n�ի�؂�	D�w����%���aB
 � 4lb��U�ݫ����ni←H(�A�́9��,X�#H-����1�"�f[A����(>a��]V߸{tÆR�{E�8l�g�d��k�a�g�� ��i��=�#F��
ʮa%�� �FE�ʁ��ǭ��̾�J����g�P�@>��D$�+	5^������l%ۤ��4���t��ZO�<���Ѯ�(�g�	A��r�l� Q����Is�.)�(�|X~���V|��\�%��R%��7>J�tpۡ4xK7V���M�8��]�7�pV�~�򶠴T��t�kڠ��j���n\�,��4x��Xfd�#��Xk�A[@���0	��_�1������5k��m;,{e��~�=1�3�s���o�d�x�v�-/��AH����T��Ljv�`W݆��5Y�E��N�3�\r��傋..�$7ė�{w��۶�%kV�՛7HQ�>���w����>�����W��뗕mG��=���}����c4!;�?�b��lJ���y�l9��,޼�<�����g��Y��4!;v��:~�l>���ܲ�,Z��,^���ݤ>��?�y/��
_�x�7�j2>f��}�;��������g��Yr2���q�t��v
{��cBX�-����B޳]0(��J�L��<yџ_?v��.����u�3? ��b@�'��D�過S�C=��*!�E�G�Dl���CaV{B�/��j?��p@�ޅ~�|�l����h���a:��7u�Z��p�S���/5�]�Xl�<�?���>�h�[>�v�Yt�[�Ց��4�j�bb��ңO�^H$�7q����;�����a�e�|��I, ݂~��>�w�~��_��^��}v�A�yڈ.���4�P�����͔������?Ww��u��p�0$GJj��Pм�RW������-e(i����[=���?�����������˿�w������_|�۷����������O�����/�<��c�C9h�	�s�@���64��ɲ5e�i�S�u��>��ܪ�
J(J/8
���
�<�JP+I'ጵ�Y�D�CI@X���v���4��P
�}�XS�gY#)(�(f�Knh�q���D��5+r��j ~(�|`�Ƹ~���z��A���וu��zaX�
-_��,Y�T3��eq��^���N�Ld��H8��"=)�aB�z�h�<��� ���9]��A��#��&w��`C]Ã�%����wx�����=�u��� ҄�:2�G/�0y���?�Ay���ʪ��4Ѣ�<$:�}���7�7�z�<���3�>S֬^�t�&�� �U�b��v�N��E�LH<Q������u�&O._vY���{�9�Ϸ��Gq�n\_�Y����䭲hՒ�l뺲f����7�/?z���������n��=k��c��c��R)�>�<F��<'�w��񒉩�˘Y�ˈi�щ��)ǻ�A+�[�-{��AV�ǎ*��*o,}�<��K��7_-�6�-{Uα�֯\���{�}�{�-sf��3�!#����ʺ�p����@���~���tl��	�`�nh��2�Hd�n�D�j�a@]�m�^�H��e��N'�����xζ���L���"p�q��0��v �ٝ�j&��/q6>_��W�4ft��+d�t������ �n������3f����@F���'=��������1����m5`�>"J#�]e0v�<�к�d������#c�A�&l-[�/@��|V����?���o�Ϳ)_�җ=�����`��q��_�J����ߖo~���Eo+.G�B���'�����G\t�~.x��u^�ܵk��ni+U���J���O��/��R����;���9�2i��-�j�+Gc��\w�u�j��!r�[�|%��87�w�n۾��X������+�������z!Xd�\b���apD��Kq۷���+��6�������St���t�`��|^�!MPw��-3�eeY�"�+&�Jg��{�qq\��g���('_m�\h(E�G8�5w��O�7o��"Θ_��Ż9���%����[�:k��.��_��|�kip�Qip��
�ie6&��T�\c�r�bL]!|Q�0z��V��y{�H<�-#���y�}͵�.�F�V��'����S׼Xy���.�̲�}��'GYxq
��+r��B�������r����ϛ7W��3��� Ǝ�	��2���J�d������1��4� ��ƕy�$2��p�x�eŊ�e��v� wLϝw�WQ�y&t��v�ד��.oGq=��O=)���+�S�I��`x���]��q�A�6m�TV�^�> ~ [�eׅ��Z�liy�����P6n�X�n�Z�j�B�K��ר[䂉�A�[З\�R��σF2ŝ�������e�UW�����J���e��e����4iyH
顲vߖ������&�4y�0��b�q�c�I�WF���M<-�I�:kYx���H)f#4Q�D���|�_�_}nMbe� G9P�4qAn��"�$��f���gN�o�v�G��<��n}��ݠ�Zw�f��W}/B�w@W�D}���jX�9��� ���tȁ��m|!��{������CNg��1�����g�R?͗��GyB��UN��,Ca�߉�^N��	�����v��.]��8�4����H�E����_B�f^�`�0+��9xv?���υ3	�ˏ���?&Y�v��3�9|�N�/T�h��G�w�к�Bv�n��E�_;u�/�w��-�E>5&�BS��6a�N���ݜ�U���(L�1�O*�x�q=v�^�f��Jګ��8��zn���#l�w�O��ȯ�]�v<����q!�8�7���8nz�;����1�����Q�k��m�Fܽ{�����;���!G,�%�R��j�X��r��	�&и�N�GAN��W�z�M7i��ԟ�nkh �8&� �ab��~ao@���RU��*%�WV C���A Ӥl^eR��H:�'�>R +��s��,fK!d���%��0��R)�^e�N�+P�A��*���S��9Z�9�Uh�t��xJ7�eƃK�4�4�g\ۄ2�闩#g��FY,��$�\p.� 5�b B�{��4�y~qg�gi�:[6*h������LT8�4��� �>�_�)i�f,� �Qz�NG�%��䒋�u�]W^uU�������Z��ZM�P��Pb�yB��{~Ut��*��jp+�\�g��Ԥ�|b�4>�+�oD*&�����mxf��i����%��K�F�M����EǑ?a�>�aV^�<��� tz�t���8wZ;���������k��.|���ƛ1Q^�T�����%�/z���¼��K�g?�Y��Oj���2I�����2r�I�0Md���b�����<�����mw��c#4�qFw��uRvW���V���ה-w���w��{7���[��=Z
��c�����H�{�x �f�;��Ǫݎ�/�&H'�+�'�+G���{�-���M(����<V����]a��]�JY�ycy�{��y��ݸ���ю/����s�s[e���n���v뺷�~����&7�U�1߁!I�2�t��ִ��r&������x���S5����z�_7����N�Z:��0]W��p�8� �do��`�ƪ���;*���]�/�q<k�&|,f�,A]�H��D�Rpe��B�w�cF22���!m�#hE�t�Q��^�1����T{��"�~$�B.���?��p��L�Ʊ�P�CQV_E��m���f���g��ue4͕���׉q�~�^Q��G.�x�Q��z�0��r@�����W7�|s���>Z}�_+I�m�������?����1��o�av����0,(F���P�T3�z&�\���ʔB���x�&L#E+�*�w4b ��l�3�RX��ѣ���0�8���5>o7jV����s�#�9���%�k���|�,�Ї��"�������'������O�?����|��X��~�H�bݤ�"eV>�h����k���W��M�d2]`�W��`��y ����L�2���5kV��{���G?,?��O�O<^~��_��Ȏ[��w���|��P�N�N���K�XR��eu/:�q�4��;��8�0� ��K�`�Y{Ъ�u(5\O�{ ��Ǎ���IB(?���2Yce�/��+���_���*_���7�����|��_��˗�����/|!��_,_��˗��_�˿,_���������Oz{��䗎"��0��d9��l�c���C���x`��ީ�*m�̪=Ϙ>m�ߪQy(B��'�A�֒[8�t�D�	G�JZ|.x�8^E�s �����˖�����/���U�Vk��K��ޑB^�j����Jg�ick�A[T�8^��Q�� �U�&r��2M�F*_QF���{�E�<u��X)M{�/�P.Z���\��l޽��:��l?���jz`��o��r|���IJw4�gE��L��dڔ���g�yg�.����Y��.3��M-Ea<)aES��*��c��������(I	.�_�<,D9޴uKY�xqy{���5��%;��;��=�7TP�|@�Q��<k���#ŕ�GȬ�����@�]�!�1(ۯ�_�\��/�T��v_�� +�T|4NYĂD"4u��.�u�ֵ�֏g ����Ҏ��cB+��W�}�6���!�m����Ĥp�ڃ��}-�.,��{�����g�=�'�E=�H%��R���
o�!����� �D�<)K]��8��/随��2T�)�o��[*��x�Q~�|����^�{�&��&g"�zWR#X��=����[�.s�#�,a����zV��.�=#���Gy)��*�U&n#�F��#5拦�*d^�^�v���A;�s�̎]c�9�6Rv��؁�L����{x��b&GX�@ވg^��oXpeV�$��y8@�e��ي�SeI��}xQg�^^����6ڻ{wyE����o|]�ŷ�+���3w0y���e劕>����I��C>�OL�$���.F@#eAa�������YF��RyY����.�b�j�j��5M��]�t�5�����ʖW��a��.��%�g�c�	�֝�^��!XW,��V|��-�m~��(�s�����>!��o��vgw+�Y{.�c��A]l� d*vL�d0���d^�dۨ-�j��q��
d)G��A����o�L&7n���ʜG^����=�m[��~�Ŷ�>��*%�M��.��Y1�*Ϻ�G9��mYO��!��_�FlOqn��`u0ہW(�$�R _8㎼�Ѧ�����u��W�@�B��y@����':�n�Zv�/���Β����+Ֆ�/���8�_Y%f���)|�I#��o�8�Ò��j7�����{l���K�M��Tλ`�FVI�l�ZV�_S���^����㜵�|�&�c4Qù\�p�pr� �RJy-�8�4c�2k��r֔i��e��ie�������ӧK��Q�̘�/��Ѐ����bń-wJGy�J
0�?��r���8��D�ų��횔������'�,�4y������+��}��h+q�< ��[������f��i���;,;`/��.��1�|&Z����I��d"��2n�����Y�Q�A�E����C ��W�8%DY�'�Ͽ�煄����Y~���`|@֬8��"|�g�3~M?c�
���Aq��qz0LT��������u��_��U�b�û�
���r�r��0F��y x%�b���w���ib����/Ly�d���X�#���,����ښG99�0y¸�ɓ�v��@���{(�Ï�f ax��	����6���=	V+��0�����y���ڟ�\ ���4�c`c+��o���7������/IQبFrX�����k�����|/1H3��^�t�]��H��z��k���q�&�\x�Ő5���{�/����цX9Ma�l�4�e����|���H�� ,B`�C&3+g`��+b�!:�"L�F�B�L�L_]À�գ���-����ٚn���N��������Lz�@YR٥s��Tn�Jn���8h�(~�/GǏk�ZD~��� /t��yJ��g��O�K����0�Y�3�J��$d����M���Ag�3R<��`�&y�_a�S��	��:�=��}�y��+����n���r��W��������9iV'���j�+����ղsN���9�碣ސaJ��'8Bv"�؅��>W�p�gL/W^�зpQ^�ڤ	$G���Q=X��&j20it96���4�K�=fE�b�FJ�XL7�L/�w��2c|���<E�j��2ej�2mj��a�dV�YI!:UQp�
/J���Q}��O_&Θ�ൢ����W)w���9��^xQ�4Ex=7K��n-�Ԩ���n5�i�Dܶ�/10�Ay�m��|
Z.�����u�mM1��a�b�y@O�*�jh(x�L��U�|��Qw�fJN�|U����6]�x0�1��B��_���X�7<��Ƭ�4���zn�o\v[Z�[��������ݱ�X�Oh�/L���m=�B�ݺ������f2P�B�b�?��R�>��/�/�᭛����>2­�k"ې��S�u<�-�'Uv�W��N���\<h��"�<�߼i�����?��o;`�������/�s�	^�z�ͷ�m�ӟ������e�����n\_�|�����/�_��_��|��rڎ�;�|%����a�e����n��_gb5��P��� �Ǽ�Ɩ󫯾j���I�2����:9����`��t���hBzw1�pѹ�[��3��$�푆8�r�Y\��s��z�F1S=��v�/��И�EGf�y��)VQ�nᙣ(>"!�)!y�� ����jP�ܔ��y� /Q�*C�ŭ���8��u6�.|]l���!o4�.�?�.���������}��I>/	�� �+�'�<R
�#��tx7$l�9�͙���w��o�f�y�E�L��<OE�0�GF�lWغx�@� �����{ʧ>���G���g~�3峟�l���~�<��#���-��ˇ>����#�G}�|�ò?���������xS�M�27I��|�~��S��4�s��Fq�j��*p܄1RzG��Rg�?O
�5e�d`���VLv��)ewSٸiCٺc[���oQ5Y���qe�M����q���R�	�C�H�[F��#ǖ)cƗ)�Ɨi���P&�	�(�IjÓ9�%9-E�}���j��B%�ݪ�У��;j��2v����c<a[�|iY�f��8�,�?��ο��2g�\��G�>D@zTo��=7�1~�PESж�a���X�1��yV@�E yG���xƌm{��Aƒ�R�.&�n��Cu0�ϭ,8x��p����$���m�n�}cE�G�Q|b����L�@qq
ԑ�L�M#���2��� ����ӏ���YOk�0m�u0��S�	���,α�]H�|��ɿW�U�`@�~>0�c7��Lށ�,��8����`x�8aE:Y'���D_��;Z�Ky<���Fع�i�����2f�G��m�˾���I�VcX���`�c�0Q3 ��Ux������{氷UaX�ދ��rA�:p�[��Fk�/�ț��}�ۺtB(��e�|*glP@�$7�.�~Y,<=��<��lx*��E �$ؽ:�8���v33$w(��(;��	~Gԁ�Sޤ���9���Ӿd�vf�|<<�痻7`��5_�/AC^c?B.0�r!�Uc�n�%��zqh�<�,�4�9� V��4T>RA�G;: ��e�R
�h�KT�L��d��R�0�>����sD��-tn'�KV�@�A8A[?0e���"�WثKIEz�ӠϘ"��g���F�3��vܻ�� ��d�)m9�}�y�2��_wxI!;�w˱�}{�H�N� ��pl��
����GI8��䏻��|Ю��|��l��)a����g��*7��S�/��v|8ֲ���r�ǸFl��6Qr#Ew�_^@�rFY=^a���A�q��g5�2J�dW �ӻLИP���хќ?��!���!�(�<J�T8̽��Y'O�P�[!�w��5e��->s��w8?7A�0�M�x2mȺҞ��`A�H�h���[k��>@�� �NIx�#s�4��/���{�����Ƀ~�C�#^��B�.�����<&�"2r�ǻ@�u��A�����M��b'��}<�<M���S�����ņg
��|n���2M�5���YV�L�p��<!&��Wq��'�+� �󻃮��oF&�}~��UH��g�%���C��VfC~]r������Y]Z��V��L�$8�cg�K��=�ܶ}�������A
��#�L��Q�L]�ӈ]i���u��K�f�]��E�|��j����d�5�l&�pe`t���`����(O�8^
W]��3d^��9�`{���¢D�3� ��[�q��GᡣˈJV���8��j�����+m(�/���°�y�-��Q�^�zu���k˴iS}�N�{9k�I܃)W�0p0��zG�ɹeV�(;G,���f	�;i�Y���������p�8��v����[8�H�&N(��_\vy�b��2��_~YY�`��q^V1헗W\Q.��2�Hq���z^p��g��k������(��z�e�u/?�ҩ�\t�2ȳ)o�A6���lq�d�lY͔�e���"����k/���'7+\tх����#W�]|�%^�t/�8�^zi�7na�Y��Pq��������s��d��Ag�\�|0�@A�y5���B�B9����7��������?J��U��ry�C�yt���F�⫼���ϊ Ǌ~��_����z�C=7�a��n�� �Z?����䚶#*��ݷ�J��f�ڲn�:w�[�n�≝cH|X���X��cI(|���:�oQ��փ�0�s������b!����«��L`�������e���e�~ɴ��C��M�@>u|1al9���Q߸�B9/�1[|t�R؏Ӈb��(V���A��x��|�(
+\\)v���r �D��h�B��5yQ��s��W����e�����ٶ�a�Bn��5n7?pF{��հ�O?�$'�2p��8�wo �^o;{����1�5�(���v)�	=�H��'̐u�/\"�S�?�:����ת?ާgv�N�P.8��r�}���%G�/�������n�j��iȒ�r9f�gS�D��&�ܡs�n�%�H܌�g�1�ex�@�p3	�1�q�������+F���鏴��ǈtx�U�d�k�d}��e��%27�or�ָD��'^E���qIiP��G�Y�՘2�`���1���������e$�u���Y�:�߫��w��^A8o��lB���Ј��rG�6�Ǌ��n�,���_�'7�E�S^��s�������_䃃�)F}�c�]�w*���*#�L���iwBa�;|r~С��+r���\��`q̔��Lಯ'n����:/�ċ���rҧB+7]}�U���5ҩ^R?����i�	`�>�B����x0&�\My��|��lg��&�g�Q�βbŪ��o�����P)(n@4��8+Ql���Q~,�*<�P��Do����t��7���B:|�s�cǎ�B�����O��h`#�B�����͠ �� E������~���U���C_���<XRQ�^���ݲS<x�_�g�}�|�ӟ�*�_��_j�]e�f`��9s��b2�UM�4E�ֺ�
A��=���
�%.�-����|r(is��)��ӦM�pOQG/(��ڞ=�\.ңC\ %�	�huH�ݲ.����Ł<������y(�b��V2�/҇�Ç50W�rr?*��#;L(
Ń�y��p�ޅ~Z����8��A7_�z��G��^�������A_?۷o�W�K��Qt8�B�	���4����L��M�L�Հ�q�h��ՒҴ���<��#W��6k��]e��ݒ[nh�͙9�xJ e8Jt��s�7�ආ�M�{g���ǟ(?��ϭܢ\�r��}Y�<�N�P��տ�W>����(g������4;r�[�Ͱ
Z?:���B�,1�`b@_CCqL�aPÝ�'�K���Gʀe�����Ea{��'VH��C"���(=�P�����A�m;U7+�L�;�.�o�W�MU�LUO_FΜ䳲Ǥ�)�PD��vP�4�i�cF�)��M,3�L+S�ޏ�Zm���3qu�΃���{��k/_{�U���UF�i�2��q�x�G��]q6�(3G�/c+�V�-cTe�^t�?*q��z欙j|�cc���^~��_�-�6�"�!��3�:p�_8�Y��Lj�Z�����Ν{��݅e�)jR�Yi��O�Ԅ��x� v�X�~�z��ePajӤ����h�Q��1�^xN�Ν�##��I3�]w�[~��]\y���_L�QH*M�b�h��w�?����9����p���L �?�h|�ž��3��V("Q�����{AI�19�����I4>O.�voS�oj��3�M�����"�6)y�'y��>�]�[��@�iEW~�'ͥ��~�K��������q0�F��G���,���݋�>�	�~B�sC �r?��I#�A�3�^ ��'�8(�	��S$�� �X�H�) %Z�q�;�+�am�(��.@?��{� ��u�ԧdHr�+��!k���<V(mv��3������	?ءd��w��� c$qh[�� &��v��ђꟴH���o��]�R_ʤ�����?�g+�����v�ck�-f>w��+�E���������#�<\.��ғ���l�@���o�J�c
� �`�gB¤�4�$dU��0%��?��C���x������2g���{�)�o���D�W7�h���X���p]F���A
w�����܅��z�����뮻փ����ʢ�޲�Ȋ���u��R޾d�:n��9sX�/�sq�~7����&�^Imĳ)G��-��ZqmE�
fǔ��Q�p�;G2�1 ~Ѡ��ի�‾���Ꮅ*���Q���4Ff�ؽ#�#��+��C��Ӓ�"���qQv��(2�d�z�:����6'B��7�x3f�X�`�.;Qh��L�I�֍�u�1��
�3g�PG=Ɠ2^fDYY7NN�����E�Ը���N�y�S;%�,`��z��Gg��.��|�$Vw=���7��` �\f��[^�u>��kزekY�rUY!�:XEa��Hfk��E��0ݜ��s�f�_��iO>������ 0��j��1�@� �$J�:�e�Wp�j�Q�ؖ�[����v�@��޽|5M
��2>�E����`k���J(��[o��\s��eޜ�^գ\�zMY�xQ��͘q�_;�(��ɋ�(��d�������W�H�U��^�](Ӽ�Ɨ�Pl����� ��1)�|u�z�	��HkV��=��U��t��wt��2Ay������M��+�>�U�"1q@n�����m�̧�Ozap=�/u:,��ß�7d�W8�OÊ�Ꜿ���H1�q��2�o�g��P�$h#�r�B&>����� �f&V\sǮ����YD@�X�/ҋ4èiV$��5�����~H�.&���?Xp�i��G��|�M�HS�]����)G|��j[��x���R�X���c���-�U���2B?%�Y���cslA��q)��W����v�;���qL���}�� ݜ����1��%�Z��q��1և�V�Z�xbb4R�)S��ϣ�����]��[��b�<+�Vhk=zd�s[6��r���Ue�C�A�Z�#� (@׿$I^����#Ә�Α:�V~kx[�c!��̘�t�v�h������D�J�5I�T�,�E?r��H�	���5��.��b��Ցܬ���wB�K}\�
�-����{�7m]t�E��i����@�}�F�Sx`�je�<PP���×�3&�$�=_����HfH��j%a�e>+GX��fJXYY:�Y���>�6��̿��2$�*�p�3~+ZJ ��l̓4�+V��e˖:������캱w �Γ/�� R��Rͪg=�'�� Ғ�4�|H3y��)�e��&:�~e7:yVQ��6n���0V�f{UY�j�;��*+�˛gʿd�+D\���ry��48ˆ"M�D��JA����UJ
��93u�m.	�����uc��Ѱَ�<2�)�Y���Q�F�tT
��
�Y�ee��5d��nm~2x�M��\׋���r��^�a���9Ιs�,*w&pl��Hǂ�`zu�v�'�>V��>lJ��X��L:l:�����RI����4�6��d鄬��{���yi3�]�+Ux�%�du���vL_?�d�_� �C����)�����z�-Юx�V��2^��J�w�L�R�Ew8jQP9V0a�D��@�.4sN�6�L�����@��;^�)��Z��-��]�퓎�Nv�X��h=��.�;h�q�W�ډ_�
�� ���8�ff�B=�\b�h���Qv�������:r\ʮ�M|b��ڐ	䟉3���x��M�L
NE���u�-j���o!BPgy�e�� &��;�0�TTB'����I�&�P��[�<&����@��$�Т�Ι=�\p��~嗱�eo���v��	%�V��u��u���b��$ɏ�P��m�	 /Us-_*�(RC��`Y�bu���/M�~>�J!d��+�|���+��CƘK#n�<�#�C���@�h��\1h��@Pָ�J�qW ��ca���+�<����>����9Ɓ.*��3c��}f�3�[1�&m:ڸ&�bA#5xn�z���s�q����/@*t� �ڣ�}�q�-�?ڂ�X�� ��w"~Ј�y"���]Q�(�p�#$\G��^M�&��!��CS����d9�ϡ��F-䗲6�#:rm�x	����i�
�'�.���iSO�����A�@q�-+�H��*�JH�B�)s ٺ�#��3��=�X��;�ӿ������`d&+=W����������/������Ҁ�@G���L��˓!�dM��� >	�H�׿~�����^�'<+��Yd5��� o��Cٝ��xӊRne%8���= I�V.@��)��?X5��.ʮ�өd'XUH�!�(��3�v�%�Kn�x뭷�[��o�!|�����׽M���r�3
�+���p|���x	�R,&N�ԓ7�s�᭏�Xa�~OV�B&� 4�.��O�mK���	�+��Q�V���ȳ��ͪ��y[<{��j�_���'�OZ�%����_*���Jy��W���W���/��w�~��2wCt��K��L���CٍΏ?�F��>�c� ]d���$��&&�J-g[Qn�8�PtY�E1 �;:(�]�E�{WvcP	{B��]�1е�Kxt e�ɗ�#�'V-���(}�M�s����f�� �h�'�u��(�8����P�C�J^8�5��r�=w{u���D��Z��T����*��x)$��J�����[#��]�S&
.o���\���Q�A��#��������eQ?w�:���r�pI;rYU.�pT=EyHeޯ���/%�(�#�+�5�aE��p��W�F�&x��ˤ�	��m�I`�GE��lǍr���И܇Wv]�u��`�X�O���b�3ݠ�1��c���i_r�v/i����5�l��p����#?��YF����¤��ti�H��ejw�����|B���rL��|��a�!�H�<R �9��'L�<�@���~�i���;���ر�lݶE��&+a�=���$�XQt )�Ȼ�6�< Ƀ����o�y���\�3���`�
"��CC�e�a���b,f|"�DL�H;5�X�@
3����\E�n���I*�<�w��)o)��.��}F+�y7���=ֿx�6_0�E�P�Q|3�P\��q��0�{L�<N%7u��hCчP���G����О	��USM�����[�9��u&�l�̱Xn�Z�>��~�
HB�T Z�ly(����sU%��))���1ȣ�A4��0%31����;��H��]rI���;ʇ>�!��-��?*@�ef�4�܀�a�&iP^ٹs�;fV�b�45�οa ?ҡ�A�(�6��������V1��cD ؚ��(�[�ni��� �S&O�
+�;�T0#b��<���"������3x�iC/o�/�j�gp$g�C) �/�	��Qxi,�(R���P3��
%�I�(�Po����
�j �@g;N�9[J�ԩqnز �^Vu����@��;���L��+\��d�ȗ&��w�ꅕ]��f��倾#��N���b�$�(}�6n�
7n4�Ό�qL ;���(�1Z��Ʊ�T4�.x�nwe�����F�5�XEz��R˱�io(��X ��ʯ�|�R�K(�(�����w��8RD|����OYq����FdO��\�{9�G��>�P'3g����\{������e����=0a�wāOăg^ِ�g rL/*Wŝs޹Rv���u�π�J�Z�diٮ>hەƕ���H�=6A�x)mue�9��]=�J�ꎮ/Q0!VG������N����6r�X���}��8.y��Hr���2E��Pv�#{��	#F�%������\����\�IC��ǭ �k�oU�5-	Q�v��m���'Rv��͵c�e�$@�L��������; 9�0�q��
vchS(#�첓�lq�̥�^fe�IF$FS�.I�,o���]F�u���~�D�m�*��`Ļ!{ԏ�/��u�S�]� Vx�R�h�Or(��Ue*</RA2i�R��޽C}�N��4u�I��	>C}2.��IY]��&:[a*�����<7���HO
�/�����`WH�?�%|C��z�M��w��	��W���=b\h��9xCޑ���7x"�͍+��[�ƶ���s`(�(�3�s���4HE7WY	������Uчc��}�J���G���-�ڴI׃�<>Aqx: V�KX����?�>*�˟�d~�#� �b��b��T� ˤ�2IC~)�9^	OI��WXg DNN�Iqt��0+�_�wu�W�s�*�*!;��|N�f_;#�ѡ�s�=�Cx��q��l�(T23.^tzY
&nx�'˓O>Y�}�Y+��]a�T�P��y�UW��}H�J�A|<geb�dX0��&�ۢT��o���r����{�}���D�ԧ?U>��ϖ?��?�Y�r���Y25]7&fg�4�m�C��
7����T�?:'ν�L;u�����A��	��1�X�D;e�:mZ�<O�&e�,���}��gϞ[f�#�N:�8��;:��1
h���NA�G��1 ��@r]���+g�74������ƃF�N�s��a�KL�4;o)���^���1��Gt��|t�pPθ�{{I3yB���A���,í�Ti��m��H��c��c�l;&�egРsC�v�s� ���tU�������~ut��B3/�:�ikf&�Ed��-p0PWAc�A_�نf�e��7�k��R^|���s��������\��B�����f^���`�ωv�e���g�P��p�Y��G���.���y�,�3;F�ner/ד�щ�B�c�5(�ЀXT_�5�9*S٩^��:u��f�r���?#��"3�
t~*P�c�"<�A�`
0 s��<Mx��vڭixA���պ9sp��JؼdQ�:��.��3J����l�L48�
�ɯ�=��?� g��T�����[����V�nxξ�v�X5��Ph#,�"uG�����8�fz���Q>�Ε@C�cue�6�d�?���؅�&�� F�A�An�y0��tIq���x����d9Y��/�.�_��E���D��G=���/��j{���(Ҽ�I�<�wxH=��U�������X��|"��e�䇎Riֳ�D��;�΅(�\���]��`r[H��z��:���&ԛLҌ|ɄJW����EV�YQ��g�n+�(��d�W5���]8���: J��)m�w�8�z����s�Ϛ�0�U&n�lbYx�U���p�[��>��h��;a�y'H�����^Ю�_xtݵ��j ?���Z8+�,÷��"ӆ �e#f@E9c g�;��d���;ʜ�g)��¸���l�g���`�z�*g%�ϴ2;a�䋉��}��Z�Ty��V-d%- �2�@��|ݍ������{��/m\x�E~i������]qŕVbt��H~$m(4�a;k�,�Gx�yQ�0߂(A1�Up��S�5A-J�7�h����UCٹ t��mʷ}�v�5�{�VΦY���";�/f�w�ye�y�}-H"��s�y��1cf9o�|��2k�6΀2�G�u����{ȟ��C�t�>*�e�������%�ߔ�ڻH"�oA$4�i3XU�i���FQSpI��ml���[I�1νƋ�����3�g�gϞ�I����Η�x��k�1VP�X$Ag�4�P�9����>��0te������&��*+��%�*��Y�f���E���W�!&�c`7��g~�z����Rt�tbC�AеW�q�_;�_��> )u L���>}/�����^�Uǖ,�N$�������t����(W\��\r�%�oP�X���{��5ѩ�)uҘr|�~Vv�O�F)-�`4�-�n݌�#oLJ8 ⱋN��1
S��>Fu��r\��R0Ty���1��lD۬�JQ޳��gew�&�hJ19���~���$��{��(}�!M(#����Ir�1o��:L p?��Wv5q����)��R�C�� �%���3�(�2�"xg��G�#�����d�ˣ��QVgLW��>�+�OS6���)rj���8_=��
k���/�&�Ы�2�m��d�r�**2�_>|�b�J��&�CX�L�*F��4S'�ݘ���mE퍾:�۷�ݱ۷�gvio(Z���,*l�)��O�Zy�	oU�EJ��9�[��?��"yuަ�r�=X�U��j$����M�Z'z���G?W[��-L���ȿ�g��޸U^���tl*'�r`~f|�T^(�� S�*m_��oa���@i�4��������a�3�F&h,���N�-��b`�׌�o.������?�$�
2z��t������g}��������1�c��'��3�s���g�	���U���/}�1�$��:5��e��5�Q9�Sa@�䝄 ID(g��;΃�>T�;���o?[���4�r��~��f��ls�-o<sr��~b�Wȉ�`P_�|����@/ɫ�	B�2&(�z�L�3���>�Q�֘�l�e�̘ȇ*�JX��m��i%@
��c�Q��(��2�"(+� �g�C`YmD�奺\�����DaC���"�h�q��y]y����5D�]{�ߖ�"[��&
^�����O���~n�`�>�4���@= �0�(�`W�̋���QL����D����!ǩ�B�P��$�UW�6&?��x�����?L�n��&���r��_w�F���t��?�<g�!_�����=�И�n?߆aQ$�?Պh�~�K�+�,)�H7lԀuȝ0���ڄ.L���4ߠ��V�5U.W�"���[�n����{�N�����d���P��K�^j�n�z�Gёg}���3w�M�?����bMx/��/̢D���D�s�os����ء���&+�����W�̲��k��z�;c��rn�8�E�A~�ᯁ���������G�������륜�Z�J�yPe�'ew׾2N��$�ቓ�>�G>��JJ<2y�d�}���z!h�<Ci��� P����p�O]�w�^Cީ�J���&���`��b��� �(/�+Xr�7{�����?��B6z�O��9g��r(����"����XI�	 ���s��_�UK������Jό%(����N��(�vЭ�=�����.G�V�^��i���Th+\��X�}
`���FH?C�S��¢���.p���ւNė����J�V��Ro�OLK�ӡ����6 ��z`L��(��uaz*}i���׆�o�z�u�C�',�L��[�`I[� ��<۲���<����~W�Ȓq
9gg��<��7&8�\Eey��G}�߅�賹q�_�����<n���׽2F�>z �e��6t c�SCy��#��n�_�������R1Db.PE�fm7�������d#�Yj��72�UJ#��OV�~�i���`4�\e`׭]W^~����~U�z�M����CQ|^O�J�Q�A������}�Y�1���~����|�+�G��������_�k���X~����+�(�è�j44���}� �����N;��m"��ٌ��4w�
G���J,�=�3�mv�����E�ȏ4�731�g��t�!/(�FhK���%ϐ���{	'H/�h�j	T����2r���`����0A
�z_��;x��׹��)�[n���(?&�	D�$]�p���H�Y�4%,��0	�t�¹��ͤ#X��s�N�7��0ٜ8��v��0ڕ��6!d���nKd"M\���1��
�N�>K�,��uL��FFa���?�S�n4KB�X(<q���W����li���f"����B�H����#���~T�����N��������r$L��tT~A��2���64�+1d�`a{5xN<��!N��b+���2!'��Jf��eb(���ی�a�TZ�?�t�u�0�:[ ��0!�/�z����;K
��Qc�K/�\^�u������M�k���^VMd"���=�-Y��&:~�Dj���s�Ѓ���~)�������Ǿ�-�-t�%�4�Ş>ċ��Y-f|���L���Ũ�Dܪ��ƞ@5�~�	�@�����g��������ػ��� ��/�a��?e�;�-�
�cȺ��D:�:�ߨ���C�UAF��c�W��X(b���+�K/�_.��E�K=��g<�Wg<���q�)&;�q�6r駻���z��p�4	��v�Dxv(�g*ǝ)_Uv�XYR��&Иi��>��,f��g��ʛ��x���_�\������2ifcw�W�jl�(�+�S�:��˖�+��\�x�	_�ι�'�x���*�=���&MW��>�|q�b<k��
�,vI�۴��þӁnG��3�BS���ee�tb�Q��
�Dx�
�l��U	x�`�8��J�-�	F�gY�+��c8� ���C$!���,��:Fɇ����c�7�U��m��3HL�زar��������h+Y�p�F���'HY�c;������e�� ��KmeDѥ>��3����s�=Ӷ����9���[&��)$ϓ��sb��B:(kO�J�J��9����9E�e׉#n��U�<e+ d,�f��@X��ӧ�,�Ϸ:���S��<7�N2�A'����TxE�a>!|���~��;,;g�VrI���yaV�
�
]�G�8�1AIR����}���c�H��`�+v��rT���P�$���f���d,���Qp͟Pv�9�O+w����fͧ^�d�g�_�]�t��եe�����o�S�x����+Rn_y��/���#�JE�|1�%)�\���/��|���cW����.s�x�
�e��6�|��Yų�n���N�*���8�$��3j7<�.A~=�r�O���[�V�h��6"#��pi��֖�߯'N�9����s�Ō��=]�c°i�<9��3��	�i�'ܢ��bDv��x����U����~���f���9ȇI�1�r��!t7��0��X��)l?玏��P���Ic�@��.��s���*��ʝ��-�/p%6/��((ޢt�h�	�	^"�۠���J/+_T
��A�2o���y=V�a:[]���n���l1�'�tb��ڻ�|%*��O	L!1��!,�U.>��׼�V��AQv:�.r^��`57?�eU7������p
Z�v�ؑC������ =�\�o�$��#�@�����=��[v���F�r�J�IÆ�9Q �	�K�f�
���3hJچ2�����`�zЏ��������h��A+�)�'���/���ɀ�UA�Q.z�������ݖ%�^5�7�9��u�V���i�!���V:�
��l����o �~v��"9Fu�-����LG,�g�V�lx��YC��FW��Pt�j��[�U�Me>\��Ԥ����(S�0�����üZ��9������M��N��0��A���� g������0f}aHC	��;d���@����U��=�a��i��G�$g��8�@^�!���|e�s���m�v�����^g��u�#7�0�5��^���)�?�����{��W��%m^��^�7p2#zrG�6�~��C�3�D�T�&��A�JG�f�jo��O~�Cf�yO�p�	d�'���+�uX�j���zb�I)�� �<��m�<F��՞�p��-H��.�T���+�(��C)�OC�l�V.e/@���@MP����>��U6�9���~�M~����򵿯~�k�}�+�����_��wҿ����o|��M��?������J0c.i�U~x�|BO�� N���`Vc+�ݶ?18�*+@���K�4�[A�R)����O~���������O���/�E��~�\q������¡�����J��'ȓ�A3��)<�">�QX8~�r�e���&�9�DV�x1�s��å��~��W$a������)K�8&�\y��C�ci�i���������1g���� o��	�p��zU�p3F�
��޽����*(s�ޡce���bl�>D0�p�?_�ڡ���e@;�^M��C%�2+��҂�$^Y�ߺ8��h���r��<��l�@��Q��Ñ��ؾ���8ct���<��9g�o��}���ۧL�X�%.��KT(cȚ_H��05�����sxuHf��F���I��&]�.�-�%&��U�^X��*�,c��*��3�����,s¨�^������}V�1��o� ��v��}�}|�o�K|}�S��;�ӟ�d���{�E��=�2y2�A�At6؁�Q�D[�����xs8V���pl��B��Ū��'���*�?��	 }���9-�ވ�٠�`Rh�x\�i�8���c�C��>������rԲ����PG��qCu��)�v]��E&2���b�_��;ec�p���)mb;[��k�=`�b�W��v�F��_МqR��O2�oӛo~�U�@����Go��T�1�H_�۫v�B�%�z�����}��֋�e<����7Ƀ&���6Cbcy��G���^f��'����O�̝�'���������Nx!v֬�f��!aX�!Ҡُ�Zj���!�H��@F+����2��2X��Qb��T1�������ڛ�D=!絢�d��r�\DҿD���^�����	��~7�	:"�(J����O��OQ�<�l����_e��O2h`Ke�ZaPFK�n��A�Ư�a��AoMIo�KcDL���Gh#�c��8�����/�_���?�a��w�[���o���'�?�i����W~�����G>B���؊1;~�Xm�ki3��j+���5,w��+v� a��Ã
���� C�uCS➍T�`�)��"�3��|��\O�����s�l���d4dn@�d�RPh����&��}`�.dƽY�Wjq��>�o��{�}���)��{�̻ˍR��47o�ʒʒ�55$/�G�EC�`����;���F��|%.��)Rnw@�CP��Π�W<�	��ٝ>�J7�-��Y1߸1�����v�me���Oˮ^�FJv��&M�{S�����p�� ��̦2~Rj�Y��!�;���u�ˢL ��0�GL�)OLv&x��6�m�V�ǼѸѼcu�U�Ӄg�.��~�����e�������wb�%8ُ��5p(Xѭm�-Q�c��a['�˕f����̬�F:��|^U��W~��Lh�k�3 ����Cv@��)M��NQvYͤ\��q"��x�������@��6�/��r�i_��y�n��顽3�ô��Qo(�����8>���:���/��1\%��9*Q=#^AϘ�* V�P�x�(h�	m���_G�W�p�ZeU"���n�W��1}u�G,8r��V̔�H��/���td�0(M�'�����L��[�<��y~;v�2-r�bJ9{�w��)4f7���.�'f?�\�<Z��i��|)��S�y"�go�7؀�$���Dl�nڰ�J/��L2��x �Eo�#�e��v���4��)7ڟ��ͻ~��`�Z^H��s�_�t�?v��D{�%3hpy��%�n�ц^����ʩrP���p+�:����w���q�LJ"��"r�֦��A��x�J�I~044�p~6F���k���U�� �`V����7�!ķɲ�e}�C�F�����Z�.��nٺ&HN��X���t�V�KeuG�C�	a�/� �$,m�#;�|����B?_��x>�6�0.򑮐�-�t_�tc�q��a�Ib�tԠ)�����M� L�s�й�g,_{�u劫������?�|`���{H9GE��ς���x���p04��w��I�ϝG�t �O%�X��r^��������?������a��g_ϟ+����rg�9��
@7�.�C(B8pa�-0���UP2�'���R�9�ҽ'�y����.��3��)+}(i�������~Y"qɒ�d�b�J�ИmX�fr�}��:�`
Jv�I+&ʑV<�\t�S���n�(Х��&D	`��2��s�믟y�/V��_�{�g�ӿ;w�>������
/��s��}���-%-�g�M��d�S��1����iX>��!�U��Ӕ�X�����/V�H��P1�ռ���I`���Z�!���3�	�ÍI��t��զYe��~��@=:h�l�ʓ2�Jg�G�ILg�{00��1)�
{X��R��(o�G)q����3��i�`��6����#$/��3��I3j���H2�tE�ό���S5A�Vg7��ђÙjǼ�@�x	)A��wS�'�|� b2���to����G_�%ZC^XIečcDL0��*)e�/�C���r��
��ŋ�)���#�t����E�W�xWı�K�l/��g��F�Ty��@M�Ӳh��S��4`���^}�7��p�ъ��%>e�M�?:�N���?b|�'N�Y��{G�R���5�!gZ����u%��o8U�:�I����e��N�����<��3����� *�?j-����{"�Ƀ��W�#��1z���z��I�W�3�+�b�����g,ġ��������'ܻ���O �L�u��H?�~��)8DR �����5q��)gr�Ί7�ݻ�ya��ɍ�A8���C�;����~!Jt1�]�l��7�Q��g��Kf ��ǯ4��tp|��w�N��9cŋk�X8d���B�GV���tq>��*vk�4�+hP6����	�I�1^SV�Y1��|����P\�p���E��P��<a�s��Ϫn�%��]~�qmM��4+�}u� �j{�@�V�2����D<�Δ�c�2xͫ��Q%ǻ��5|����3�1	�K^�)����$Ѿ�ƋX�ӆ_?�}�����y ���fW򅌆=&��[�)o��n����p~�<�*1�AI�S��|[�4&^+V,�r╂ի�+����h�N�$&ñ����sD��B��lis�BaUw�rt�>_�5Vn�����h3[d>kJ�o�\.�����7+���~D���#��?םɍ#
GF���wL�� v���:p��>r�̘<�̘:�L7��~Ӧ��$��Oو��!y��~��L43���"C�c9��`u�c8��Ij�=�t�:#����dH��>���^�_Ҥ��ĩ\\E����+婧�,�����SO=Y^x�y�o��˖x��/Z�Ѭ�X)�ݰkf�W�����<��r]��w#^~�%+�l3F���?�v���}��}�V�9��:�� ����m���Zn���	W�g��ʦ��=�]_���>Aʃs�� !�G�K���2bV��2vL��<�w�撚�D>���|7�GK�C&!�>T���i��2�џ��I;�O��#�xowR8T���ݦ�օ���!�<�d�T,����`PH
k&���n��d��:$A���2�X�ݾc�_�b%��y���	�/*�F�y^\�A�����m���ٸ�e���I��o��7m�m�.$A�	0���m�,^\�q�'��w�S����Sa	�կ�Le���pQ܈��vh�[�m+�*�����a*�C�m1ܠ=Wum���Ơ�+��h��P^�W�0���`f�����	|a�[fX��
��%�Ȗ��\	I�!�; �O�xq���;U�2�t3��f�L�@d�׭1a�����h�T#nw8{���-�����\%
��=�+g�1���H:H�����L� ��r=!��	��"n�8/�H�I�_?m�6�/�$�_Ŭ�f[�QZbrA
ɫ�mxE�	wt���X�E�������V�P����z�Qm��߫�[���o�"��P%s��RxG��w0okEP��X��V۫489^q��դ����6��v�1���4>V�H�>A�w��2q�8�3E1���"��F�&�B�u���%��~]���&),ُ�ʍ�n���4+�)�LDmZvPt��%��qc�ی3���qt�ޣ꛸|�&��5q�j>p�(Pرs�c����}��A(�~Y�L�e���Y�� �A<�3�ظ�����q|�{�&x|p	Y�M��'QWā6�/5�Ħm�᧫��L<?���>T����C�z���ФY��?��:I����ɫAtMc�ޅ���Io�����6�܂s�n�MU��P5!�~ @�9z�h �����)z��W_S������G{�z�C|�A}���UW]�� ����Cn�,�+��2�4��@�B?4�Dft}��H�����	���B*�%kVv�XG�lq��(ܹƋa�Y�j�$u�\�G)8�엗�P���.C�<H�S":8o:6�@D����7�ӟx5�C�(�����oe`�7J�14}��׳8\a�ʅ�Kǋ���:�3�Su${V�c�S�`xU���3��A�+y1e�[�*/���T=Ka�1Q�0���Ҹ�-�-��J_��	)���X����ʞx@��]��'���7�Ս�)�и�����=Vy�(Noܐ�/��7�01�cL0��+0>�̙O�.��Dk} �����v��w*��/�h+����Ξa �5a3_����1����! �®�|�'1�#XCW(uL�QL���RH6lX��˖-�Q>��B�W�Y�BC��y6N�B<;Ϛo��m�b��(Әب�)�|"u�ۑG��»O��^M��*#-c�DG���`��=쀑'��s�z`)���R�T)��MD�R������/+ȣ��H)�#E�(�×�&�gSF|>T��.ء����PV�Yea5;^�O8˶��n 'T �hV4�%�7�s��__��l��fL�P��u�����f����G��Y����$?1M43.�oЗ����?��7=�mm+��tRWY��2�����c�%�i��z�5�/_���<i���.��ۓ��Ӄ5��w��3a �C�#�pQ��L�3H�D��2�{���{�o�}yBW��������F�%�ߙB�5�,��T�\��1�n �?g�[6صC��z '@�2hLh�cy�{����+j�����|������|�S���g�g�������=:�W~Y�T��t������$��W?Kv�K_9,��2ix�J�h�0�{��' e+Ł3�W,X`e��x)�sb��q^�U^:�q�ǹa�|}l�:�]��YFY�A�����_�»F_�܃���"#�AC�����r�}���n�͝"3}ܩh�2���4x��s)�X����I����M��k��""N��7N"��8Wh�RZ$�|�pԨ���)�^�;~l7q�Lu�l��`ε��8V%q��z�F�A�AB(;/g$8d��Y=f�Էzt��� <h��?E�_�v�*;U�|%��2h ;l�R81P��Jc#^�Aʂ��x�l(�s`��F�V)/�!��R��iC^�o4;tP����
|�zO2�eB?�7����/{��O�(L�U�(�A�G�>TG5!��J��[M�� ��FȨvv~'$�@�xÝ�;���̲��$y�,M(�;�}�.+�^r���W^qE���[ʽw�S.��R�\�S�0A�.��/�����JS�L$Y=c�>:M됉r�Ki|S~���C�G>^���  ��IDAT�RMm�Wl�Q�m�Z�o�QFK�/EK-Dʮx���NP�$�(�~�ڪ6�Fш�1h3��7^�4nB�4Zr�Y����`��HwD}��P~7�]_�,[Q���c��A�msn'�����;v������+��xm~��B��p��\���P��1�T3�E�VQ�d�?�e�!m-> �L���г;s�Uז;�K���ƻ���a��u��I�'
��1�ܑ곸]�����(��k#���--���j8Z�~��l���>Vi�M2�%��0ދ>\��$�]"^���,]v�e�R#�������=앲n��;Iԟw�P��'�G�U�ޠx2���6f�dO�̤�t�{8z#��'>�s=�ZA.�d��"3�5!ix7@�C ģ��"�ӎYk���<�����������cƣ!�IE즜.D>�od�lک@�����aW\����#(�ۢP�k���~�K_���Ǥy�x�8��w��痛Ԯ��r�w�[o���z��,�]w�Qn���r����$�7�p��i>�[�&zu^ى�cK/�o]�p���G���`8���hSH���s4<"��T�"A:l��8_%���q/���7^Ӈ�Yq`5��Xq�Bo�,��(X/�5�OD3�G�޷o9���D�R�ƛn�'�.�,ő��P<"� -:n��&w�=�vi0�җ,y`��ŗ?� �uz1�yv�Nx�'w���5���
��(2]D��S�~訉�!V)��a�/?�N�fЍ��&�אkHam��;H��AڦC<Î;剁T�zPn�!Ø�7M�|T�z!E7��,��C�摴5���Qz���|��SaP��<"1�4R��=�	e�+�<ɍ��H\�c{�Gp�sض�[��4U��a���7o�'���e�]V���|�|�ӟ*���ϔ���O��������>���O|�/�>��#�я~�<�����/�*:}�W*�09Y����f���{�c{�_�ŗt�7àL+�r����՝NPcH��(Gv�+Gw���.��xnm@��%:��44X��[6%+#�rT�
�.�5AQjc���C�s��]�s����:x�+��w�*��n/{w��1J�N>1�,ҏ��3��|(6G���J�`�r;p�S��C�&���L����Y����������a�{x�J(�#>&t�U=q���s��1_Ǝ�����RJ_8N� J �2(�(��yMs ��≝0��J1&��=�a�#A�3ߵ��О� #@ܿ����M��n,�|N{�����M�\��yDĊ�S~���4	��븋���_�h������P͡��s8�?>M.�e��9�=a+&�1[{E��%������j�@��IO�&u
�f��ع9aٲ�>n�����*>z��e���~��p�#��2���8�#7�.�x��ؕ�^�p�%DS:A���'�1� 4�U\VH#M:�=4X!e��+T@�=ipa{u��1�l۾�g�x��x�����*���/�����ֻ̘�t�wb<'v���Z���@)�y�:����/�]�W�8��R��}��b�l���v&��ͩ�Z�(Q9!���:t���`Z�۫�Rr)�鎕=�7�Uv[�->�X�Pz)�)�]H�C�`%'����Z�j���d*��p镇�a �ĀC��0��#��Ppc0�W�Vn��F>��LZy��o�j�z�Y�1�%/OڰU������Ʋ��o�ӑ4�W�����[ƪ2� ����׉)�/л"����o���裏����r���{��{����{�k��:ǝ�:�h�-��,��V�B��Ɠ�[Lη�b�m�c�����C��t4gw�S���.u\e���q�F�q�� ���R@��B^cE��x����R�!��|�=��9�	��ATfV�GQ�J�����[���]���*�R�Gh�ٳmG٫�����҆�y����.�k�&V�Y�/�<���;�7��~��E��P��{���~�.�o�G���.�x��Ɨg�q��@�P85��Ɋ.;4�K3z;`���0���.Ys�|���a�E�@������׊��F�I<��2&����O��G�U�j��Nud�����A�H�Dp��~7�4�R�΄�n\����{p�f<���.�_7����؄�k����Nz�u�~4T��\z݄O`���o~�>�����?���7t;��	:�I�jd���0�����f��]A��%�C�ԏ�S�4b�9�I޶[�x���.z睲bժ�~�Ʋy�ֲ~��P��n߹�lڲYnq�+���$����������������ۿ�y�]"O�H�6�4 ꊂ���,n���L��	�(�|��f�h�e�����# �h@]��%� ��]���;,�+#��l���BR릏6�a6��N�r�/%�bn�������ns����څ���&��c�%
)H6�D���P�?:�~�ҽ�a \(/�2��1p�ρVh������.I[��*c23:O̞��������6�vzy$�ʙ���X��\g��'�O���
�4���c����2y"��$BN�8R^��Yq~�3���y������!t����UZwls�G�5�9L�i���|<%��o�:�uk�z��V��I}�/�1��۶K��%���WY�Q��IΥp����M�=R��eve˻X��҇I�{v�?�
}��M5�\��ǥX+�ރ�Ў������ݥ�^��l��2갈9tT��*{D�>)�����(�W]��̚9�uɑ��6�-۶*��s�v\�l��=(7���g
��5v[�vCʰ8h��"`��p��B�)�HV���/ye�p��e��^Tٹk�&D��8�Pz�ͶF�(7d��MB�_�0q���?LG9��ؓv�S� �
��G���[쬰��8��v�Cϸ������*CtS�ɑ�L��"@;��&L�)������^�h�43�3�Ӊ����]{B��OW�y�;H_�d��	�[ӿ��;�ޓ�ܓ�.]�zH��v@☺�m
;�g�9Q��9��P�,b��o|�[�_�b����+)��,_����o���� ���+;�|b������n���"�"�Q����>�mf.��LƁ��|��5��C2Ō%��3Sp�,E��^�,Qi|�f��-�%K|�w���r$�7��|�M#�
�����w�xТø�{�xUx�L:��O�A�ʒ��@oE8|��Q�L� �\r�%���^`5gƌ����u���l\I*��ƴ��4O\^2�ʵ�FS�6R�'ti�8���#,�Xl��RǪ)y[�i �N���[�{b6�E��p'L���l���U�S'��qt�|�moٵ�O0sV6�kkӊxX�C5���5FC[B��� g�B��>�V��b�e�2�4�/h�<�I��;���o-F��M�yE�!3���<J���>��L8���&��2�'�P���l��پs�=���JZ�j�_�DNI
�B�Ąn�\$^6�,;�|�)�@�1E���M?�_}���8�noi��_���+Vؤ?⥴xK}�_$Ý�������\!�����P(Ao����Ы
*�1ś��L{c�6�K��k(���I��*�R�����Q�Sn��a�{DHx�Iyb�-7(�B�Ҡ��m��1R�GV^�ھ�ڶ����)����q"b��1e���۾�J7/�A�^�;�r�#|v�8滵�K��e��T�K���:�< 6x�nv�-{���� ��_�����p aegq�EO���'�#1�DE���=z"W��0&bCyS]*i�RM�b_ ;�������j�`� ����#��$e�3����B=c!��d�>e:�an����D8�����<���2�V|��j�,>K+�:���x�]�}��>rO{B�}�����9��U7xԴ��uO}�0����9�:n��_@�맥�>:�~NV����.�6M���A�f&I_�z���)�����j����~���=�x��g���n�9u��פ���7nWJ�4�E�;�Z� -	Xɏ����#1W^yE����5���u0t
ӗ��@nUpɌ%i���5���#E�������	�U_O�7�B���_�w�W�Z��bk&g����ʠ3t�X��<U7?���~�7�Q |6���=�U<p���k�ٳ�rr�=�����.��
��[�P���":"��M|i��6�$ǉ�խ�Lt�;!+?�(|��5�VIn\�ǠɊ��L�/Z�
(:�;��t�S]�=)���s�
A�k4A�;3�.�qz��B\�IM$�R��l��%`Q���Y/���,�N��
�R�W�Ոs����s��q�*��.d��G�S���4t�e->��]�t���z��5~b\=����)Z�?Џ�CQG��P��@�IK��ԏ;��8B�q"@f�͓=��N���Gq���g���g~�Ly�ɧ4)~޷1p+J.+	�D?���㥿���������~� u7V��*����.��s����s�Z�9�*;�6)�2�Ti���<�AM�*�v�)�7o/�6m+Gv����f��ce�R�ޗ��G�ڲ1z-��Q����
��]8�Q	�X��3�t���bJ���!>t���9�0O��y���E���&(���W��|��"��{J�2S�yw�u�鸾+�]��R�u�@<����e��Y��ص��`(���j��#�@%X�mƃ��*�Ad�K�"�cu-�@���~�]A~8$��.h�����q�'�
j��l~�f��t�If�x���	�!���3�#�{&q�'^�7���څ�w����xM��ݴw{Լ�z�t�'d��� ��VEwL�� ��R:P�����)З2�������Ny�2�s�
�l�-���1�M��������VJ.B���-\�Ǚ	2�`FHU����-{�̎�1{��r����7����;o���[wsi���I�KS�H���Ͳ$[����(���C2A2@�5pl�`���o'QF�dK�N�\$JERܷ��}�����s�}��y�n�J&�y�zj?u�ԩ�Su�ֽ�����V��:0J)�}�t�
_�U qҴ��x��!0܏�ɉ����{����W�W��O�I����?�~�7~���O�t��|���c/�w٦˼�{�%�-\9I�0�Cڨ�j
O�����e�I�|���Iثb��1С8� �.U�C]KH����"B�|Fa��!h2VtQڰQ�d�c�O�m��?�H�|-�S�B�L=�ⱛ���(���I��4:S�`�="�CZ�+�Igژ0�G<��3B��Y��������1�ֲ����|v����VxyS��R�OizU_������'R*8���`��m���_|;��<��A���fŔ�@�Q�*2ɠ�p���Qȵ�/�I��?��ꯤ�IT��e����\h��s�\��s����i�˚��;>���SOj!����}T��'8
���[�}�'|���}��U�Yq?���͛��y�D�J^ߊ>Ө���o���=�vu�=�lwT8P`1�]���hÆn�d�Ʈ}��Q;)�"/�8UK�k�t�W�r����W�w�_����{r��n�ݒ�'�����]��[sZ2zB�&w���C(�G���u��bv���N�F�(�K�������]{��2���(��\r��FޑMv�Pt���пne�}A�\�-�F��8 ����Ɯ� r��N`�?.�.�-��ݟ�;cA?���W��Q.��y��������LP8�Aܲ��'c��O�)�=&D�q����TY�� ��O�0�>x'L��i���v�F�_X���b�$��Ώ7c�Md��?�g�[��8J�3m裮S3��o���li���g�1�:�`�o�4�G����+�1�����|��O3����T�]�V�3r#���
V^d�[��_�[��0���cZ���[����@�����S�%�	�G5v^�].]j���	�V�	�1����[�ġ��>2���R`Y��_���y`�|?:P8+::!C@*��ɛ5}���~�~���_�5)�����o�F�k���ݧ��Ou��+��;�������2�O�fא]�|���GscL��e3��H�/�p.�s��l��/�e��#��]�L��~���_�_��\wϽ_��Q���&���M�h���\־�L����y���(�y����[o��)����`�c����E2&t���.ғ�E��L e2)PF���e��eBQ����7S�	P���	~NCK�`O��!_���_��	g^#^�W�CBLx}�Ae�B�xfe؃������f��Ms&�&�i3���I���3��cxL���e�R|)�l�'m��r�A�J�7pA//�����̲S;6��.f�[��h�[�I�����>[@������ڼ(�R�`̵�<���[o�ڭ;�<˻��8�3�܋�}�V���q	���,:zR
�n��cݢ}G���w+������[qDy�K�ݵ�;,���v�{��{�w��Ko�8y����6��Q�7�ɢ�E��x�������]r٦n���L3����� d*��>f��� �*�G��A�&|��m�j���ay�Uq͈����D���w��Rf����c���p5<�~m���X�|0�ق�e����i�iH;��a���(+�T5�?���=���r��3�	:1��io�0�y��1u-�ߒM�f��\}�5��~�g�_�.�?H���_����������g��v�4c8�ۥk�/�N�Ud��R�k`�<��`�kmT��l������?��L(BQ0�l�Mb���~��O}�#݇>�������;o��V�����Ї�����w��G}�-���W_��r����8�R64T��
;!�nq<�e��\g�y�)��t_��_��1����{\&W�=�OG>���>�Xg��e��E��e7����H �e�<-����Ɓ�+h#&)�z6�����E��O��5���eQSn��c-%�H�L�qʘI5�L�Ʉ��/��]/���L�z^�"�P:����&�/��c����DoP@�O�CQ��hLl2��C�L����a�T?!mY[	���[&�<B1��9v)�,X`�'5�A�C�ȓW�L��.�&����>zΨ�>�D��	~�w�J٥�r��~76� s� e���p�����$/fY�)X��� /H��<�T��3�x����f���ݭ�ܚ��HJ����|�r�Q��,떡8�:QDcK��ܭ��Ǻn�wX
.F��z������݉{��;�u'�����J�M(�(�·D���Z��]���m���o�|�o�`ǜ'e�f�(����Mj��D��X2�'~�P�4L������s@�=����z��n ?�{dPlswo3�f��?�� ��1�o�wlGqտM
����Y�EG� ���-.�S��X�1�)��q��n4�j���Vs�y�P2��Hܮ_3@�k��'P�*������O�Ӽ��ƀ��`"�������9	��6��mU����O�u��&n�/�"�F��Kw޻��ǻ�����>����?��v%��v?����~�'ߧ1s�/%�)�S��0�C�N��x3)�n�� zL���WfAew\2�`Ё��	�8��P�q�����}6�~�ow�������@w��[�M�_֎-h�� }��t7ܸ�{����}�c�>���>�sb�O��ǚMz��c��T�s�"�;΋so�����r��3?�pw���u������R/�=����P���T���\��ۄ�ur����"���E�	��M�(d��Nhb���A�0>�,�W
M��@h��S����(9ԁ�*��1솏G�9�X��<��"�B��p�.��M�l�� N5�CH^x����4|[�G�N)?���P:W�zy1���d6u�|�LN0(�cC�y���Nʱ�P�����1��(��᛫9%ks��INJ�G���0(���	����K�E8�GۋImRB���BH3�O�$=�w/t�bc�7a�G{���YV��� ��Ad{d�+ڑ����k��
�{��o�Eh`�?�n`�K���o��<�T����vo�uk����ERD���ǻ�uk��>�����n�ػ��̎���9���sз)߱�;�c�����νRt�u���vRt�y�;r</�	������򛅒O^�Ev�bj��>��K�W]u��n��3u`�������,�0ָ(>ү�����ʌ�^7��g�q:�%e�&��;;��L%�P��k���2$(��F�	�?�fg����^�a�)OcC�R��"}�'$�#`NC�f�ܸc�3-��Z4���h���iW�4|�MM�ޞ#���I�V�*�W�lzb������̾�Vn(��x�)�i|)��g�1���i���ۗ��U��5^��5_~@>י�s⚟x�G�ɦ�р1_l�6P|�Ʀڧ���h�	�9{����ǥ�������|�[��n���q��r˖k5�.��>�`����v�^%���]}I|	 i��\�ʧ�)��f��ص����� d;G�Y��������>�Ot[������+�e`P@a�
�_1�᪟w��]΋���k�s��0��1��8v����K&�aP~���Ǔ�{�ۻw��c�r��/�iBa��L0�0� ��onH7l&`�f�P�d���̡���^�A��"��Ne��V�:|D���c���a�92�Iw�v�e�s%�{k����B��Xa�W�?e�����Y���i��
֜�^�ż�
��v�H�a�������	+����³ ����5��$Dn��Y�4��%C���G��Ay��ĭ�^0���,nb�B��ʰc˽��|k���޽�m�[��8e`	r�b��A�}�;��s�~�t�+)�[O��< ��&�9��d^�E�Ç\n����?н��wt�^v�_,���7vؠ���2��>!>�z2)���{�; Ew��ot�����u�;y�h������I���Kl�e�G&�Ƨ�9bvy� ~eu��eݺ��u�o�ܼ��p�~pecg���?`�K�v��gg��I�j�Q1 �,�Ƞ�!�xl�Kɓ�X��O5S�aS�2���Rt���q��T9��4�7��o�]�h����X�>;��h�59��qb���%M��aV��0���������s?�~��_~�ݗ�|�o�z�����Ž�>����������}�.O���Qm��X� �ś�s�����ӄ���/��[��g�}�{�s]��� �:^u"�Mx��P�r˧��+gxD�bI��#h�ɝ�RB�1��C��:����}�ŝ�DEƵ2��)(�t-�.��o��6u��,�4��5(�o��6��`�������B�jk��:o�t�w}P<J�A)��g]9M���j� �WK-\VbG�
��"6]�ɼb�@H��=�2Y�5v
��Bl7
���n��$��0(Ɏ��*M����3������B˱��W^��"��Gvd5ind&v�@aTg�p&�_�q���&�L��jx�^�|��X���7�Qb��'����e:�w�e�ä�#;�Ֆ���Nv�S/&�Kn�k�����N���4��>��K�5��P�=y�+]W�l�I�q��{Zd�R���ݬ�ι>+E�W_MpMz2/|�	��qMW��Io	��{������6(HL��5�+GNy��Aܑu�;e����w��go���g�5=������;p2|f��O|�u�Ƌ�����]عo&��B<mN�sÌ�;���G�D�^��[BD��=�~��V��/^�U>�Z�t���E�-B4O�;'�~2�0����{X<��;�(�hf�Q����C9>�1��ڑǁ��s��[o�I��e�=cr�����_z�1�1�j��S�
;f���
L�r:>�Pxʱn��f�w�5����V��+���+�z����N�4��XN�8�q9
lT+��v��8��c��9%?��e���Zz���x<s�!��{���[ΛR�I�6V���_��6�mg8c/��Vr(Y��>�n/�Y�klbLbna���V��v))�Zk��<���'�Ѧؖ��+r�� ��In��`��$L���v+^̗�0OTx�p����E;��YP<)p��g�f�#l��sE��8᡽�r��[�7-?��퉬�h�� ?���;���{ꩧ��=��e���'���������Ow;�ow��p%g�{l�w`L'0�7��+lx�f>e��-�U�&e��)/����B��1VP4�"�f�Iٽ�λ�+6_�vVӱy�y��]�+R��~�ݷ��-_8��#�j2~�۶m�wx!�	�2�V��-�[i^�z�;L�� 6�� ���IM,t�U+Wwo���]w�S���|����J�(wlrv��:s�t慰�'2�p@�;QT^��񲈅���cq�Gߐ�!] Z�4t��ΔFٕ i�D�-��yn���$��Y�
%ll���\���Z���re喸iC:�N�ݕ*���Y ��t'�m��ΩLm �J��rNݨ�p<��[}I[�+<��_�T�ܗ)�Q1�Qv�8�@�g����5ɓ����ueV����\ygs06���> �����?�S��Z)���h0��kچ��҆�q%��!����� ���v�]N��|�me��fB82Ɨݐ�R�R���S�j@CNIK|���ʟ6Y�ǭ�fԐ�� ��&�9d̀�C&}�l
���(�,B�/%�r�d������linhY�E��W���.����z����<W]yEr�կ|E��W��SB�����w���n�ͷt_��[�h���۽�;��`��Љn�EݚS�;�X�Fߤ���,%���x%v�q�M�J�q��S�t��o]��;w��n-�vj������{%c{�w�4N;tċ��7vW]}uw�wt�j��d�GQy��4�|�7L�d��<Zi3ڐ�����>MC�pı8�e9�
�˷I��HKԢ��ֆ|NH��]��n�JV��=dmiQ&}Š��?�.����R��'�(�(Q��cp�(����������Dэ�dsl|d�z�"jCٖ��oFZ�e̯^�M����ez�W[+�U����h4i��@^��_H���7&�}���������h�y+������$��3e��9&�M+����8��ܴ}��fC��>�U8l��ÔVm�i#�=.�Ǌ+m�l@��9�����׼��������L�?�|E�G�Q	0��x�Ӝż�����ޙt��ő��ywv�|饗�T1�s�;
JK
N�V��X��)����>.e���Q)�$>���%�=�Pw�=�t���g��|HZ�3���R h� �� 4w����+V&`P�Y,�C�mF(=��<&���>�/.U�۾}��u�
1J�\��r�-�e�o�#anh�6Z� ��g�:W��W\�/>e%|м _(K#��j+0�όDGr�Ni�+y�F���+}ăɍ�">�x޹�"	6��J�
>��w��~�r��#�w��� &�)��5IC����],��O,�h:_z�%_V��.��ԗ�p�TS��8�E���_v�v�&��$Jip��we�"I:��r���;���"ń��֬ew)<b��Q��+���Q�������$67rQ¡�Ӟ���3���!�0Ғ@���0�4�Y�Fzvi��ս�����%��������0��/��Ъ�P�ih�Q��b�~�}�[�U�p��7$G���A��F�K��#�(u����e����R^|��S�/�w��_���q�*�?v�Q �MfQM�=m8��	�?�v�)б<I:o���B�dV.Yѭ�����E������؟����dV
���=v*���o\{nw��5ݚ�˼���׻};vu'�Ni����c��W]ӽ㮻�w����7���r1��m�T�α8BҎ��40�ƞ���ss	e'h��'ڌK�w�{�s?��|c�s�����8]���Iw�+���J?.��ȃoޱ�_v��������i�Ptm�/E�ڦ�3�	p!q	���P�
�cC���vk��s����1�c����q� �NU���
�^2d!nL��}&�??̇oV��)x3��
��vϗ�l�6;[�Ua��,�LO�=|�O�8P���U�W 9�ޛV��D#���q���fq�&�LU#}�ԕ΃�Ŧ(��-p�ḏ-p�E"�n>�# +��C��NB��L޼���w����Pb9;����u�|�ގ;4�Es�]yt+%q�&T.s]��:OJ���Ũs�<8�����<��A'�1v �
�>&Ǐ|�#� ٢���z�aک�L���Į�B	<�أ��`Q������=�;)(.{�4�?v��K�"���ĉ����05h���&Uޮ�>�fB�]�jMK�z�He֊n3Lx6�������F
k���#�n�'�*;qk�0�͹�P���Γ�{��l�A��,���x�����}+�ԭ�eS�2}���a����Q��h(,�Yd�4�v�Qp0U�s�=O���3�s�k׭u|x!ި�L��L�|7�����u�/��;a���|l)AQ�7^qȰ8�m-����F?�����m����Da�.|��FY�L@�7n�h��ʮ���m�.ݗ>���b�p ��Rp��������$�h}ahóꄌ�h�l�:����Z.�x���D:ښ��"���:��6���XX�X�f���
Æ��Z�t��ip^�A��4)��:���8z�[.�v���R\Տ�Y�)�?"�.����tk��^�R
�Z�Z�k����v�(��.���v{����m���S��
�9�z�Жk�������o��2��D;���(��%�g�~�{�׽����Vc��oT�ih#��ӱ��y���ݝ�W�Am3(��3���Il�h�0�`"����`�bd}��,UO���U:lp�_l��&r�ӡ��_��3�4����U�f�K��݂��?��nT��D�}~���P�*�R&2�О��C��Rʛ����]q藩���dN=�F���>*2�4���/��Ǽp���]�MY@�����?rρ��zTɡ���x־^ٍ~煎�h�Ie7s�������Q��������8��)
c	xQvy)�r�!�/��+���q?�}N�/_�a�C��4���T6�i �W���E_��<����}I����e�6�Ґ��Viv오�蜝�)��8�3�!�N&l�1�9�Kp/o�s$��~���=��3����n���v�7Zq<tHJ�&�Sl2�s��ʠ8e��"|��O�R(��t� ��13u(zPN����F&��uR.Q��	�v��^>����q| �(�|��_���9��]��]�{ŊF�xL�g�Q����&tsl��ɋm�5 r��Q6H)_/���Q�W/��1Α{���M)/�B�QL�*M��R|��QP"Y��8��u�:��W]�]r�%���oܛ�be�������K���n��=�Y'3�י�J42}�R�U�㠸r�G}3Ŕ�O�'�Wٸ��C�K�I�����Rvix����=+eW�p�2�K)������c�B��,(�,���ԝ���7l�.p}���*-��F}V��� �2�h�5���.���c!8O9֨��O*�	M �������G�#u����NK�]|�_b[.喏A`���Ld���p]'e�7:�R8y�����=��7�w;^y�;�{_w������\ټ[p��n�-�t��4�'�,��6	�ɱqO�Yb�vQ�R��q7�O���djN ��!Ȕwv�i���Q�;���c���X��s��W����@�T����Py�aiC��)���=0B9�`L�X��̉�1vKL?�(�áw�b/��L�ߦk�{��gy�6(2�s��0����`>��l��g���Bx狫���4��oz�J{��{3���ũ�Rt�3��3:V��6��E�\e7;��%@��<���{lOA��\��eXD�
�2����g���J��y���� : �-	6����v��݋��ۯ�ݗ�\2ᲃK~���Ñ"&7_/�y!l��x�KY�L���O��G,j�����BY�~�g?�Vʞ|����h��7u?����'w�m�_��:+A�E��1� ���N���]/k��p�
�e^�L7�I�Q����͗�Ѯ���v-�����uםݍ7ި:l�b��
o=���%\&�2�0��|Q��b��pz�c'��o/c�(�gk��rejM�0�F�8�ɜGZp#C^p��삣�s����鮐��N*�ۯ�p}Ҧ�ROnA_y��ng�{Vn�_s͵VV�����kd�+��n��n���-�������Ʒ�h�o���dp�q쁊�����g�խx�ɤ�1���M�� ��DY��7�{Y���Ӷ܋J�P
0,n0(z(�(��

6�J�� ����oA/���_������ �oYPq��_�Q�d\b�L:�c�iԕ��|3����>�`�'D2(|���:����B�8��e�Wp�ĂIÝ��`��w\3Ǔ���f��?�1t�kot{_��/
ܻ�;&%�75�C�Z�<�ॴc�9���x���_�^~�����^��l����70�Z{��[o��Gs6���'�3�ğ}�����i��8�	���_��M�[t.��XΞ?��fcIh)���?,��]0�^�O�d�o�q2�� �k>(@h�A&�x+������(����Q��p��J42�����`�Rv�3��V޹xڇ��a�/{�5�YX٭�$F��nSvQhzZ��+?�"e�f�:P����{3����*|��󝿲�7bˏ^���sZ��
߷g����,9!m:��Ǒ��y�y#�sZ��p ^$��Gqc r�M��e3�cAe�ɢ?���e�O+�#�D��7���0蟁��V{��MJ�� ��&8��ȷ��4�Q�d8�Fe+�9؉�
�sw&��!�N��3>�{�ߚ��W:)�>�3�C~vo��FO�L`(�4�[�d�q�ۭP�^>vq�M7�W��5�tv��c��2��!9÷T�;�{�h"l�?�<Q9nr`�Z5�h�g��c���(�����	����m�N-�"�BEvkW��R-|~\$�V�LM�c��0��"��L�k`j
��'�QŒ]J4��-_�T�p}��dgv��\��2�9nw���n,�*E��l�)u_"eW�ʎ�e�m�w������%J#ŘT��l�f�[�b�Q�y�/�d�ߤ��s>�i:*��Y%WR�:%F�i�������H&�~ C����6�Ճ��|�E�ք���gj/����m�x����H��벳��]n��(��v�ŗZv�����c�2�}���yRn*��OI�f���`%ş�G)�͵e�yϻ}�g׮�>_��u���*��]�ܿ6k�"Y�17J,�7��f���W^�^}�u-l߰�Ɠ�פ ���+��Wȱ+�ˮ��;�ww�E'u�?
_�o����8 h2Y،k����`�*�"cS ޞ�6Z�xI�Te0�^��Oi�箝��o5���z@c˶�^�v��U�7��ܶ���o�7T�
#-��S*��Pd�E��-Z!�7c8G�83���⛝��TBFt�s�2�b�x�F٧YHI&2�(>� aH���ǉMgi��u���M9��"!g�5�(]�Y �����1���+���c��Ӿ��U[SG�� ���5vBS���? q��J�ا�)��1e,m�q�8�I��f�{&�Moq� ��Qj���yV|շ�yV�A�e㉹��#$��&���S��"/�5��\a��ڼ2	�C����	̭��FI��/��C>A_�|�?f̳�I<��	�O�؟�r�N�-�������Hc'�8��7ކ�bw���`<�&<sz���yL�8��1�js��ӛ F'���g��(�jg?=RQ~�\�'�ͻ,l�(R�C�z��˸��K2�i�h�L�hDV����I:�>��}ᅗ4���>ǭ�,�0�ʏ��Sq�)VJ��N�r����~+���|<F�*��~��*}ڏ��qb7�*ĮW��sʏ4����lv��i��m�c�=ֽ��RH���iH�C�)1<:F�`׋��tB�n�����}�����P6�0P���\�ä̀���Y�u}iX�ۿϷ��6�y��w���jtWv�Y��a�E��N��ٍ�v7��C{�Bf��c���=�F��KZx� "t��Ώ��6�6��
����P�
(�93�N��I��D�oAUZ+�2>�jUS֦����F6gd�cS
��y�� �c���W��#}��	1��j�g7>�X���x}�9�xJ}X�Aox� �ןQ{�pB	k7�<�o�;)n�!����[�����w(|�V��b�\�����v���x)���(��9�-�%#�͓Ώ���ΝV Qvّ�5�r��b�>Ϡ�	�������.T[��' ��vխl��ujʐ+�����Wc��&�]f�<>C�޵k�oA�l����9��'�q^��]np9���H�iS9��������[��c�Y�	(�(L�[�~�Q�zZ�ˈ��z�;ӇE�Q�=$���(�����)vP��.���Ɏ��Q���k�D�R)(�[4V�q��b�"���,��~W�.WG���ہ�xcB��I>����]�n�k��5n����q�Ԕ]�ʮb'qٞ2�0פ�h���A�J1���|�B�ԣ@r���d�\'6�XY��z�-����[+�}�(����I��e���3a1�\�_�a���Ǎ<���7����>+���"Z�3ND��8�|\�Ys�����sl��
C� ��&���d0�������Ҍ�5{Nٽ�B �^4$��-}��=i�h��r�� �t}��W�)��"��0��ޜ�f�b��+fA��K����a(�(��;�4�����gl�������)W��O�yW��<m_X�}�e+CL|�}c���] B��R6=(��[n��~ם��_�J��I";7o�Q����0�#aX>�@�;#�jE������k��1&�@�٥�*'���̜��|�f3��ǼЃ��}��n�u��3�>��w|�%��O�EAA!�Oƚ�P�^�[�ϚF O@������-E��xfz����Lu��(�1����CG��p�Gx��`T�wlJ���j[��e�����Ks\�Ez��bE�yHn&�h�1ǏQ>�˜txlx�!-ׁ��Z&�쎥3�ncC�kr��%�F�51iCuIyZ�R)�~��R��Q�#�]�K=����	2J���xG�ȍ�H;`�',�B\���r�SF����O�%7UO�,L���}@� {��D3 h[vF��
�C� �T���O7���Z�n��F��B�z�������G���{��.qcݮK��(T}g���M���eE\2n{l�>��r�^�˫��hk�n��}R�u��i���T��Re�Tf,I�����`�Y~��|�Gx2�yk�Tc����:����|9��2a ߌ1����*X��	/"Y�+|7�|��6q�gt�㔶�E4�,�5�'����R9���{�=m<��-���$3�H6�灳��å�� egwٲV����m0��¸� e�|DQ����*mJҏ��.0��c��e@��X�4�(��y���o`��8l.�@�}\=����xC��!��&�܍����b�蜦w�����d��pp8��5�L�8~����c�g��0�����=���p�`�_0E�`n�$�*�N���y��6'����C�?�K��S�+%<}4T�h��F.2�E��>*E������0�������<��x�^�1O��/����{�a	��n��=ݗ��e+y(�@v�J`5�{2τ\;��c�K$|"��}�<(]?x��,���L���&i�ŭ��*�Gޜ������=�*��vX����Ｓ[�{AhS�d�3�e�胑(�~�u�]�ϹN&Ν;vj��i%���<&�q�<`���)P<���~��q��Q_�r���5��x @1Ҍ��_|H_6d��
Wwq��Łw�d��yw2
�X�$@�?F���]a��=�,�~\ԄH~T�ڍI�]O�t��2�B�J�o_N¤pf���a��L+
MF���'�)`���rk��`�晌k!��,JS�� �3�y4��DQW�+
�l:�;7�2(��:�Уvg�ќ���(��ɎH�*Z�8��� hC�q���y���R��� (�������9zD]X �ڽ�e��E���4��#|Z!��g�y�Q+�,ly�,qD���ow�|�;=�����t/����4U�!.u�6	C���R�����2�#�xD�I7(M)����&fQ�݅@b�C��}}^l�X�z���x��e�o��"�hd��;\�Ƹ�E�+P��s���c|�愕�r�i��f��l�(G}��|�?�X��l������/;�������g�`�>���1�g�ռ�O�����¼���9*�q#���F�e��C��S0��u+���շ��x�Ǉ����' ��Bm�Dh��<�*��Q��GcZ�O56Z����Qx'�`\MQȎ:i*�l�,UO�A��1\I��#����}��n���_�5��tD�����D��{L�Ӭ���!
|��S�rDޘ�q�v��΂��B��sP�}�;��c��؃���a�z$�l�h�5U�^x�~��F��o��q�X��8r�{K۶oO�=���Rd{P4r�.?s�Z��c�+��$�D;?8��:��cclPB;�1�3��ηw7l�~~e�Ǉ�?��&�c~|e��n۶����ĝ�ce�;\�ec�i>$��vw����D<�d`~���o~�~Yj`� oȳ�ʋ9�Pt��7��#�01|������?�������NcW��,+��A���f�ʪ��n�2΄�NȎ�;�#s�W�e�q�`�8  ��˙J)����<&+&���i?;d���}�;X4�;&Jvf��'/�>�mv�ʝ��J�b��X��e����R��e94>�Ǡ^
381(L���m�i�&R��nSv�ɳ0���~��B:�/��6�U��{0��:f�'/qh m��`�G���%1%����F]�rr���̥PF�U����+7���e�lv���_��
!7��y��*/hH�py��|���� QmF<6�2�C:7�G	EVy�O�9���xZ�o��9Ƴ��}���8�DF߱}��|�>������;��)u��l����ӏ�4�`�iy0�g��?�ͧ삟�%C);rmW�k���}[��b?6���b�L��r�ܠ(�(�<ة���l �+LX c��C���0�pƝq��?/�y����'F?|�w�����nϮ�^��]��
mL�@�b\ùP� pUު7r����(e�M��/.ew�ƈ�JiCy���>㺔�v�=	5~<��U���8?�r�I�8����F�1/#v�Ӛ4��#�W��	���/��ҕ{Z�Mڸ�\v�99B��^�M�4�|��+��拪���)���jG�rўE7�(���4$u� �c#qؤ�o��0rɷ0���8�3g��7����=�	O}'�A�L�t��$��8�1
�(rndŖ�sY���u	:B�]^df^`l�6�|3�2k!=�b��K���-t�'�4��D7��{<W��O�C�~�T�0�@��Tv5��p���z���N)�_���;�����Q\�L�a��Ղ�G��@�9C�r����<a��b�2�����/���&?�ȷ|f�
�<��%�j��n�W��]�AXe~��_���_��W_0��:Mz�Ғ���&��c�P灙�i���*3�P��d���/vu9��s�N+7��V����˺5(�7F:���6��Q
<_������r���y����B�j ^�z���?�7;9����������[������ �.mB:�H����&�`�~ؙCx3�qX�zr�@]�/y�7��B;����Ȕ Om�a��|���J�;�/6�I�d�[q�@��������atR��`8���+�ݲ�vhL��>�o�]dQ鏫�#+=��PJ#cy��`DK���B�NxP}�9M+�qC&;���?gd��.e�/�M�d��X;L2k�U;��(���so�������6�8�<�h����,����/뮻����Rv�o��>���/x��'�^z���o����f�oàD`չ�M�Q-x=k�3�0�΃?a ��c����W��ęׅ�٠;(Zqv܆�o~�� ��lʣr�71U�v��s�I�����j����&%2�y�L"��m;�k��/ǻ��rN�v�|nRmJ�.fw�c�ؙ��~)V���Ȉ��=aU��f����#]�0yFv�q64R�Q�3�Dٽ�;��x��f��˒�+~��R�8.�F?���%�	i���[��=K��S�5^�����m6�m��i"���_�'h�e���ׄ��̧사ܖm�Tv�-�9]�S�����w��}�$m�3�l�0�����/[��	�sZX����2�2n�-s}�b�[c'��{�(P�ҵ�N���W&�P�f�f��@�� a�;Ngٝ F�w��T��e��%�@�@�R�؉�5��2+����Z�16~��\�;,I��Jm:�즍�I�'͏;�~�v�q�z��o�c��G����#���g��*o���g��"_(�|�����Pv%�<�Vl��8�T��k�D�0�����n�����J����w����Oww��f�&y<�=�!/up�Z����$)��s���EG���?�}�K_�n+���d�0�|j�L���	��&�j ���/:),�~�0����}�����(�bP�AaǖIEe���3�<�½ :ÇEJ{�on���;�+4�p�E\�&�����4����V�/p������ދ���x�j#)*�t3�0B3�mEyGy�ԓ��q�A�ɾ
l�z�%�V�4�r�t3��ٷ�;���+�e�j��r^�Lv�L����p3����3���I�ש�t,�d��Lx��r�R�d���e�m<`0 ���C�F��@���T>���:7�W�&�a\d�eR��(e$��@�~��'�s6�G�|��'�'��p����������]޿�e� �Uo�#w�)OQ�=}���V�?;�<���-�_'����{��~�{Q|$'��<�oH�=e������*E�G�\���}��E�$E��xgA|�!��x���o:z���'�g	�Xm	�� i�z��ø2,���%9~<���Gژ���_�P9o��?�Q<�����v�稌#�����:aA�qc�6�������k�`�X�˻��v���'E۶��'Y���_}��"�7d͊w�	��yC~��dMM�0!c�M�U'�Oub���Y��Z=�&�B�xQh����ݴ�2�y�x�ƭ��ϸ���d����)-mTac����d�\�A>�m�ICJ������!�߸���%�e9*�2p���S8��ܶT��ӾD�G���3eh�>�*n��E\F�����)7���#�ug���׿�u�A�(���a��h��#6$j�)(~O�ZP��bE=L��1����6��7�ƻ� �q�cw �tX��N�+�
���F^�� �Wڊ'1��4Aw��7�<��q�7�z0�C�G�kal����;��h�7���,@[ϭ��x�+���|ƞ~N�X����z���@~�����N��#	�T�X�EN�w����޶��暫�WvIx��k�=�I�P����w_��W{�2BUL񪰅V�����y
�����{���C���::�_/�@�'{�a�t���9V��ys��_�F���W�7��L�b�bq���J���^�E��(CJ��n�OhL�0�Di�Fy��O�{��u�/~���_:�Ɉ:�l��]§�ķ��G�LL48uc�`7�{�b�r�r+\�ŇPٹ�)vŹ��o�K���/Y��f��vv��}��8
�ǋa����^��~K]�7Ji�%�r
}���Qge�Ց�	&Lv�P`��Z��5mȀ]�R.;I(Դ%2�`Q��漍�*�lvCQv���������V��B�Q�%ڥ�k������wi�4�ҳC�b�ly�҅��+����r�zp���#�1-:��s�<Aa'; KqΖ���7R�1u��/y]t�F�Y.%��rG1���]y�5��O��?� ��C+����WK�D�����׾����}��CS�a�03p|�2�3�<6��,j�I^�P�O��)/|�zK[�g,>dM�e�8; ��v�6>��$>�7W5����K>�X5�#�$��>�Ԍ�l	$叕�
?�1� ���i
��ry������joT+d�X;�K��H
.����m�a��0�wUv~�w�_zj���9��!jG������d��������|)�o��_+H�aq����LWe�)�o�����o�p�kaw���T�66�)��ԫ��<DA�_T��Wl�&hI���Í������*4���Ia{����da��l¡q�o�*���܌�<�{E��|�+~�t��g�d�������n�����.cS�7���V�Pe`�x�m���i�!/��G�w,��e�hQ����m�q��?�Cd��ph�F�v�&�{s�&,�Hq�2�*�(<]c0��c�m�3J#h���(:_�es��"-��#��1zh1j�<��?rH]� ��IZ���5�7�ܼ�{K�Ow����6�W_uśTv%�/������ �g)��2̸&�˥�]{�uVx�����(Z�j̊�/��cx��ǖ
���t�����/�.�|�@&:��À�G��/:�O��>����hŎ>����Kcq���]������s���OWq��o�Q��}�s�˯�����a!)��Q�� 0��2�d�4o�3��p^a�L(��m�U\|�ق& ���3e7@��#��;�,0��}�QFСc��]�hQ�8N�.44��(%�|>˭rh' :6]��J���"�QL�|ʏ�N�Z:W�ކ�C7
9�
m�B�� u:�Nv��	U>;�C�<�k
2����i�2�D�x��2��%2���6'�4��U��c��.��\W��h(0�$;"Qv��]�β�2������������ݾc�aʄ?,�hCx����.s�<t�t��r~V��>�C-H_�$�"� E��S01Pȍ�?��K��.{�������p����7��|�?zwZ�g٥�L�=��2~�W?@�N'm�L$����&8��->x7����������	�M�IQ�3���R�����|�Wl����#_�ҥ��?Gix�ceW���./�ڮ-gO5ں�ƥ���ˎ�Aj.��:P��D�_���1��mn�D?�E*{8t�8�t^6���o��e���%0�2H���;.��1vL{��n�������r\ra������M���dhT�1�N8�C�AD��@Ѳ��X�R+P~�O��)	���*���~��*�-���O�USn����S6��]�'<k��ב)��0^��Ţ��Yp�G?`���E�s�����q�4#դ�A�N�5�7���� �~�F��k���VO�q������2Q�����rW���|Γ|6�S�OXK�T9Y�'��Ӹh�sn|`N��ȷ7B�φ�2�#��F��J�F�m\�y�٤�+�h��!K�jV���M��O���]F�0 ����ή����}���n��{����@����}3�]� ���x�/&Q4�Qd�!���|Η��>��ww�y������5t&_S%%�g�Ō0��������#v�P�N���K@*K|��ϝE�4t��������t�tFV������7}�AD88z��}�{���mE����#���:�]�ʏ#������2����������R�5����!����d��˖�H���UJ
O[pĂ��i���>ܼ<���+�8���|�f�(�w�]�w��!Z��yEZ�E�o�oK�����J�RH��EX�ujc� �$�#A7e1Yr\�~L{�Q .� �q���#����ڀ�!(!(�x�L~h��n�2M��Y4HiNN�#Î�
-��|�s���\�T�/��,�Y)EѤ��r/0�t�"�ϤcqH�9v�b^��@����	��q[@�'[y�l\��Mi4P����ԧ>�6|��O��O}T�Ѐ|ӎ��xP>L�ҎݤS���_ɂ���������ģ����E�9Ud&��7�d�M��Z��\^Զ��S�*t�,	��� ͑C$;js�Ʋ��Jݶh+|��D�$�B��<�A8HPY�ag�:؇sv&��(>�p|�[��]�e��0��1��ӌ3Sa��5�4���8HUUk��s�FJٍ��D�J{��C+��mG��#���<pqqW2%�L��� >u+z�qa����3�r���N~���V�L�>�(��xO�穖oP�������EX>;͓�l���PvՖ(�|�����1�9�S��"�#d���&�����\sv��榧�kH�ํp����O5�%�d]}l�k-@ .�L��i&�3 Cej� !/I��5$�	�o�&��Nf�/lv��`�-��9�<����<2d�6��N��R�G�]��f�j�4+��z(��s����+ZBY2��"SC�t]<���� �<m�"K�8y��ʮwv�^P�=����Sv)��n,U$�e�_p�z�<v۽w��X��6/l\}�5ݖn���R�a(���	|���|?�s?|�,��t�:`eN�-�ij�؜;�8�	�����X��%��[�Fu�Rj����[��%�Q`Oy��>�����w����؏�٩�L1�#������1p��;4��A�\��vx�΀�fE�	�i�N���X��*4h.�`GÍD�S�LX"=В�I��hw�嗂��v%� ]��G&��J������萡0>M���'S�x���/%�eP/�+_�Ɲ�Q[P��5��2�[�����Vt��2�B<@��F�>��@��b7]�jw��!�ϠA�"[5Xq���������G]i_ڀ څ6��L$�c�>�ˇ�"y�a<�����^ъ���~�۲�����?����M��6���T���M�&�c/�}z��&aEIsVy�O��?��!�-��Mv�����\m�ɮgp�#!���E��T|caDaLb¢M�ЂK�����}�����Є�!%�(k���<������3&�r$�����7�U��~u�l��:�v9��:\�f��F��=?�/k���_�2%�j+��{��D��U���I\ڃ:����nT8�9Pk(� G������U ����͆4&��n�Z����E(�(��'�w��^x�y���_��>�%6�<F)���B�e�|�ȵ2�	,��0�O<�Q������~A���1�4a�z�8�N�v��6�	Ȏ0��ii������1�R�ڀ Ȳ`���|�he �甩�4�2���i`��qe�L��P�ǀ.�c�_OdYd�)(��hWm�a�z�P��Xܫ/��|6ߘ���3���zqȢ�xGP���#Kmh�s�� ��v�O�xZ�����q����m;�לI�}���|�.�����Pv��h��~�
s���iڼ@�QP�@yI㦛n��}��ݍ��*//�����#/�|��O�:�Z��JR�qE�ʠ��9��y���P4�I�d��x�ۢ'E��_�n��sc�:YS��D(8(�:E����de+^�[w^�����̺���r���V�h��E=~�]&���2rf4u�3dѬ���2ٴ0[��i�4:<t6������P��qgp��wB��Io�
^w��[�i#ʇ~�AoH�� Nl9N� ��L@�O�HB�ۤ_��N��`9de�ʜ�ۙ@�N;x0Q��|�(��M���s��j�)}W-Z4@� cqe7�_�\קԟsP���=�2���~�R�6��(lL.�����?~������R �'n�Xu��r�4�'�Oٿ�?�Nw��*�b�o������7o�c�,���o����2� p�Hd%.�T}�N�V���a��r<ǯ�����O���ـ�xc��I�LL/ۄ�i�C|�r�~��K�_&�(E��#H�Kv�d�Q�W�C|Ix�7� �N>d���o����k��޼���Z�N���K�x豐p�&<��B[�q����˗���t)B�6�|�v�/9YD� v́�>hKZ���kF��ie�
f� ���4�cPZ�W~�U��(C��3���؅����8��d����g��}�i��9JG��jng�4cв���#w��y��'�S��`���Ø�����lϙ�c�ɏ}Bs���D�)7�r���}��1�2����w�VfA�=�@x�0w��ZR��a5�f>	V�r�>���B�o�ˢ����1�tN��^
��L�)��%}�O1�(G� �Rv�#����-VPv�z��K�c8�^�}��u�@�Z���VI�K��n��˴|��y��yhː��e���l�p,���Y��ήVm�6�Y�.QaT
	��J���A���c����+�|G/ ��q�1!�@�9	�����]��-���j���%���Ҋ�	PA���'����pS/�U�����+��~��48���/�'��^�g�.*����\}E㏕��� an��|�@8[���
��N@� G�a\��/Cv�v�4ܤ)3AϨ>�gْ?���@0Oac�7v�50��]���4�f�%^�L��H���M]�ɪ��l䃰�x�d���� G;9�[�]���
��o��o��]���?�g>�G8)��}aw;0�=�8~�$��#(t}�{�?��q��~����5��ipi�F�_~5I[�8��D@0���[.�+��*��4g���Y�~>T %Cq�cp�fFj�:���-;��]��א�R$��Qx���&&g��T��D�
��Ի�a�
I��hS�ʹ�|8A������1U���K��6����J�#CR�r�
��ѣz:S �%�>�.s����������O�q��z(R,|�|�AiM���fW4��~�Sn�#�(z��!�Y�w�%����#�񣇻���n����u{���1���xC
��u(�,�/�t��Q�zQ�����L����������� 4Q�8���:�$JØ��:	�5����N���Ru���������cd����d�G���Y*�m��2(m���gs��5�'O��.<�v�/_���h�J� �<m���^X�{C�Y��Cug� .��#����W��櫌�5}�j�{v���Z�V��1��9)�#��V�܊_�>Z	�Y�������}�{��[o�bz��Pv��z�;x�?���k�Q�������n�Y���� �'	p��(����ώf�J11i{e�
��hvazf��Q7���p��B�ȭ�j�F��XSv��?���L�R-C�7�g*�J����Ws. E�ybי�yf �����O��]����lcd�:#Sz���$-P|�E�앣T�q]�cd���s�ؕ6	p؋�\	��')�B�ap���)�&�Gi�]x���JI�N/��"��㷺��x����/�ſ��.+hn�`�`�#����1=���'����[�I�w�9ɟ�2.���bW�`\�*r��g��Տ��m���8Q��7����1��E��3�c&R.��] ?�����e�JV���͗o��nÆ����dZ��V�2��IN�,!���<~�SJ�+�h��>�;&�F
GZ���kP��UZ�1?}2�`���3h�(��e�X��+��/*7�����p+=�%w�_B�Ij���sy�� �T�qJ�FP� (5(�(L\��}�;v�*�Z�o���C<�z��׭D��`n��x�%�c���Rְk�s���Dox啗��.sꊕ��O*G��� ��9<�N�x�'����JJ���C��Jڤe�c�R�o��P21 Oy��pP����j?���EO���K�#�<��юZ���"����2�96���;�e+���'����7ڔ'��N�G.�I��&�"�_BW�7^���q���}�W���}���o|�փ�
G�}�	h�Ki�����o#�����z36��r����_+\C+N �(8���#�v�OمI��2m�5=�A��ٵ0H�6l�D�|�Ð:	�]3�p�Mc�{s��g6Y�nԟB���Ǻ�_����������+e׋�%,�K{Z��wd�+Q�g�8K[���/�� 2������ַ�˟vg�[�����S;�(Q�zA��:�����9��Š3����s2;%$P�L��	������������R�&�d�v�R����YPe��V<V�J�=q�h�j���W�����~�'�����}��c�[��&��}&z�p�	>�o�;�E�yg���v(���)��� ��D�8�D&A���F�ғ�6N��0�_�*�P��-�k
R���fڞ�{����S�b��F'�^�K�򪫺���c����x|6eOy9�T;_d�ia�{�9�>r��o
�O¬D�84e9JVS ��y3J�y���@cd�o����g��\��K�
��K�l�P����c�����qN�c���]N�s�JN���&<�-��;7
�Z�~:̕@�'G�rL�{�O�dW��&>$rL��.�#��{�4SW��,P���G�X��e7J=/�c�B�G�K��FV���Qr�N1�ɦ=)GlvF}m���V��C��g��
�����<��5�	Ui�.^��=�v6o�l��&�r�_�� ��q�0���xn+�����.�L��E;�|��3�(��xhy����|,<Y}`�x�n4/#�Ӡ좷<���w*�	��PSt�:���,ѯ���$��e�n�^zwoǬX���g�B�����-��J |��u%��|����.�U�V�4.�ZA9Lw�LU"�m����|�y��!�R�s\L�V����B��e��7��B�$5@Z��!!���T��g�[ ��5|N�0����j�-I/F����$y�|g��2s���0�� �d�l2h�& oɅL��Ig�d�{���C��k�H�2-��@y�8��2)���-e�՘P2�f�+TW��}&z�p�90�9Kf1=0�'H��p���Ή�))mF9�t(@�>"@L�ť��C��C���G�ab�aU�P��0�]Uނ�5?.�����8�v[�d���_�v��TZ���5�E�v>�@&x?�_&%X�3'qk@ e@s;�����l++�����}QL�A���rtB��G�h�"t�h}[��~&Z��T����)��%D��C��D-@�l��(E��n��������������D�8`��<+���ɝ�g ��p�v��3�we�"]*%p���y���:x�{���^�/��Ʈ���#\h�+��'mB�ʾ��-�-7������/|᯺G}�?~PJ��	_} ��7���mv;��n����k��;6���@>xt��=!����WV��^��_�"G3���(�+��&4Q7d�Z>�`�_�����֎ ���Od�|�ٌ�=�b�ydA=U �������*��j��r�#\O�-���qޚ[��K~�Kq\����t���7|g2J2(3�i+b^j���]P��k����m��8�������(qȣ�ݭ�J����~�j�a�A�?C����

��@���*��](dUȤH8�D	4�[�(~(��kg�"��RvŃ:�p�X.E�ϥ���1��8��A�e�lj*�+3�~������L�KB!u(�y�(0Vv�y����tmZ�X�����ǳ�=������݃�����z� ��5����=�܅h�p�9P8gɫA}.��� �Cv��<	���p��n���sR�(��?��L ��	�c�9��9�r,�!���[(	�/�A9�&#	��A�*=�/�q���u��)�M����%�[�ߚ{���e�Q+�LxF<�ˇ³��J����K�G��
�	7+�|����0�hCQF�A��xnр&^�b�C��+�(~�4Yi��w&���( ��O���x�ܿ�Y�ԁr�X#�E��J�u�G�,�@����{�2 ޜ��|N��4�j:nZ.e
%���|�;�9������x[�>�
�p�G�Q�xI���ֽ�]��>���}��_�GS&wA��Ja&���&�f��||�]w�]�O���������1Mv��{�ym��%­�i�Ĺܒ_��oQP5&P7���w~A��
��]{ɐ��Uڻd+ʪp�zژ&�@?�A�%=���^�[š���*��
���	?��(�>��B_|�٧�=�W��9�>'�Hͅ�ի��Z����2|L+��H:�^q�7��͂2~
r$����޻����L;��K�����=�t>���]V1�����nV�ZYj� �Fce��
J�cL�*0�J�'��w��4�P<bƵ���d#��f�# �,�T��)�.����8׎��'>�O�����{����|�����7��鋓#�hp�R;GWE[8U,)����j��mH5@���Җ@�*�g�G�30���	��oz^�n�1�*�������4��BԆs�	v}g�y��A�
�'�iB;��J�G�3��&��4xݓ���Vr汤�C�OhB��������;�t�����=_�G?Ga�#O��e�ᭈ�,��7ٙ�a��U���� A�A�H�r���v�=F�2�_��Ĭ!-�"$$�	�
��z*8YM�a����hl�������઎A�(�u�&�F�p��n"sK'SC@�Z�l��/��t��N��+h�!�w��d[�L���B1�"
Ċ�+/%f�U���S!�I(m�(�+�RF���{���4�m���R�wiU]�	v�
j�Cr+�Z�i�H��)�����W��ʎL�����Rls�8���rō�=���PtY��G��\�q��(��?i���Ƹ�=��6��L��!]׭�"=�1�r����PS�(�q_u��ݭ�n����wu��g?�}�+_ռ�S|�t�w��p����H6��cj#����[n�Ż��C�Y���);�Й]��V� 7���"
g�AR�0�PG�2��^����1�����:T<Wג�2=�
��~�����YL�x��ʗ49ϻO���^x^���;��*Bx�g'6}�r���UUnǂ��?�d���M����q
�C&���7��\�od!qQF1d  /����4��%q��_n��6
���y�O��?�����e�a!j;����G (�k֬�x[��� 4��ї{� �Va�+&�'0��+��� _k��r�s��<�����]�CӢn����w������|w饗v�����=��7��V��my9��ND�(J�Ҁ.á4�i`��o�`шG����z ����t�R�� � �]�Gdb>����ݗX(�$e�v2}����rf����l�Lc<��4�j6�|0�#��&�*���/�5�U����/[��*���+7�iX��0�ho��JǄ��~����d�����6&;�QXq��f�v�ؔT{Ό���`�G�fR0�N�i�$�d����� ��J+^�2ׂ&�@u2�h�R^eH^�����2=�A��*�l(<g�	Z�9֘f�Q���~SJA�H�����Rvʴq &u�.
Z^f�ba��;��Z&w.3�A�Wt��GId⧞Y�(�h���&������ч2�>$
���e��Y��8i�-07{w��J\�p��^ �ؓ��lu��-i��i�=�*l\Vƈ�Q�]����@x�x��ω�� ��V���.
ܠ�r����o�rz�}�k�|�۵�u-h�Hi[2��褝�K����]��A��u�<_v�e>��ȷ���ݷ����x�Wc<����О�JA�˸y�=2!� 
(;�}{�1���O�`��Kʗ�N�����1J�9���oy�����Pv��+H�ؾ���Ox1F!���0�h/ǅ<��vӦK}�5<x��vO~�{!��ס�?J������O������c��ᚶ�;�ǌ�q����Sΐ&�iuR���Ƞ����j���K�k9� e�����=�;t�Hvv��.BSZ8
��[Qv��VP5�;D��o�@�։�|�C�'?�I���i������_븠_�K����'��
sy�G�7��7ϒv�g D��E� 4�0��`�ۨ���QPQ��Ҁ��B@���ʟ��A�`a�f����A?.�<����v�m��ۼcP/P|�, Q���,U��6���'`n��7S�0_Z?e�,�t��4��c�*	����_�nݺ������S?�d�g0̈́1�C����,�d��=雳���?���Q2�h���4��MQ��|��͸��r��7�L�=�=�ܴP"�)�.vΙ@}��,`F��x����ӻ��'?�q�6"���H�FW߆��G��%���Ҙ�8�| /��E�[&�lЂü0 ��#�(��)�{91��{���F)�Nd�<�ytҴ����,8�R9F��H8�D�5ǁ�� ��������6V��_����A�]6(<�Ɖ�ñ�O�m��@���i!g���S����~:#��<?��Nx��&eK�̺���"�&)��?�B��k���D��eq\@i4Ryd�X��ǢPHyEj�1(X��+�.;���%>��.�CJ2}�zRe0��W���z������2�p�+\�(	���a�؊62	�'Pf���պsԗ9�m۾�G >P#����ChK���Y���=��8�����U4A���}eG�2��_e�p+֫��;8��7܄Tx��r���������E$c	|�&��n��ۼ��n���nQ?	���9Ń��t_�җ��ʮ��͠��A!Pv*1�����ɔ�����D�R��XX���g����D)S�=��KOWl��Ds���#4�Y��{��?�}�c������{�Ǻ;$|�xī��]r) L�h��]*eI�,b����"�^��:�ڒ�P��8��_@G�������d��x@����;.s�czIGX�qv�M�|�� 7pz���������sz�����.���#8{�.�YP�O t�S}�6a�6p��Ru�t# ����K:vJ����[ݍ7���C�g&���㯲������_6��8삱{�pڬp}�<	6�'}v\��K�u
e�*��{d0�p�vA��G�4;a)��(uI�1�bTO&dv&��$�i���A(�2�{���,��أ�xj�o���jP�r	�ݧU���*�n=%p>2����Fp����S�@�c�|$\yZz��SJ�܂\$�|���#d�^���x�׸h�L���ݔ�X�V>�}~9\^���DN2�YQ�0�
HK~C��!-o秬Ax%�ջQF���c�i���Ui ^̀�d&�@�&r�#��ⲻ��P�8��fڡ��n �hcT���;	㪟����V��? ��]b]�6�'hn�cg�4�9M��/[a~g��52��v�V����!�ë�I�S'��Z =E��/���,s0Qԉc.жZ
��g�}�Ŋܴ������[tʦ߅6RB�	��ܖ	��!/�0�.�<�-�m��Ke�)b`"M�$n�*w�j�t����˘A��%n�8/G7���PT��/bjG0(�K|��_�b����o]�!�03]��V�&�p7���ـ�5�H� 0�31��݂�FY4Й !$癷n�ڽ�����?��������*�O�Y"���BC��rs�h4��F	�"z�(zL瘯Cm*l2�$L�� )��5�M���I���� ���LŏiO��m�gT���ҊK���.L�m���v�̂�a�v�&x�>}��xL�������z� ��s�.ӂ���@�S0�����H�`
ڗ7[���������'L�a�ώuz°+�=�q���AX���J_P�p��� j�ǎ����(�?���n�4�Y�)ӡ;�?�>�#V�@NR"�GF�~A��3����A^�8yR��[�k�c\A�R�iڹ�c0��\&�R�yY����y�J�Ĉ��ӵ�<��:S0��p�k��& 
!4��|�
�\��A��x���8�h���m-/��`�L���+5��S�l_<6����jː�0c"����4a���i*��k�S��m1�`��;���f�������c�a�'���2O9���Ҷz�'Θ��jyg\mN�gG4g,kG�j]H�6�;�&�T�I�����j��#����4������g�d�#4��+�e��ݜ��f�&���l�����
Z�վNOZ��!� ���d- ���&h�i	��}�Ź�:�nJ�B\�GE��<�gc�tSy)��UxHk��V�l�猤w�@Yp��x�&ms;�g���m�ص��$w��,�Rњ�G���
���x8q�� Ѷ�׼�Y    IEND�B`�PK   ���X�,Y�/  �/  /   images/6adb3134-3cc2-4380-b4ac-017fb4b87c19.png�/WЉPNG

   IHDR   d   O   �`�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  /5IDATx��}	|\�y��ν�o�H���-o��n�`��pC!@�@�&�mR�#�k�פ%�$MKפ�#!MHXfI �z�6�7Y��K����������ܹ�H�d�/�����f��9���;���3�t�S h��uj���c
(Ht,,�~���<��Q�P������2=�ay�A��A�<g�(r��d����P�2d�E�.�(<5�C�4����|���T�~��V�����n����&s�2=�a��U����:b򠡒�s��r|���h���C�7���A�{ԕ3#^I�ǺF1�C�����A�Y�Y-��L^`��T���:���F��_Z	*�C�E���k6���Bq����י ����/���%>����i4�c��s���U��7��h+r>�K׋n��p�BX)@,���;yq+���Hg�<�n u�e?�6�^���5� >����,u��p�u^�� ��ڇ��Ë���\�ƒEn��^���YB\��e>��ǧ�����āE��y�j�B�s��3���W�O�/7k����3�T\�����eT-��7V⹶Z�s��:�0���L�2�f[�H�.�$ԺGQ�M�ݣR&.�����^�HH��-6z�����7�ۣ)����t$T+hb�^�S�	���n���K�N�>�")8l�\
|t��G��ʅ�+�I#�͋)l�߭���qjK���`�W���}�S��l�51@��	��i�����{*�)�ת�I�l����.y¯Y+�} 	'Mfp4��
*��ڡ�qܾ�.�@N���i��r�Ց���!7^xa�!&.4Rt6��������.�~���zz^�Š��%��Ƹ0��D������#d�qn]$�}�����6����f`�k2-�K��ΞnB����Aj��]���Q{�ڿ�Ձ2�m��i��Ldm�VZݩ���j�32�"���t\��/��HLŚF/6�`�4�x��0�y	:CZ�y"t��ǚ/�\�;>[Y�����=�c�@Q��u3jk�\^��JOf��=�]�-�)�h��ĳ�������;��:\��'��M�Ѣ��XQ��ble��+�<1"�L��e�������p�3��'��oQ#يߟu>��!E��yE����w|e$c�B�mg�+��dN͒�v�m('yZUj��C�A��k8Elo��L��BȰZH1"'����r�,y��\	�i�LZ.	5�T�L�f�uI!��H�f����/o�x&>M���Q!�{���(��Ǻƍ{I*�@�<1Z�=1�=����p/�!��3u���J�0�ډ�h�Vy%�{��F���p	|n+>�Z��E[h���!�գ��r$�$�d���m� ���׽�h����bAs�	���6��v��{������;^"����5t��	����b
�:i�I4���
x����J��<������i�?��;!I�����>�%����N��ڒ�:Q�99͊�����-k��e���A�k)<p}#�yomC)Rh$��
�gD��Xq'Ό�kl.���Z��cQ6vvag��V�Ő'�{���k�_��´ߘC��"��'1t��p��Ⱥ�T_�^Y��|�W��e�Ǣ*D�|��x�6�i�D2���ru�N�E�'5���^��W�k!�H�h��<�L���AHn��$�z�l"�hUI��N�.Y��Ӎ����V�uA��}dU�>�}`s��j�8�\��ҫĈ��#=��ƍ_	�On[�t�]�s����t^���	�e�uRdU�0�g��VPmm	���c�'`w����b�+��o-�-7,Ɠ{{��o	���EV�v�hH�X(`��mVd,2��I:{�l)u&��M��4[Kv�,=K_�-䗴�i�N��,�un�Lm#�b\ED)"�����u�~\��xk:ۏ��$�g���&�0�9�s��N�/�@?Y}�t�@8�I�8b��J
"�g#�XN�M���>�����x!��ݎ�=�|�H �A�f�H��A��"���k���+������B
<Nbkۺ �deu'/�CX|��a8��nzjz�e-�/�Չ�CJ98���Z���-�|���6��G�_��<�a��'P�\A(Cc�*�������jb�h�W�-�N�%!?D!�ף��z��y���7��&jMm=��T�{:ҡ���Ǆo�jo-���	���D�b��YV�X4��>���\W�ܴ��*�_I�Ej��ھ"b�$���7�暏!��k�*�5/��3����[s[v_N��B����I�Id�8I9V�c	��=$�di���Ǫ2"�ڊ5��vG�Cf	���BC.����Q
j�#]9��_�E��G��2�4�UKJD��XOLx��	P��uc�D�|v��/��>�1����q-M�-�s�7��C�$5f�u�V�g.~����&�$[<��mG�����j�9�S.g�?��D�	�;5*&vY6�J���V�n�zF8���޿��)�!�q$�K+E8���'���D�2TBcdT�����E�0���k��9d����1��ǭ�����s�6�땅v^����g���h�c���;���O	��ƼA�ӍkKQ�ds�8�G棓�1&^e��곃| �%O�N�D���8�jӲ-6���C��>��[o�J�����4��t�|V�le]��}��"�J�8|���'��Lv�91Lĺ��Z�9�ڲ��)�S�Wa�d<m�#�W�w���#?iC:�������J�����و����>Χ�doߔM�q��v,Ƴz�xﴦ$�%k�@K;�C:]���v
��V�3�`��N����J��G䙓�H�Q\��8d��F�%^�%��{�C��M~�_��'3�`οO�Cd�b;~:��Ѫ�����M)�s�a�*���<�")�#9ǀ��Y0?S9�ы�������A&e�P~�M��@��A�|�HTM����$�18��-R�.�n���� [[���n�
B���a �m���>LC�%���2l6Yp�B��Pꬷ�6|`]}��'��`8��sɸ��:,i�t�xq8r� �e���!Y�P�cgd�l��}�}�����2.�#�^=4<��Hً����M����ںb��pJH���I#���綻�;�#��ԟ��@���%����x{��g*z����M_c�4h�I30�т,/^�5;���/,�"���~6��l�	-��B��5rL�J�D����:)n�90��J�D0��lXn��������Aޒ���,%�e��z0��m�,S����V�@�*��'�'DD�0'-",mRŰ%��D�;A"���ܚu�*R҅g�݃��~�lK��}�;�W��m"��-�E'�}���Cᴷ�'���Zp�{E
W�b�\	.�y�?5�a)�(���`B 1�m�S�j��t^>�Rr��5i�J7���|H�܉[7���K"@�/;��"�%��@�E�֚>\Q�O�gӗ\�A���Kv���BC&�Ʀ�d%��:O�l!??9�m��7V��3�ʩ��}�}߿������ud���d�ׁk����`EN�O%����ӗ�T��ڵ�ca�!,p�\�&9s)������Ȍ��"�`�DE�S�U� ��h��t���&���	ǅ��dg뇿���Y�t����"����3T����Yl~]��M_x[�{�T�vE���$�٢[�Ȥ��[�r�
��,����J���#4�r�u�(�t�Dׁ!2@,l`
�躹����z���v�`�X�~=Vմ���������-5x�Ȍ�?$�%��8.;��ce�ԣ�uS,k�����r��v8H�u�9�D~��j�>�ֈ�!�e�A��jc?D��]{��j�c!C��%Z�jjD��;3c�	G;=WCV��%��x��Ql�<�;���ڎ����`��pIipA5��KJJ��T�Yܺ��$��DF�U�?d8���h�t��w�oO7.)��Hځ�/��.Î�
���A�"��g����:��e�
�a��������ۖ�"�ꃣR�=�v� �X``�-�G^�ں���D)F2[D�0�# ���%���$\�q�_Մu���ʇe����[C"Ž y����z�w�	��}�m-V��#ͦlL?Ă��ƭ�����\��Ǣb�9i������΃��Ø��"D2�q��JO���+�+,63�6$
Ks�����Qt���}oY0?$K��g?�Y���y�Jz�zV��W�pʇ�����>llrbe�5�0.kP�b����gT�%����� ��Se��C�L��n���0�lJ�jbͷS��dx�&���&��/xr����'^�i���@���B����.��92N�>����&��i7oj"NrL�;q��3~����Cp�,��G!A���++��Ή/|�(\J���f�u����M�۟���^�LJM �)��-�-8v�<AUU�������i�Fq�h
yjL�xa߈���ɸz�k�]�,q{K���'V�B����O�ˋG9|I��@$��=|������V�e���9���P���2�k3���S6\߰Ϟ�g[kң5�+Mr_"���Q���<Q��c��M���j=�w��R)d�Y�=��#�Z�1��_}/���t�A�'^&�R^Ȥ��3v��Ջ�c�>te3�T�@n:{R�D��ٝSV�B/�_�74�a�˫gS꼊�\GM��%ĒFH�;��_)u�ȞϽE߽TO�����ؾ�B���ؼ�T����<Z�c��J��S��,�k^�;�iY�������t(M��K���<I3r�����
�5���x����![F�3�X\6����G�	���m}�wߔ��n]2�lHCx[X]��Z��E�sG3Н���*4��K��j�`"er���,�B�1��������S����x��1�pvk��Dސ�WB�}�ˈ ^����x��xfsNϊr�7�{����2���YlɎR�o+u�roF�>l5e:.	�`Y�*r�\�l��so����=�9M�39�7��E�g���
Sav�bE�E$V���*^m��m���J���HP,g�=�G���m��F��6QEy�Dےj7Ҵ������.jg����BcťX����jrH�h)U�i������bH���H7���cW����rko�@�G�Ϭj.=l��J�'B��}8��n��>�Й�����-A�(�ߊ�X �JŮ�ʄߠi3�"�1�����f�|����NS(aG��&�'2xv�0�ݶ�4z�zZ�%"���jq�0�cIr �8��7.�(��
"_�x��g��R����v�ڛ��na�����w~��`=�,΍�;�NASLO�߉x��?��fE��T�#�7��N�W��_�=+�����*�����*v�9W3C�f�6�iM# ;[,�/��G��s�e�+p�}GF%�Nv��w��z|��A���I���ֈ�t�c^=l��{�kă
���Fh+X����S�`fV�d�㜚��X�D|\�."�y�9���d���ϩE&oan�Q����{�����S���}��^z�L�WX"_�ܽu�t�9żGM��w�𥻖�U(�E�Ǉ!�
r�8(f���-��
�X?�n��U�8%,�������C)�{4����/���Z~�j��Q���(rv����6]��l�F?Zj"����_��Z������ ��(�[�������؊�hNG).�S���MM����x���*�c @DY�H�x�R��M��{�BFȞ�(X�B�X�bR�LF\����S����2}Q?����V2-��_���K\"b�~��zGT�92��(Y����E�!{l>��Ӈ�mQU�2���N�f��]�^��>��ݍ
�8�eE����!ʄbYo��ؘ�V�yē,�����%%n{NTM��2�*oi��j��𤘫
��7wT!���{�rf�JC&c_�5�e\T����Z%|� x,�q��tU�����X�ձ�/������~�Gw�d������O�¶��Īz���`E�zi��Wgs�����yi!��Jww�8�zy�i�h[&���ŚN�(w�pw�q�F�S���Kq�'����ޫx�x��A8��?ӄe��xj�،cbX��� n^��[�H�l�����v|��2A��ye�P��	E�r?������Z��K&�\(��K��pb��
�v�c�R���A�Y�3)�e�O�e$�8s��K�Ê�X$����}	���)��[�N�
�v�o��%G��|$A���z�O�>R�ű��c|f{�^V��/��x_�A҄d��NB�>&��V�Wo/��51.��̅�TҪ��L��N�'�y��PN�9�\ʅr�~�?o����z|y�[��D��v?��zF���!���n�!�{Ƀ��&T�J��7��fˇ�ZɊL�;V���.)���g.-s%��?��}��.���	:�b�����:Jp�;��uN:��r�o��=[�ב�����9�i�o`�j�ì��d򂸋�r�����Q�yE$��3
r��85'�C:ēy��������!�[�!C�t_./
�3�A���EBپ~hX�����!�dNA&�H�Eo�4O�Y۔0y��K�e�&�F�S��cY;w��w��ϟ�C����m9�]2�Sy��A\�܃�yr �i8�2"�}ê'�Be�R"���sL���D	�xƆo������h;��qr����"%��]��l/!������O_�蠭'n�0�#��f�Q�(9�ϝi�v.��EᇤKo�W��)��&cvQ\�kID�EE�+��ph0��%N|�*�n��h[�y�����c�صe�i����W?��fnXyq�1��>%�r����q_�́�c�<A2���a�P��;���Q�g�5�ZW�2�E�w����^̖���0�	�Ϟn&á[k�џp��c$�-SB��_�l"�a�q�{�o������{k���|�t��C,���R��	�i�������p!��v��L��i"����d���|�� ����)��}ĉX{��}	qp ���Pp$:�-�&	#��{ƅ���q�qUi�J��9�|t[)���<�HQn\���L�K��x�l�b�u��[�����3�M�^|�b2�i�z���_��-�x���:D�S�9Qpl���?YX2����˖�R\xQ���Yq����5�v��q� ��1�2��1<u`�V�����7����MBBr���=�!g���D����i�._ST]���&q�[/X�g�5A�֗�zp�յHfe�:bp+�9�w��d��b�}���O����/mq���Ů(9yYrm�~�K�<�!s0�U��MQ���c��q�]Ǯ��0����b$Aʝ���OƱ��{O��d31�nd�Ƈa����/��ݶ�Y
~�C� �6T�"����[[^�ǒ�>��"]�`r���O�W��7L�%+V����������h';$'aE�1"�/�n�7���(��q/9PY4֖������y����xdo��S_�dׅ�	X���ɽ�s��L�Ny!z|��|D���(�]f�@r֐w�mXĻ�F0=�Qt��az�R�s|z���ȘW�Ʊ��MX.���FB��|�P���%3b�HK��􃭽��,|>���J��:��c�"�#Xj���J��(�,�,U%��u�7;E� �,��U͈FGG���Qeγ455���Q s&��w9/3W��$��;;;1222Q���܌����K�GIdG6f&��z;�[�*�ļ�[���6��+O"��"$�&�(��1Xy�K8��j������%�VE�&*�xTE�V�XҐMO�\;��?�b��HLf�sr����b00�9L�Ç���;v�@MMf:ab.�����8�~�m�����f�|ppP<��ݹs�xΔ���M�R|�Bq*hY�7��u+$�t�9���A�D���$lh�������*�J���[ODF�p��	*q��5��I9�Y���a�WY�p��. R���2	ŉ0����m��&��{�����o�!����	�O�09�����>��nq�|B0S�,������QR��Q7F�Q8%38l�X�ɤ'��9r�!*��WU%��GCy�Ű��P�NTO����s���0::*��!���Մ������ݻ�я~T��� ��8v옰��.�Kp�	���ؘYCCCx��q����gf�"¥�v��6`��(R�QÖ�p҉�|%�6�=k��~d,18�pQd�gs�99TU�57\G�%!���z�*t�Ec��evQ �Dpz���_��=�KtS�I���F:#���{�왅�=La~��D����7�pN��:�m�)������\XYY)�Kkk��xQ�F�A�b9#qǈ1��)b#S���w�-��>*�����D�/�u�6�*��O|I�2v$,��^�����TJ��q�	��[M�<�&s�+;��!���&�y�+JP�"��e�*%���x�<a�NWΦ����A���
1âm.�!bu�#�pӭ����g\��DiooǺu�mZ��(��Y݉=���^H��N!��H��ߌ'c�#c݇�3:������[���*���5��b�M$��O_?�3*���(S�՝#��'W5ͩ�GE�1��,�z����(� ��2�*�i��e�s�����g�p]B�a�p~�8�|����cNai.�0!��뗘Qc����'��Aj�E��\��4 _�{�1���N�|k�4$`#��Z�5��I�X���(��O�#�,Ɩ/^<������p�y���#80�Geun���8ъ�`�5Ib�ee#��@'��&kN;3�ӯ���s�t3v._�X���3��m$5��&��$��l�>�x7`4�8{�{�7%���S$�y�U�,����!
2����H���S��:+�+������DVހ��͚U	��,Y���^;�o������@A�g�`�^T�2��&��(�I�}�Xb#a��{6���'���|�a.w ��W��;!���;����Yw6A�:zi�V���62A-R��q6�j��X� ���24�}�����h1V��g$N�Ԃ��a�x���_%M޴Ӎ{��˅�6�;i�
5����j"���Z�\J�	���Ik��%K��U����Q4�K�I��L�ˌr��%���bM�$�|���YX5f��R �8(Fꖏ�\R�)��YK"�ϑ�v��<��"m�Y����8~R�H�Z(c�VY�&{�6����2�R�5S�AF(�l�B�	�LW��3�Ȟ�|���"��M�Uf4`6���g����~�3���
�\뼱�#HC�K�g#k���e� -|�-��9�˹>{�Ӻ~��}�fE��C'�|�oj�[2I���F~���B��K+�7�)RqF6��ʕ+��?���y��1_����go������9�L�s�Ԙ�1 "$s1V�ꏋt-���%���b.
8D�)���IU[���,"�Ń�m$sǩy��bFy���V,m�b��Z���Xy��VH�&uCw�kB���_-�3L0�OCfoڴI8p�!�	���"r>�&��_���l�.�<6u-ZtVl�xөQd5�q�<9D�8��K<�8����UXM=�)rx4Qt%�O~�k�Ӂek��U�I�)B��"6�+�-�AzW2��ۥ��WU����cN����.�8<� ��á
5y`�}.OP(I�G]!�������Hd��?�`�^`�����糷>��B��F�=+�X�$N�qf�??����C��cO�H�*�4�q�Հ��;�U�L�E�n���5��(c�J\�m$2���ACBw^��@�(��|�|^8����'���s�7�������D��Spxk�8	�eS�����,�|�?��Qt�8I�O"�E̉�lF�y�>/���oX���?\@g���F����a�U��JT���o�%�uu!.w��S�2g�P�.���@*�an%����'vW��KC�E������PF^EC�~k����Y����9#���qĆ�!/90�mB�|)B�d�X��#�|�S����18�4rEAG�������*%�#z�8�#����1���%xב��=2��K��������dR���JyĨ�י��9�MLC����CGDA��A/C���8A�,�gaS�q:�8�3-���ڭ6d��W�XYU���|67I�퉐��dq���1"Lu������*X]���~����o��_�����s~^r�3^��N��L}rG�l�WjA-:��j߅q��� *e�|��$KU!Rl9�t�DU���i(�2R���5��aKs%*�;�>T�C*�3����K��<H�7�&y�i�10A���?���ש�,�������a	Q�C�9ƥ&B\館�`�sx���Oy��B[�	%�$�G�pr`��ehZ܄)����8ׯ��W�yd�k�y�Ζ�3��&�M�_�q���$���^���q����l�E_܎�ֈ|y���q�ςO�����5���~7~��f��&4�;����y	�Mv℩1���*&�3����9�o�)*P��qĳ2F�V��8��K!?I\M�3��eYQ���2}�	�I�/�~��	�	�1�j�.L�"�p
�kX�I�R��%s_�!�5ij�؈��'1�r�"�1p��d����N���n�v=e�8������ZU,���赛^�i�N�!���J�Τ���-#θ
%\�"�lwp�i���Y�01�Bvq��"��8�X|}z����`.n�N��(���Y'��z�84��Z�	��<��)��2"F
�����MH�z�IT��u��R��Y�.���Ru6Hs�"r�3�|{ɜ�e�)��!w�`���p<(p��ӻ"1Oc� !�๙��8�L���1�����5o�	��C�{b�L3�a����	�z�$���CZ6_�΄/����%c��@�r`�Z���ԑ�eU����շf�J��7��.���56���BK�����	�H�ˁ�؍���)��ɹLr
sG�kkk�9�?�sRD쁺l�;���3���H�SG�(�H���D/��|��\)�G���z�5�����V����1��G��i�5D�s���F@ҋ(�H���C;ӀW/#�+G8��D&�""-���2��b��s.���@����o�'%��ಖY��ӟ���wS��Ǩu�8P�RB����P��J�����t>1b�d��c>�x�pJ󾑔��cnh���d���y�{f>�kD��'b���JE�s&��Ñ	)��N������D�\D�:/i�x\�u��A������,��	�E��|#/�G^����z�̞l�	p���S�T�%�/�ǣ�wl%.�@�9���/;����?;��)��%�
�*�}ٕ,��A�v�}7)����T.��2$�鐊G��1�ߋ-�QT����U�F�|,#3���2�_�bz�m'�>Ŷժ����:����1���(�ܗDy�M,��yF4�(.��l�s��s#=�S���G���N~��e<��,��M�wb�p���77"���R���A.�L���p�L{O��Lp�9�#a֕�b}0�jW�č.cw�&jt��׆Y�2lV�w�9'��j�K����4�ޟ���Rb�Ԧ&��ٌ������W�ɝ���>>c�O�}�	¾�vj�^fDZ�9��Z��}3�?��?z��G"M$���H�KV#��R���;C�y�XQC�/�z+��۔s!�To^�&z:��dX����q7]��.�?������h����(��u�w���"S�9��� �"ǿS��O    IEND�B`�PK   ���X
=)�.� � /   images/770fe9cc-a3ef-41fb-abe5-14f6fd7b0eeb.pngT{T��������	$w�0�]$@��n�e����u ��9���^��tW���I��h5yTRT  ��� �  , ��Ȉ�o0ϑ����ݤ�����e�3
PA� ��z9az�4�_����s�t�v�}��@ N;g73�����S1R ��(�Z�+�x䥥��xv�jw �FF�pG�x��Yo�=��tBv?d��1�JF�2�17��"?"�`�>����I큥���Q���?��#�k����=_�:��=R5�cb��ҩ���4�c�
aa��h@��w���G�=�V'�wr؝�j����i�ᰅ �����7�J{�r��A�_ڸ�b��S]c�'��.`�A���=�qȨi����1�%�>��ck�.�cȇ޾�O#��̶�����]�U��o���6�T�����_4[�w3ļ�QHG�~I�o{���K�Q�P �����/8���Xf�8�iV��(L�����ɤ�G�u��O���>iy��׊���jc��� �����0EU���-|(���B(z�z�����E���#�1xF:��/�e����j�M=��������^��@_��|�M���>��.�g��Rs^�w`�rH��f�6��|����+PKLA�������S��l����aR���-�65晼�L���f�R����|�{����:%��Pu�����p���6D���#y���6k6b���9��&^X�Ӗ2�?s���8���ğ��J��諃�{�C���a��|(�mmc�k�A"��Oٰ�����=�+&�q;2�{ͣ�7���l/����.�����������㴯}�R�́���x�bv��4ď��>��N�S��� es2ӥ�<�l���"�l���.<0~��[��~h�b��ֻHɾ?���]U���S~ �[+�/��<�z#�%{1?�֦gw�> y9�K�7"|a���\�}()/�5F�m���.�=��h��O�?��(yk�;>��N�X�!�� ��#
6�M$�H�$����yl�8УT5ڢ�ϳ~���j�������7V�u��$�� F$�Y�31��Q%b]~_��6~v1ɤ������6�Ӿ�˻��s/]d���XE�?	F �2��:���|�}[K�=���oJ��3J�a�l�Ș�Z��
1R�2 ��9p��oF/D���$�LO�^r��&[p�'������N|���q��y�ъ��lf!�z{���a�G4�a_-r�On�|�pp�iή=7�x�_r��8�X�yj.U��h�Ĉ��-9��;�4�\k�2AUs�;<z��e�cQ��$�K���[�B=S'L�b=
M��X�A�y�U���_3���~~y�ण6�դ2�, S��.�$�5?�:͚9.,��s�U�Q�~D���CJ�w�ɝ)*�������Z�����	���-RL����W/���Y2�o�4���}}�y����|��N��t��ZpNe��C{�6<I��	�qgʝs�4!�K*Њ�iS뛉�c�LO���/��n3�4D�"��ഺAd=�^4�[\B�|f
�@���B�%�� ���iDv��w/Mn��N���K��锉VRԽf�� ,x�(��'�kvh���+�=������y�6,�s��ّ�@X�T�h��czmƘ|̸��~i��DO��m��:��ھ�d��Y��%�_�=O���_��t���=�@��P�O���ѥ�������9vi�z)�al������=�|C�)!G'�����tOe����i!{ok�th��7u�ոMU�=~o����m�J�C����^qC_�f�5�ڣ�@�]ߋ�}e��ش��*��M�#ɅS���I4c� К^�q5�V+#�U��'��|�6&�w�J	c~je=�����&�_�6��c�^�}y��m	����7NN��/8c����1�O<�?MF�z}#�"����f`����6�OM�V��3��R�`�xؑ�"ꛦl{��t_�;�,����⊏�(���
���ק+I�?��������hQQ���O�����ͅ������]�x���q?�z�6~�R�P<����]� ��+�P�Ѡi��%�D�RQ�o��w��"�Uw����C�|^��B�������(odD���y�~�͈���%&��Onzn�Ǿ>��G�O�
7�爽�]QDK�oQLl�H�����fm���B�f�׾%��|^�������}��;Qa(hiiI- @�c�R�G�l�C�_�����WVbz��[�E�܏)1�6��0���4���>�f���yD+N/'+/����<$�q����ѽhsg�a"{`�fbbbP�tt���7��Ƥ��V*�F���Ê�+�[��2%n@B\�N����ѧ�L��(@�ʊ���<h���(.#Ks"+y��.�Z���s|á�h爞~%�p���c��@��(��qWX}	.��K���gd�ecC[i������]^%��EM�l�a�⒇�)�k�_�w-޹�{>�]�DsM���[q�q�[����XD��8WW���<���`�o"4�����9�Dx8��S����ll�wG�$�s_��58L�\Qf��<��K�O��+.f�/*��>�67�e'�]-�Q's��~glL��ʪ��~w�����|j\�^��Ϥ��F�o���=��ї.�F��x]�¼@��7T�78�Jїdg��(�ô���.-,�8!�pAEEU�-o�O�5K��Y��a�Y�2���0Zep��̪W����3����p9��Dh��	Vb��D@����O��;�ZX����!Z�ɝϟ%�/�� �Bї�!�`�2A��d�}�D7�Lgw�b��]`NeW�L�QR�t��|3����g�{�>;
�BS�">���"gJ��z�q��H%�`�C�F哐HΧ���zϋ� }�1E)���J�=5y�5�\��{PNCW4����\�fZY����?��>� �!�#Q�~�PP&��2Q9�S�-�Iٗ>���>��j�����i�?q��s�s<�EE��'hHe��� �c�#S�����?�6�
/d�:��S8��1 �
��%��'�On3B5�$���]L�䯕���{�4�F���Yn\�iɵ0O7�c����\�t����/c1^���A�%,/�K�4܎��=*G��p�4~��C�Q�6�0�.���ٛ����0�.�ui�S���v.�Ikz�|� �;$��(��nǟ�^>}���X��]Q������r���v[� �>b��cQ�R�DC��oPM��_f�Ǧp����<�ޜ�{D(�����d�A��in�7�����)�"�{�85�[p��B�ŋ|1�]��aY2����
��r��������'����j)���� ˀ��Y��:��s�$�F�� ߙ0�f�w�Q�?vL�B�LI"T�H�"^�q
��W��S�8�6Գ�׿�_�H��=	���S�T���/�~<[,��h�Q��XFܯIb��k��:O�Wu;͞�e#T��ߤ�;�.�ʷ�\��QD1?W��a�)�G��*���Դ���	
C>�:��q�(]@�����;�~!A�����. y�.���<�"q�_�_/�n&'����>H��k[k�/@f��fD�K2�u�d�3UD�+,f�'�����l�J<�g���4^��%�+P��e���̩_L��\[��1]��TΏ�"��@}���n��J�1To�����c/w�K��_�i���_��<jr?��3��_��U����ekj�DQ 9�뙿�<�R6��'
U�V�;��g���hB983A��&���uZ �H��n���<x���ݔ�u��TK����>\�������>�XE9?b��oA5���K��?��/-�x�>�܏�@�FIz�9��?-v����ǃ��^�]��t!z�o�u.�F����v����f	0P	�!lk�W�P��	"nh��O
H��ACU��ydL��}�~���6���-d��ᯇ���缯n^]�U����&��{���;�E����	�@&��)�M�F�օK$S�Og��6�`�̜�*ɁzEA迏����$FrM�z��:G\~���݃ӄ�.�0�[�/gY(����>�hN�P�@�uYP��	��M���5Iy���'�As����oig���.��O��ɣ��F�u�����áUJf��RǒF�T���X	�����@妽͋�=��Y�����ĕ�H��Nli1s"�%��=��[L,H��u|+��J ��{Q�|f~ί*I�H��R2���(v�����-~�C7;;�_�;�(PK,���unh��ȇ��&h�R��뒎�$���Nn��F�/�~S��̱��~<K��N����W��r�;�ЛC��8sY�/�jMɋ��՛�i;��ɮ�.���0~JV��n��x����*��(.+��䊫R�}�1]L`Z�$�p�&7ᖶ:���G|����ٟ{�'�珯A��}|�{|�o�!NË>�ί�>��'�W#�fPTUss�!��ٺ��9�M�o5 �>a?�ٽ谿�2g�s�*��4Q�վ
�M����Z�N"�ݚ��_������a���;9"N��6~��颚g����_��P~����B��E��c�UTA��0{ۄޑp���>���H8�~(�;�4�F�ǌ#`P���}Oڶ��tT���ډǨc�~`y3Q��!�K�޼r�#�8�하�޴����T�}��̘Yhw�մ�����`��ڴ>�MҀ�.cIJ�s˂�zv��Sw�X?23��B�l�>)}�B[�x2��syB�j�qI\�yD�	-����o*��������f��%JCw�8�D�.���eK��8(�/?�p`.=�����PYu�	b����j��]�^��}��񂌽ޟ�̈�9J4֢��sf�N�_fW��ٔ%�>�C?$�]欙7R�RSZ���`|'V[+ZH�K;�������ţ[�v?��@�t ����&�u�Y�JhҔ������b�gѡP#���VD�X"�N���n��s~p�`���42�<X�p��	���]�vaq�����o�^L��sX� ��:8k�ݗ\NN�rѿ����o�Ym�^�l�0%;_8��:�Ā�ܞcZ[���J��7��R�?���X��m/���4�گC���w)o���n�}k#֭�z̮%���m��ء���1���+�ޟ��`�ʎ2#wb���垻��X�|L ˅}9^i9戏U�a���F����"�ǝ�X���Ó��
�+[D	u6j��ӕ+�T����o�	L�q
��<���+��H#�o��y"���-�S��H}�g�$2���A-���Q�7K���<˻:�}����x�-�ϛ���^�����}��UN
(?bPF��*�/SՇަ��T	��XE���MQ�!����h��v�r�f��?�W햟�-#K�%k�ܰ�+Ej�-�"�]��������λ���%FY���W܏��o4���o���35��x��Te���ν�S��ua)�'d.���+�͔��������rh��d!d�)�O=!FD;`?~��#�e�R	N,|Bα�J��DQX�G�FC��� �ތ�5Zc��T��K�Lx8�P�ӌ��ΫD������f2��P�?����Ҋ�~!�]9�P����2�K�/���@�kY�.��᪐�����_I3r��ɛQ}��&*��Tbo����,��@��������7a���B|�wC�߱`S}�BZJp���V�Y�N��7c�Y�J�2����+���fQ���,�q,v�j��L'�-f�Dm|*��T^Bo�Coc�hQ%dn����E!J /w�v���A`2���4�%1������	�ge�a`���ò�י�b��*~"y�s�4(��$A���-3V��¦�P�q吣� :����Àt��U��W�?����D1f���e}x8Gb�5���e��.�q������=z���~>N�=�X�6�� d57`���غPZ�_[�\�7���:'��K��;ڡ$��#���z~���Y�*�Z�|����w��2*Q�7��a�����;@}8O���H���F�ڥ{�{��v�RA��qmS�j�!{��Q��q���3���� 	U�)�54r���d�\��-��ꀓ��*�;Ҙ6R%F�Æ3�i�$̍"�	 S\Fn��dӑF�F�{�Ɏ�(�{��U�BD�Q $�8"9�w��r"g=��3�F�'\a�v�M�μ^a�cS�Q�.�-R�̆i�����*zU\�p�o̞CH��e�l������.d�с���:�^�����JRR������8��	�'���ټ�kʭ��bp��O��������Jш�Ո<������N�g��_x��I�k�϶���xY��M�Z�|���Qz|�S��W$� ��f��)J�eNk���T�q�����C�im��� J�0��΋�C��E{�[|{�:��Xvx�;�_��
�D����+Q��d�b������s�5Ga��*
��#$�J�w-N��Rz"�{��l���6*M���Y����W�ދ}�z�k/���� j����u��l͝�%#Υ���~ĚcM�o���9�0K�w�{��_c�j�D�.��3���XG�!��:J�{�ɠp�ӛ�e���mEC%�6ܵ���M�u��aJ�� Ow��Ӿ^y!�(4`��r�"�U<�i�̯X��0b�n��A�-jɽڀ���������,~PU�v���-���&o66���B���@hm��t<���\��^a��i鬣 	���@k�:�or~T:]�P.s��}�g!�����O<���h�,K��C�ؐ��� ӆ�a�҈'���ud͇�@
l�ⷰj�m��P5������֋�=�ʈ��6�P�����q�?�e�����Kj��LP(�k���[�$��.��x�s]3����h\�a dIt�h �<2)&��T#oq1��L�� ?�8�)��fW����Z�q9�]�2s]SV�ly"�!�����Q-Rx�:�r�\H�d�-Ze�&��h;_R������Kxo/S��SѾ���/�9%s_'=�Mw@FK�˟�x��vEg����σ59�����v���"t���-�)+'P[���5���>f
Ԏ=����Ol=�'^��Y��q�~T���y����T(���/��u��H}筍��,�lP ��^�l�DC��h�H�x�Ɠvy;�����[ �����a����<a(ڄ�(;"�"Q��Xn���ޓ��rV�7]:�UY	��o�����]m-������٭f����۶�m TO`�E�vq��)��\|�{Y��2*v���w�0U�p[�N�1�����Uw���AW��6�+�����7�0�����xzb;�R�z� aj.U��p@{g��������7dPP��cfH��S�cx��Dh�惬x\�{�\�es�ܺ���V_^� )�AG]��NVE���O��c2�"ʧWoy<��N_M�*���J����J̥.Y���dJ,�)�b�<Y��jP`@�w�N��j5�9�,eղ`���?$;a�����r쮴M�n����6�t/-nLc	f�D�z#�T�&�������r}%�� �ŚC��Pv�t����n pmI�t
5�];&Hv�"T����q�^C��Jo��J��0���6`B<�nE2 �V��ul1t�i+ �^���}qzs�1�7I��U�%B��	\r�XTv�Ͱ3,7-��K�f��T��,��UpM#��@\�kkw��B
8��#�Rw�&�qV�ٷ(�A� |M���v�w��f�QX��a��%��� �ȝXZAH�(��D�GAoS�u1$���Q�b��/g��sK�Dud%VӇ齟����t�w��1Pw@R"�6�]�P!)-Y��[ɭC����]>���ͥ�����8k��1�LG��q���L�8j^1��G�u/z�<�TJ~�(�C��/�4l,�E��B�o.Y)ŗ���y��]Z�Ł����e.���tE�����F�&�����Wg�ۆ�Q6��|e}�Sh��zh�xX*ͷ��XQ�ߠ�,��!������%J�{vaF���&<��9pa��K�`4D�ͷ�M Ӵ�mQD�/z��R����=��-ʨo��s�Q,e�h�Z5[w,@ް�����v*�"WJֽ<�&�]�,�țZ��T��C"#��`Mf&��u�&P^N �{%[c��ϫW��&	pY+��T30�&�xf�p��P���M1������.�)+l�hh��5ۻN�Qc-�U��'����K��xr�j7���=ˢ��o���}NU��?���j������X��0��ĽY�Ü�l��fqp�8lt����UZ���17f�|>aq�4m�E-+%�v�â�r�q;����7�o���cE6����W��`���#�Sח����&��6���փ*!5�X��ښ��[���酺Љtd�*ڴ`7��ž�|]~�礢���Xԍx���b������8Í�ˡ�Sk����X�\B�\���)s���C�s�<a��x �����kcש��׈�$�e����E�y��u�5;KCg+�[0�\�J��.����y ���T #���F��Ǐ E��� �(@u��uWK� Zv+���V���q =ӳ�w˧W�o��򫮈�t�kB��?0�8�ן��E�iŶx�-�A 4ɳϏ�S�]�t�Դ�|�r�&�C��֖K�au+-��X�C>���mMJ��ˀ��鱞B���$},Z�������P6�=��e2��k+C�%<�*<O)埐�j�捵b��x���m��M�S��ڿs^ܾy�J/�}����>����d3��ؚ"9.�q�-d'��8e�pr���������)`u"�뛼0ܕp�{������	}�ޚ�1�vǩ<�2��<�+�X6�2����U���>�ei�8�G�?zԍ����<m������&� $�i%��N�4�<
�uX�(�2�(���)Q�,Yņ�y�*��]�G�p�!�`޻������,am}��q�垑W�Y)�_�,� I"bO�&~չ[UK�����V�(���27�"�1g��V�2���c��)9A��M=Ҽ��!���;�j��3� -�R��Ε��e��'���V� �?m���%��G���O��<�:�hi�<b˺Wdg[�tX�rp�,��2Ϡ��K >��ȫ �d�y.��]�����pT�� ����n_̢��T�����J���������Z5�$Z]�S]�z��w��n<R�L/���A�04�� �������k{w"�%�'��b�B@������g�Q�f+.��L��v6���Dr�Ro��U
z�5 �$��C�t?���x�@y��sIw�B��f|���XK&B~[���$�������'t��2���Ǌoo�;o^gg��"�����0I8���J�i��u(m�L�_��5_]��q���W���J	�"x��x��HU U��^�:On�}������{ns!}�A\"�O׾�q�¡�.O�̟T�|$�u�)�0�>zMǕ�q��4�ҏ�ۜ޴O���
{��"b_���n�v����dāq���c�e+�������柵{��%bC��3xҧ�n���I��+�ݻu3H<%�C��H=r쏈��mH��{[y��j�x�M;Nʔ�:Q���5��	_h��ʟ'�7�P�_T�bC����߹�1RS��{�����''�t�"��Ϯ�A0�na���E��D�ouN/�q�^56�Sw��S��E�U��Pc�h�ki�����N��Iݛ	-2�
�_5?@���?�{R'� �3�
��>�x��4K����s�>3pĂ&\�J,����ٓf�]i ����qi�o`/[_���*�e� ��-!��52S�|��*tx۫�-���f,t2� �Ǎn���Z��0Z����b��٫j���W�#��K�FS�̇A�ڇ(�Cٜ�T���Gø��e��~V�P��*R
T��g� U����+_:	�z�QS�/�$n�e�]]�D���-{�A|(��Zʠ��/pF���S�![��Q4�l�M��7�1�z7����q�{*�V�Xܓ�5���M������������3��:��<)~/H��byX�$�5���"��g������>ڗ�e? �Ӟ�^U> 6�[��O]��ߡ���Z�J�g�p`u�jQ�.K�{F��t
w����u��`i�9D�Jʜ�Y7�u�Q�^�.^Ig*�1���=ZQ*�")��h#۽2�(T����@��A�~w�+.������JrG�h8���)FH�5��CH�?�r������2t�:4���0���7EFE-c�ґ��vc~+|�L;/������&󍎈�ޱq
	T�.N�E�]���y�W�S
�ڂ]�������]�i���2%{kde�Ν�;�:���ޠl���<<���Nq���7�^4�Bw ���{ kN��7�qg����ƾո��ߌ4z�@iOE�@��1�k�S�3�#�q.���]���*���1�Ahpk"j���Z���ee��a^��s1�2���鰜����!nr�ׅQ��pc�2T��e**� ٨5AT���SX�B���j��'@>w�2:+�dzE��7��s#�I@!�+���Z�����������S��JK�m\������S��#P�j�����x&6nCG
[$�8�H�P�1qSYZqS@�1�~���ˬ�#$��Ʊ���cE��bƨ�^E���eYKq���N�s$R������o�|^�:Х*g�杻|m�>��.L����Iλ����(mOw��*�H�O��gt->ݱ %eIG�.�/ ���!�ɑ�
Ul2��Q���ܙ��LX�2�����ᇾ�O8���0����o�.��:8ܙ �w�i%�E�
�w�e��Z����������Zr+($��b�h����m]UWs#��N�+�C�+@��[�õ��E����3<�	�&Z���[;�W܁&�ۻQ|�,я�`�~
�F{6���d����O�B��A��(Qy�Wp��9��|���D6nʻ̄�4%vu�ռ#3tQBq�jp����e�N {���=7D��@,X�Q� ��ڇn�Ǜ}�V=�,t=�W���\P��~��Ts���������k)��e���u��r�D���$gw�l����(<-?["O�2!��c��k���1�M�B~^�OJ�y,��t�p�pռf��~'G��e<��~��.���ڡ7����\�u�}��DW�d�}B���PH�c��BC\k������?[om僻�Y1����7P� m��b��e��N���0��z�L�*aJ/c	咱V�qdFG*m2��-�,n��,+��z�8X�A�6��<��n�~��ϓxh�(�.25q}Z$�<X�a10��U���'�R��]�l��!9t�{��։ա����
����Դ�z�N9�i�j�j;����4N��|����e����ڸ��q3�l?�� M� �T��k�l���doa?����tU(���,Ͼ�j�,㞍x�k%^����Rt�������~'(��v�\�\o�8y�n�VN�Y�Cբ�S�2l@"�y����� �(T�D�݊�c��a�UzU�ɮ�B����J_$�?�а�b�]pF�Ȁs��X]��.bj�A�� �S�T��d��:���//5�n4	�/��j�4�[p��#����n�J�N��v(�'��q���S��й�u��-�@�[����%g�K��J����g�,�L^��ڡ3��@ֹ��N�)�\�@C#��c>��#���Dr�����P1f����/}���b�7� ��!g�W#��F�0b��2z��1��ڞ��z+r�1r�z1���¯��y��r�٭[
f��>�Zx� W���A�;ה�i!4��v��1a�zI3����{N����A4*ʄ*J��9�?5ڕ��|c$��?j-�ɧ��x$t}���f�>8U�ދXH�f5�I��pϊ���K�!}�ʎ�wSq#��e���R{�`���OI˼GeZ��=;%}1�N�VU
�K'N��K5�ë��0�K�n{�.
*����{�/��flL!���~_V��A��؞�Y}��:H��M�0���g�9�t|g�����=�-���%��sO�x��Ǖ�
�������`�&��SVTo��&�<��8�=�y�M��ٱ0:z��D��6��V�� X�S��.�3QƼ���B��ܶ#�MT�����+t�fk�s��P;1���� 5���甆��:�P&�/Nʟ.I�[]S���ո��UvO��������<,��Kc�6�v��2�n���l�E�v��Z��*���~��O��D������VzG���6u�<Ꞣc<"�7MZ�U���à��dm.�d�Q����6�T�����W=�L�K����R�Ļ�HC��:bl<3i�|�cl[����~9��tGկ�%^6�[�e4y���F��8��'|5��ޏV��wj1+aWl�z�L��"�9�NG���o����r�z�����SG2 �~����*�l�OcY��up/"�n�潟s�5٘�`������?��׆�yɌo��ޤ�����E{�oӔ>� �iQI���A��hgbR�5{�P���x�?86��z�5���b��pqu�Q�vk\��B���O�c���
f�|?�����Z3�bl���%����9��)��`cs��S��� ��lG��ZA�ǖ&<DP��OM���d#�O
��{ې"�n(ʪ!�w#�/��w�����.����r̶��έs	#�|��U�3���� �M�Nd���!z�q����q
[�e��J�Z��'�lSkS�c�XJ�]Tg��k���Q=�5��8�$�A_)5V������Xl�7���QJ��#b"�X��=�>}�!���M]P�3s����:;�fh��^T����&Q5�P��o���V�+�ѼPm<�J��ts��dy%�W|F�o�G�+́> ����H��"Վ$���P���}�Һ�vMb�x��{�p)��.�`�5�S?0ߡ�&h!{'�J������>�塓U"J�$��ɭ+�j������֣��:�܄�2��j��+��i�<����vf4�c�Q��GJ���H����X��p	�G�^DV��3!$���U�~_��v�1��0s�+x�tY���C.�HoJ8�W7���cN�S3bkN�	��w0��~=L��]E�|�L�g�_k����*��$��	
f�_b�/~9�	��[�����bn㝢�q���Dm���.��(�ΏM��ώ�N�,d���~�����IA)���r�8�K�dm��p6���k�������;Q����RJ��է�[0�ʛ�1�~���i<�������}w�������⯓��I��MG�N�wӁ_*eML�/C:�<*��g{����a��HJ%m�q6p�@��Y������0r�+��w�fZP����2.�O럫��~��?�sX�!f�{/L-�x�02i����JT+9�+�w��ߜ�kS˲���6w=�2���2�u�`����Ҵ�_;��K0����i��׊�P�IW�q;�t�P����Z�}�����2��6�E9�,|;g�%I6D,�垽$����%7�Ď�n������RI��S�~��q��Ӏ��U�H�GGN�7��y��C��v���H�ƞ��2�y|���{�����sM��`��S�9�7�U�/tP֜�@��n�EQ����"��R��r#�:d��N���i���@��7%^�+�zy������xW������Ec������!��E��8(iIr�v-
��owH�-��x������7�6�B�~��k�8�{q�����s֧
a6��8o��!\����h����g��"������!�[�s�?%�K�>���&(lW6��w�Q;�u��*���Y�mg�gB	>tE���5.��`�*-������k��Q
�8�6GR��#��jͳ{�Ϯbg�K�~*k�i�2v��h��6�ŋx�G�!�_�M1v���TP<� �L.�H��h��Z'�U �x����g�y�u���X��.U�؍v܄���[9�s��}��W�E�i�qh���S��?wշ}vw�e�s��U��;�(�ބ3�!���+��/��9���q�Վ3�Tg��x��=2�#���	D6W=����Vz�y�GW:�5o�$ï���T7�����o�)�~���.��T�q��I��AC;K�-i�O�_$2�t�,�j3�<��vT���u�ٗ�a��
8�K4 Õ;5��//�(�;ܱY�}��93jQ$r��+P]:^�5�b��e��(�O�V���x�0jq��a��Q1g�CB�����9?�c�c�
J��27��a��1���yqY+�����n��/L	������R�qm8��W,@� ��Ӟ�;ek��{'��Hc|A5ӋKQ
Q��u��PN�uǰ�1z�n�a�ͥ�����ok���'����A&{�4�#6ѳl�� .HϊB���e��U&�����Ԗ� �
L��d���X�F�U�OGC:�JZ��ZA�IՙL��Q�/M�u	^.�f~�5�׺[^�t��/�Ww�r[�4%Mg�ֺ�bw�~��G"��K��J�<�]f�f�rB:b��k:��Q�3Bj�P�C���Ֆ��,���qd�b�k3l2WȰ�\V�/�l��(I�X{6���ݔ#Ӏ����ur�Dc@�*�q�@O�e?����"���U�v��ퟔ����	"��uG�R�߁?[f?,mh/�dԜ.L(������o�vG9�M���#�G��q����2�ia��k+�}η� �k�º��/�(k��k��4A�U��g����\4�(�?u����|f���<�S(�#!Y�%�1��n���f}�l���G�^e��]v�@�tK|,(:tU���6
�6�{);q�ǹ>B��G�4�K����2��Ǐ��̄�f�o,qߙ�!��֓C5.����d+b`�+���J-�k_�'�"�<�>�	�������$~u��T�v��1�wL�[�bX�B�,�S�bJP=��B�A�LLOK�J�alP����Dx61�Z�v����e�[�i޿����c4℩|�0��� ���ɮ跼gQ��S#�u��oO��-Zy�+�:�SǗ���ǽ�N�� �d0��t9<�.s����� ���/��F@�+�EY�!%����SJL\�A/�Sh�E���������v���r�?���`ߨ�Hs1ѡ�$1R�N��Z!;����J���tAj�*~�����}�����xd�J�s�������v�v�(��Ｃ�4�z�b��V��Z�� 273��#��z"ؠ6��u�qG���_�����秼���guǰ;{��9�%���6�败�?ߦ�^�O�X?߮�kkk�y�o]K��K�@��x2T�yyu,3�(y\�+������������;Y���_��U��~�*�����b���`���~r��pr"nehb����HU%��� ̛f�����G"���D.͡������]����fn� 5h��n#���_�$�)�����n���zꛮ�9����:.���VU��E~t6	�ߞ:\���h:lM�!/C�䟈},pN����QI͆�A^[����M�>LMT���O���!>�LC��H��Z �KA���)7ȻKlϭ���-?(G����}XȾ� ��s���a����T;���Vѝ��'�yD�|/���OP�h�������L��ÒO"ΐ��V��x�F�̮�q(ެ�yq	�{u�j�x�ai�l���Gx8��N�����8<ԍǎ��@�X���Lד���n�ˆ�������0���_f�ܳ�a�h�����$&^d��œ"qޚ�K1�
�!�C����nG��l�'uV�N.�.���Bd󸫄8	/q�{F�jJ��lg���/(�6��(�T�l�C�Q$|��ȕ���B��ebۇǵ�19���3�*��&wX�6;�W�Eu!��o *����Kvi���y<dE=݈r$�L����x�hK��E?Y2��H��8��d-0>2�k��q%HwZ�!�gv������a7����e���N�?�2���ܼk�2�ٯz"����B�[�������p��ro��y�����5�I)P>	��``~&��R32�����YP���D��I͜.�Z�EMݡ�f�/��Z���ܲ\4�SW2K��1|=��``T�$4l�'M��l�� .}����Kw��NU+-�ߩ6�Kckڦ>7-�: P�F"))�28�ȣ硾���\z��4�_����T.49�!+;�$�0����e��ޘ��n)��&4%6~D9�rISo;��&? �pڷ���IoZ�A�Q�R�`EU3�\�<�6�+/��Y8C�nrJ-�#a��&G���5����qX�Rp w�]�h��r'�"i��	��X�a��(/v��ڣ~v�#c8����7)��� ���TS�#Z�&鎲a~�BD�>���B	5yxI�,y�n�*��h�
���.
�-� �]���A@:����ET�A��K@��;�����ς�[�ŝ�=���Ĺ��|�h��M����:�{��Of�tOa�8L�Bdq�GG��E�M�5ۏ���3��_Fa����ȴ��\B��;bsZ��!�M>uE����e!l��t�EG�]a��V˳�(Pz�B�uw�u��O'i=[Q'����/z�&!��4vێ)�gw�\/�^m���̺�%rV��. [�j����iz+�I��	t�m���迾8�"֏N6#[�Ő>��+@�k�9�H��G�J,R��2��lI�{�#UPX�Z��,���۲�Ў���B|��LWq=�v�q�;��g-N����љftJJ=��CοdL��(Ͷ1I�Ɩ�m�)
�;ӌzN�J~%�|�>n]]>ٌ� �2�KEUīy" *��+{��q5�� �����I��P�R�'�b�?�+1m>�<�,AgV����y��̪�f�!�ˊ�K�Ѐ�\md�v��uu�^Ք�#�鑠��Q=�ٸ����cZ�#V�%�!"��_p��_���������	���^_Vs��뇽��f�x��k̈�|�TU�b$��՚՚R�o05�P��������ķ}�����s�����{���8#$�o����e�B$e;�#�z�~]m�����-�9��<�s��P�T.�I�a����.?�	c�>��\k��I�S��R��z3��G�Hj/�OOrԫk���K��ClS�:����W:�曻���n+3O˟�鋸�#{�Ǜ�}3bW/�DO�����8�	�$Q|^���N��f�O|�������Q�w�)(�ٱ�
�j�>I�/g���E��2wK���tJ��j��؍~��#��4���dE�9:��fה{IzS���\ꢯW�:�7}uP#�t3N�XQ�4����_�4��߹x�q�e�_��1��.����)[�#%|-)ʱ;e�V��'u6-�s�6�D��֟�u;�J/�O����T=E*J��S�&0ɩöo��D�{�,	K%ט��>֑J�	��w�S�V�vj�}��4�Y�CX��t&��^����)��i0>��֛v��lE0��xr�� wD��@�Wږ:Ҳ��zWn�2Du�̙�q�����Zɫ���
���������gh�vS #N�07 �SR#;F��l.cx�lFH>yl�]��r溾��vO���73Fj�r�8���ì\�<��6��)5���<]+�w��j:���b�xѱO�W�C���l���E~&A�Z@��R��1�R�4b8��mӘ�_˷s�vd);:o�}_��~j+�ٚ�w �=�y}�\Aj�9�{Q�h�Rj\٥.�=���^�o�mtȺ��7�t��L��_y�*��ey

��f\ Q����B�f�e�+��*���M��p�uh�K����q�Q�"�����C�����n2ǐy���8����i�v�k���N�q�����\��i�еMh�EM^+���~_;Q����լ'HS,>��m��ܪ��_�={��V�dt�;���d�6O��w��0ūg[�{�r0�EAn,g��ʀ#�l�D���6�I� ����ʵ�Ȧ�`Z��.�w�S|Mg�=���U�?@ē_,rA�P���k����d�3�J���SjJ|T��r�����nk&uͷ�#��xv���:�[ٵ��Q9J��22���ǀb�����A��BJ�F�;G��j�'�B�����˚�L��+\����8m�Qo[�Ť���%#��a��W!&����5M�S�����.�v�_ސ�=��3|����O�ON�}�<�Y�K	�����X�:I3�i�����Ҭ�B�˗9����o0�i�~3jա���*�l�ٰm?�d�h)�_p���im��ՙ�ӗ*u�Ɵs��=���6 ��A���rJ��4�|�J�Y0�'�R�,ԟZ^�R���WvZ�Qɮ�}�3n$d=�SN=ŕ{.�fz0w��t�
o��Ћ�R�?�����g�XCvj'V+>y<F��6�	�؍��F1��>M7�Zq��T��="b��:�YC�6)��6��2�5��H�����k�0gRx;&0�Jjqq=-')/���5�q93 �<�rz��nߕ�YxҦ�Avbֵ~/U�Fko��m���
�S������󆒊�*���}�1�.�]���k/�p4d�o>��՛�f'���^�D�\�m$V$i�xW��C7D����L�^$c~��H/�)�ү�c�<c"0o�[?jX�f����q���j|��"��ND{�P�i��8��?�)05�<\'�q�ȭ�Kqb�~0�^�f�{�l6>յ���3�X���|>�'���� n�{�R.���4�b���l��%n�Qy���9�=��"�=-q��x�-ǿ`��C��^T=f���$Y��.s$HUz�V�����r�ϙM0�@�����K	ky4�|2�_�:AƔ(���;^Ս�A��ȧ ��ʂᄖ}�ݯE"�._Y�_�ڜ���C�6L�FG��D��ۚ��)� nF�+Q�*׺kU���Z�������/ 4��m���~)u��5Tr���ǧ^/o?@��/�-�k������ȥ�yZ��'���F���c����J�����sl�v��K���Y�΃��YR�M�ii��
������?�܈D֧�� �;�t9 ;L�	��&פ*�"�wi��I��h.���E�+����g�	�li���^Y�=�B�EĚ%U*�����0�v�����KC���	��ჽ.��f��&�1�kC���P�S1�P�d���.���a����.��G� x ��3�5L�]3޾����槼=�e�!�8�S���Gg~]�r\��� [�����5+XK�*�gPlƄ)�A{������6��">ev�	W��)��#j�BR����)�1�Y�>f��k���u6��|��شV��$�^ѳ����v�m!�T�����ؐ����~���yL���P��:��{l�erU�R�v�L��)�h�<(t���nXw�E) Ѭ��x1�6;�E0���[p��38N~΁�k��?Ԗ�Y^lc��ǆ���I8������;����3a(&A; 6�WO@�*�oFAx�� &���dc�&�3Y����Ō�\5�((�B噟� ~	�
�]|��$�'n��u��%��r>u@$gℝx{����W��ɊNN}�b�(h��2��x7|WB=�N��)����'"23s0R�Dk�he�Hus-��™���1�5f��񾼛 k��%zr��xE��q�"X�$x��Mǈ�A`3��q�҄+_���,�w:\Cr��}2�~����y�k*��`u���0w��+=�?}t͝�������6Ƶ$)Ɨ��u�s�3NbKx���L��I�gC]�9���ZN�ܖqf3�ǧǧ�U#�U�-��!_���?���Y��=>꿞Go�	�S������n	��Sm���҈\8����h�Sf��_y(*U�L�*�6Q�!�����1�l!��U�q({E#��iy�6	�����j�kQx����]�}������i�E���(��4A�'��,pj���Oˊ�f�,�l��*�f�=.P���A��J�MbL��BŹ��ϙ�����|2ICi?jŦ����S�Q�)���Es(	*�_Spm���޵2E�o()�#�n��]��E@�����]�"&�����N�0���x���V�4�_�s��M��`���w�n�n�JkN�zh���h�⽄s�S������0zv��rB��Y��q�bFB�����x Aɢ�w�ؕ���G��]����aE8�vp�p_3�R�j#"�+ .��:WI̝˒h���8�����rS�� l���n���+�i	9�{\���8WV��}��N���C9���ƽ���|ׄA�gK<�8�.��kY�9�3��h^�b����?n�@&���>2�JT�ٝӉ�д�~2�A���]�P���Y|W�;��x�w�&�27/!m�p&����L�&$�a��A�����,�H�#�D/R��./�Û�`�둯����&^�-\�J뛨��_�@�p>��zj�s]�tu��Uz<s�S��54�g1�a(��q��&�$RL�/��Kx�cGwT(�O	��5KK�v��2�g�/�q��2{�E��D27�x�ʤ����OJ�sg�A �(��r,�2�Ra~�����,ZCTuz�$�zsy�����2�->S�#4�Z�<���%7��@��b��li�I�m�&wc�]O�㾢Mu損d�r�����C��V��`o��4�[v�f��I�q��_b�%ښG%zvPK�E'�r�[�7Ҧy�x���1��`Э�`��.�&aP�/ߏ~�@d;�1��[�"C� A�<��#��������V�j��������U�$�\��E�Y��W�K�
�TjyV�џO�E�p�`�Ir�\�!!��"@7E5h%��'D���U#��Ȇ%YPxUp�L4|8���۾�4K�/����)~�A���7��effu���>��L3@�}	����jl���._�����>��z,�K=:�<#�0}�g�	���d�)�C8��ڴ��]>�ES����snğ ����^ �K{��\�;N��k��Ī|�rʜ�>qi.��t$W1g23����m|����.�T�TQX�t¦���O2�E��t�4OzŜ��sK{/|3׭�fx�����t7�]�q��&��daI����T_}1A]Ooc�bɘ박>�޺��%�T���|�8����� ��3�o-@u@A4V�[� ur;!������cVSg�#��qi�A�t��]!iJ��,쉟��p�~�w8����8��c���q�J��z5n�v���d*ʃ���؎m�"�@ʎn���!.1T�xb�z���b���"�E�Y��g�w���ο q�vy�,"O����t+�x���	?f�W"ǁ�]���S�Us��ʹaK������J�vE�~q_�ǡ@�-��WR�C�p���A�Ǭ{�M7|�*�^\\iФ:�l[�������%��b��x|�'�__wď|j���j�G�JF(#f�ڂ��C{�����~�E��o��	Bg=M�@b�0sT��A�������} �MθВBO�q\( �Է<=��]vL�f��N j�"B�|��>�b�S�$ѕ�IN���Q�o��0��
G�Xϵ
���cV�ǉ��E��t�^@�-%2�b����l�"*��d �ξ�ge�!Mň���X��[��B�w�+���!sY��9v�%����� $���_�=+�[2Q[������K�^|J�U���r����_4a!hJ1k�ɂ�ǳ%虘T@�qz���6DK�c�s|�)�����t�绍�F�	@������pP�p���>�M��}(x���L|�L#�8<���.�� ��[� ��=��M�X#�nn0U�]�V�v�|Ρ���淞����&x1�+���� �q�+L\�fNJ%�Ӱ%ff�h���1�� �VvE�&�ڥ�w��=]��3T��f��m4�I��tZ��é�b9"��^����f"��w�����?ԋ :ڂY����� g��;:��X�$�����Wlϭ��k��Z�gD���Y���w��[�^�>�:\Ԯ�["�i�;H�<߫�-�5
�O����Y[����h�|�n�g�q��hg�Lk��'�i]���I�� ��DoWY��ۮ�ij�����Z?����α��e��{^�b�t��G�}����p�$�-���<�:_��ݮo`�<&�6a�M�F+}�~y�T��S"xV�W���w�d�%� -�ٌC_ծ��	�m"ܽ�����؎��ⓞ6��M�I�t����ysY��?�m:���h�5�0���U�j�]���I*����#�Fx1�������/4�^6)�ݞ!FS,�J�/\��o�Z̡P�q$�R�ߩ`Vf���i�~�1�O��AeZX�܇�]ȱv���}��7�Ppk�݈L��y_~��:Wa ��	g�Z�f�ڌ���Dn�Xм
>N�f�ry��xP��J&6��:rܗ8ɶ��;��Ү�ms����������8���e�_�鸾�-6n���R⥧f*�$� ���o��qL����� ��ݝ`0� ��T3��Y����Dc���T���`�M����Ͼ^m~��h�8<�Z~�JH�~�z��sq	�v^0�G3:yD�� ��^�Z~��U|��9Xx]���ѕ�f&R�]�b5�3�h�Iؚ�O����t�Nҍ��+��_�K*����̦�V��>2��K��؏�u_��ʐ*�r����Z�}2ތ���fێ�~�?}�؈)���<�DP"cs�������p$����z�ض��ק�t���H<Q��G��U�/�9��בE� k@�u��X��Vp2es�")�|w)5�p�����*�:��y��$O���8�u/����~`k[�O�lVH��y���Vrd�AP���_ų~o��O�,�y( ���U��9�W���V1�ƏT��tnz��;_���-,�nf7A}G��J�_߷-ҷI�=�B��A�x����fZh��*�:%�5_�u�us>���x�´T�*V���nj���"g�RvV�����	-0�ސ�[L�Ƞ�=D ��w�`iLH���W��@h�gvz~�"�]�?f d�t�MԦ��9#��>�Y,��5�O[P�bQ�0���"8	���x� ���=�?��F_}9� �o�>��n�@���������	�]��^#��ۮˡL�~pF���Gz�=%�;�a�ת(��^�����NRĖ����p �u��^d��k��%�R���|��lFi���Q���Vվ�n��)taJ`���w�u�P��Ni�r�W�C�al�{Y2!p"��t�\D��n �,�[�Q�����+,���.<�s����{Q��D��C��a3[��z��bqWjX��/i�/G<����o����5�<�fk �y����7�������*�l	P�7��=��]����.��6�mn��a�y�\���?�
��A
������z�O��=R�Ⱦޖ���	�X)2����@(���bA=Ծ��#��+Ǖ�x���f*�	S��K��|U/�����0�TUs�{���&�"R*�(�D��,k���}���C�8�����T��K�<�Nq
��}��ݪ�!�e=Y��UO�����A�m�BIf�x�����ʵ�����9R��ͿJ�N�XÚ Y���������>���˗F$���4�OR?|�!z�ލ�x�
�������ʏ���r��zK�K��ѷ6��sda��N����+ҩ��;��}l�c���Lg����(�R�l{Ĳ{5��3[�GKYQ�8�W����$,ڢ� M|u���/0?�6��\�k�ᕱ�?�D�z��GHf��p�D�۬~�28O��3���?B�r�xQ�ˢ�9� ��:|]B��֧�;�{-i��f�T�;�
AS�f}�"��}�3=r�BL�~y�(����[�Nr�&�-��	|����V�����Ty5�IO����q��U���N��x�cѨh�*�)�}�fQ?��l��V�<LG .CRV�(%ɞÜ1\Z\�h��]|�]v���6w|���r% �j�D�������@�y>��a�R�����0͜�~cR��@��r�\WOy�ߝU<)Fⳍ]��t�=�+,�������˗�r��Kf��xaE\O��u����F����:�z�;*��+x��!?�G��_Vu�N�F�A�O�=-��f�����0�Y�A�=ќ*��4-���'+�T�UF����z�d	�4����z���I䭼$�SN^�@�o^6�L�}e�����17�l�[J��w:	q��SL}ڰ�O������Ց��3�lݴ�emr���ޜ,�r�:�7f�@.���W;���Pψ�o�0�/G��Z\w�[���7o}mO20���
qRZ(|Tu ��~������a�ڈ��i����╰�����l\=K���z��%������5���4�y�Ā%dkSs`���ߪ�׌���'��*_���['��U�{W�uǾ7\�ǞO�KN�O��3pnqឡ��t�~��~��JJdh��#�g�=��R�e=B<>����p7�~=z��u�\�+\��AC8<��/Tq���I���d~��8����V/vH�F�+����#$��GF?;��[���w��jq'_:Y����Gn�|ơ2��^R���x�'��U����B! y�!�[���m@�Z�,}���ig׺�Ao��g�Q3�\�7ӵmR�*�)c��ǿf	G(���`x�庈�~|n)[G��d�'�h�9�(a�u������F�$��@$�Rmu|�.��^o)��5��0�vR�VL���`J#���؏У����H��,}��'��)t> ����
�yď
� oYy���Qw���RI�����^���.lJd$��V��eV�8��iy0v-�+��t�?|lܽ�5���xT��,�C���rRH|��H�)㐺���/q�!��82p���Kc +LR��AW�E~&=�{'*T ����}v߿g{�7�6�;�DA�gZ�:noQ P)��h��(g�i��|U��DU�n�/1+�zu�N��-�DI��D�-oM��A�3�$� �7q=���n �ا����k�n��(��^7���t�B&A���-��[�V��5�^�)����B�Nl:Ųs�T�,
 E��B�M������E!z��HbM�=D��SB
���H���Ěc�H>�g�������u��խ�]�1�0M�7;�𵎊A��C��7 {���ڈ���ҏ�I�,���|z�c=u�!�pMX�j'H�'�r��5ü�J�ꢹ�����=y����
T��0����p���V�;�?�=3zj��\S�c}�����OeC����5}]�X�����De���Q���ˬ��è�i�W���WT~��M ���=��|�@�B��{��7�Qg5��ή�<;ijh�o��]�"^?�';+W�}zp�1��)L��M�Ԟ�{׺��ee�%�	PKĭ�M���Ɍ[f��y@���_�l���܁ �އ鋰��ը��������?W�"��T��x�J�e̢w=��I�(�i�����&N'����ohi�)�j���`�jx51�B�H,DI����Ĭ��9�~�T�$�U�XH���]v�ľ{�0�o�9��8ǰ/G&[�t��e�O���A�c��駯iX�+/��%K��<c�]$Gw��C�U���'���g�,b��zR|�su|m��7�p^���B�=��w�2`���.��w �S�/?�@=~y�ٶQ���q��Hh��ZWRtO!��n��_��y����W�BV&����l����PFX�I����=A0f���ҵ۸���zVV?� q���c���]��&�I6z(խXX����I���&�G��aO!���k-1ŭ�m=-��1�/���e
rc����i|_8�������O��8ޖ�����๎�k���3��`=ViaL󥄩� ��~���58?e�"�������g��[��V��?��o���}'���=��ew��T��D�A]MҪR4�UK$)�H[�a&�n&(=�3�~k�ӪK:�0�Όv8P��(�$L��^`fr�*	%�y���Pr5�W�AZÝ��)0M�6\�Q�-���(��hFU��]��5Ț�X�ʠ�/3�W�ÿ�ĸ��^� t6��j��_+4���ʫ�d���Xk�I赒�����)���,�97[FbW��rd�,̂a�a9�G!&�ްYi�3q�pI�HJЩ�5q��D��qn%���z�ν����h�vӜ��m	Q^�N8#RM��@ߨx ���Jvr��"�Ҍ�
�?~�,�)�z{��0�ڧ�������G�9��ŝ���)�|j��T�c��v	���L�x�l�����"����+������hg1es4�!�1���7��q	3�P�oD#�xi(*M'=K\�=�O�ٮ���ֈn\9h�ܨ�H.Hi]�a��"?t*[:B�5>NV���@?�>�}c����������V��(�۪��ڤ�4�O9$���2mR.�����yvA����asں$��]�<R��J�n���SIq9a�M����pRb�!Լ�T�Zdb�C���� 0}�3�]�&�`=�D��h$QA���Vɧ�PT�T�q�[̨�/�54+�ጢ���R{��ʸ�Hl�1)a��x�O$l��J�;T���J��6��&GJ_�Yn6�O���Ω��H�*��a��&s�$a�Qa����S+�k{i�sM�4�V8��\�V�k!i@�ǻ����bt��j���ԕ���8+��J��xe���ݯ)�����nЗ�,x<��Fd��H܌{k�ɋ�3QtFd���]hd����@aU�,�*�ͅ�z>f�0���g���R�Jtg�!�z�`{<�0?����`Ԛ,�h.�n�l�]А����i����@�x	�0-������R��I)~�;\�?X��5��L�$�<�pX�>���
�\�4�8i.����G�w�i��(��>��ˡ�.ñ���r쫫�ϷV���T�쉞;��B�^����i�]�v��M!!!aw$�{���d���5m�d�GQ��7�UU�C^�G;������$�\:"��E�%?��ru�xԽ��s��4)����3+���}^��s^Q�F��Ic�ߢ�ן�<�"�@&���^��##)v��t�e��:�ϒ����pzqƼ�q�N��@ED9�9)�d(s��zР����{�A�A����r�X�a�ŋ�ö2��/�V֡G�ZM�T�U�8�P􋉯̠D1�习Rf���#)0v=^ǂ.Kڮ�aPT�^~��0`	�αB��߃yw��)?��ox�s�^-�:�TvO��Y������{v�W*��P�u��t���F�cJTv���h�RH���4[i�#�`�Pk�# ̇��'�e��w����=�`,I�*�Q@,�d�RI�i@ۆ���j3I�j���Vh�c����r����a���a�����!cn��T�H*O��,�X���7,���L�\���t����Я�҂�莄����9	�ɶ4��p�4���셩������1s�ߛ���A2v�82�>Wr�ul���3���x'wv�_[���K]�5���x�U�._��+��,���Z�bٹ��y�p�u����8c&"HȃnDІ<��e�>��+(�2`�)]ez<A:�)y�����T2�"��^�ж������_��`����p�R:��<��<� V�
�&��L�{�K�B��\z���P�@! �}N���ݧ��%v�T�j2=�
��ce��H�)Nf�\~˒�u2&���r�x�7x9(m�pN��vn��X ��k��.}8��������8�}p/�;ȧcD���d�rW4���7gڙ��]wF�&���zp��-��-�v��!�9�Ŵ[�Ң�I�Jr�HUiB.�t%CdS���åB����f�LV��U�E�.	�
p����]�ߕ׼U��bӊ����N�ΉH!�&��F<�~�?��SI?�b(@��~���΀¢;��������.��^�����ӫ�b��� O��Z��ʩO��A�����mϛ�&�Pn�lC�'	���+�|�E�j�CW�S��;���WP@�eqG�?24"kj�a�	'G>ż#�6�$.����6��Ƭӌ��|"ӃWeXa� CoA�!��tGB���9oK�v�!d5���"o��z��y(cڃ�_y�8ś���\p�1P�)�N�紓jkJdtu.��֮�d4m�@�ʵۯ���/?M2>�V�I���(����mfġ]g'�&��s �k�9+ ��{E*#�����h�X�m}�8��'G{���� ^��}mǉ�e濋߿u�P���'4�,vYS,�}Ȃ��sC�����Ӆ�I7��mu`�;�R�}����Jц�鰕��D�V0��1�4�	/{as��m���C��������~p�b�G����!ڡ$tA�����_��3��`U�qXO��nDi�a�֫w6��ܼ\�
qu;A�)��ʸ������7ιSdS2�!Nfg��LX
���\�3M2��ʀT]A'���>�h�Mh���1��ޒaj�����+�`!�7�4�����;ժ�S2m��	W`�����k��w>a@�뿆�[
,�,�)cn�i�;qcY�������>k�]X7����څ9�IPR`L�|.
��f=n�Y��4QP�n��h�$w�O -o�\l ��s�}�q�0�|�eA��;d���2KK��$����w�m������΢��N���98K�$H�6�W��� ��6""������6��ʀ�	-���Ս��w�j8c���`	��NCPZ ��3���;��/����ipP+���t�d���ua6�B�q���e-@��K�VP��A>���cMk��KlN�`��bN��NF�K-r���-���;G�����EF˝cmu��r������H���wl�`=5[�Zx�=iC-ϐ�X�٧�̰m��p�".��D�U{Y�U"�qNY��d�oq5�N2y��ZonK_�@�l��\f���&g���6"_�Jj����i'0�8QSo�B^�٥�a-����BWDJ�#�(�Q�p�cx
��SmX�/����ra�ݓ��o���%�񵂳�J L	�r�g�%������S<d�#��,C��ߔ�Z;�zs�ŝ������ۧH�K.�x$t�4@wd^�x$�d��A� �-{ �%�1��^�v����W�>�r�[qW�@�����	�_�t/��Z�׬>��w��}����%S^ '�p��A^��^��}"@t���e�4���ɶ;��v�!�hd0���{U��a~�/LZN�!M�*7{\�j�7�v7��0�(]�Y��g|����ja�OH�wg��\i��ө��="ҝ� � ����ʭG�XQ�xE�ˮ6[��;����l��Es��; r��]R�]�ȿN�ھ�;�q����!]�b�m�Tn�ÝJ��aǶ��z�j�U[��f�O�.Fh7f �^���iAn�/�7nB~�¾˾'4�-l�|n�}�h�+�Դ���5����l:ܚ��7\��B���ŗ�~]���D/P�	�z{����|25�8�[����݃M��������؎)����a�[�����33�:�%j_�>4��+��Z�3R(����X���ن���%"w�MT@Ro�=�bu^8M�:.�Y���"Ѳ ��Ȳ�D)�U��G�W'+��2;�/���ᑻe���Hgލ/U��w��,�6��q��?�@�Wq<l/�[���������p��n'��p�l��A-f���n�������c9S������Q)/��B�>8۝H=^��|{y�-�^P༶ѕj�(O���&D4���8^�Â�:��o~w�9e�_'�GpD�bP�>���(x`���*�T5��Fa��fE��21v���c���r�_�A�m�[�'�+��)s�s�"�X���x�W�N��_�=g݇#�P���¼��)�.�_�+�P�8�~/�����{f�!^�0S��C���B�C�5��:Y�C�>L-����� �hӢ4*,4Vi�A{�%���ғ��?���-�N7�e�s��Ur6��bd�{<��4��>�4L�}{�ֆ���Z��J������4k���So������{�F�1k�B0�G^��H�4�&v�����7�s��7q��$ O�'���/^��SQ�w "hk�����������K����Р�@�Ħ5�N��%�mah~Q�9��ђ}R
�+e.11�I���ryWv��1_��
��'/v5�F���W���ޙ�:���I*�k���,�l)�T����s6�������5_�X��)I����RR?c�D��W���?���¤�Tz�D��h$���#�(o	F�.��Ý!�(�L�t��}p�|W����힆�;9
~] ;&/g�1�N��r�����w�d)��~��}��y��$=�;e���kG�����Z�3;��0n�u�k�#�>\�Pg��l�Q���*����!��7=��e��!h@`��	g���8�s�^�]�������(�I��1�|e����v��QR	3��u��x��c�ó޿�R����GB�S�Ő�&B��e]���ѥ@�9u�yO�Y���^x���з�%�6��#��/�8���w~vWA����^�$���N{,LC$�	 ١�ޠeXm,Ұ��d�cB}�}���˳_
A��k��}���F���� �\�z!3��+�\X�S(?�D�)�L��hPHk�anBP�o���8E�[�`�l�;�{Q(�o�B��}S�����7m��X3��+�RJ���d�<�{��y]�i\�5�-^<>>o{��9>�;������SA�[qa߿�/N����L�|��g�uywW��k� l+�3�����`�E��plowJ���f�Ry��@B��o���@��X���+�,��І��YS��p���x`������!���l���52(	�d��Q"
9�0궅��e-�F�V��]�n�:i��a~7�����wf�$���-Ǒ��9V!`b�`P	j'h�rA�;�<�������k�k�	$F�d�5�}�������o�䶚6!G zS:���X5����_I\��aBA�]Qd�]�
��r\2d��"u��8��Q�!}K��Y�o��JvzĽ�y�+ k��9B���P&�퐝��:U~�#B�Of��|�]���c��S���<5�U���b���ƆE!19���3�{�)g�7�
�Z��3�{ï,*3;BWh�=��n��:�ci7s�-�з�Xm�b%_m1{97\��d���i�0}C�}�tM\��;���ࡸ��{�4]Q�yJ}�SS+�M�r}���M��U���p*�T�a�	�M��<���@�>���G~܏�Ь?���߆'��zU��q\Y�]�+?f���ajЊ��f�D���l��y��V_�_b��o��Yx��Z>!�pCW�b�
�L�U߳������]q�O��j܆��%+����b�zw������-	FH'�oqi�N�p!E=%x�#��9o���.X��4��$[�N��U�Pl����]y�Α��8iXI
��ջe�Y�y:j��Y��8j��"�Ҳ՝�;ɂ�i\�d��Mn�p蟸�<3p���֓����`Q�R�\���1Q&��3����nJ���q�}XwVy�vI ���* w3t`U���M4��.�v�j��&�v�U�%�m����A�4.:���J�$f���d�<C���KQl��(Y��VǍ�S���M�6�;��6z$�;XlL�Bќ
r��\�2c��N|_��GY��0��|S�M���z��|%:���Q���}���1L~<��B��§ŧ8,�2����^���؃��rr��/���Wu|p�����t�����G��<V!�=+�Azb,��GS�"D�����@��gr#w��  0�)�/e뷏��Ú߰0�*��2�dj[GӞċ��z�|3Mkϰ/a�4Hԍ׳n\N3�C���������ag3�_�������.j[�K��J�r���s�OX�l�'*��4���E5a���}�<#ꆽ�K�������z� ��^�M�Z')������U&�]_��_�f��	��O )�/�H1o�˿D��Ud��H�[�w���beM0O���N��������Ա�n�89ܒn��>.���䵼Ȩ�ǔ���������~X}�5g<��\a�X�C!�/pt=J�m�#VH?�|�T�ݭ~���C\����<Ɣ�Sd����TjKJ�k�\�g�
�2�?׍��Pn6%��խ�-�wf��M�
ڹg����c$i�H[�Sي��1�c���w�c_OӔk���a��U��ޚ�+�*��Oa:+f���Q/�7�hQ[|>���ԎY�}ث�0��p���k$}�E�-�9�=�ny�%_FL�V{`=�8D�pD�ݸ��GK+R~A_ë����K��`�mae����n=�n&��`��W�q���rP�Km�\�5���
+*�tץ
YϠ�FR�Y�.�BK��O�.��Ka��<#к�ˑ�
������2������H�/�}@:���lY6�v`���{�k[/�Ղ7V�݋�*;�)>q���| t�:�66�$���ȓ�4�eke�������κ��x����|�ss��<�׾��j?�|<�=u�!�AEٿZ�����?%��]����k�A��x�w5=P��+���W�p0��w����b�b޶�\�1�O?n}>��*5�j���m���j���PL�S�l$��믂�en�W�Z�����t�rg()�R��^��\�#�E�w�@�%��g�Y�uO
�U#�
�G�U��
��N)z��˝�/n�q�J�*_��/=��K��H���z���:��֝��\�y��
t ����L߱2H�#:��0�tٰ��G�r^5n-���mO5_/9��A��L�,��YƆ����͡~���Q�Pq-��4xp�@���[p �ww�B �����w>���3�~���Z�g�tWW�Ou�d�aX
��=��>�Ex�k߼vi�� �����T��$S�l�"���1k���}��(;��1ũ�ʪN�07�a�c_�E�����;"#�q�;��[gx��y�?%��EĿ�iƸ�0�j�%�� ґ�׀��ZR�]���T�`o��)ɫ�."�zMWtUV|�2����:<�r
-�0c���E�w�i�2�t�4.K�֭~J��KS<x��`���V9n���J]��[�D"����z��[I2�f�-oG�2��3 ����Ò KM�p�'B���e*Q���,��sY��>n�W�j}M���瞉y�h�?*���㬤VB�6�1��8���r[��&�V�~i��B��UÄ�yC����x�^�Vчv'���	��i)w1LU=��O�|;"@d�9؍��r�k��� �����;�p�o�`�F��.�Vk��F󆵙3�\��S������|E-�Nx(DGKkCG��fnш4ϓ����e�>�h�����W4�L�	2f(��j�z�gp���4�.���@��i��xc��ӆ?��
6��=A�~@w�L~�NPq��&'��:�<�W�>VuuXf���޵5xn?�<?>?(pg>� H3��@��p\�[�+����~q���8Qa��<��Ƨ X2*�i�+8R�&�ofƮ�1t6 $TV'��q0�6�WNOy]k6U;�vŧ�z���Q��k&��ud�6�1���/2@�������(5n�����u����U�����:x�b�I�|���S$"����Ԋ�N:�[���;a)|��z�=y��u2���1���,!���ij���ۣ��D�����oC;&��f��=�MH����!�"���I/pl#,(
v5����c��p�Y}(���>u��ּ(����+�,����UWq0/0]�H������;�9��;[�~��������u�S���,�Ǩ���7��GWy�#���Wĕ����m�[m��I�um��ͺ���ЖH����
�f�U�#����3�,{�z���0U����J����y�3��{i�꛳�B,XuTA�>�B"@�t"%=!��(�Ǧ���A.	a����M��%��������nw;h�\�7��/W�)����M����-�F��tZ+̈��nsF-����kx}F�tx��^R��IP��cC#+8����3�đ�|�|����~M��C̱J���q�P>��8��o�D.�d ��9�!-��q���׻E��_1<ܛbP�����'��h����b�1����l��i�8�(l�J��k~f����.�x�5IP������C���}DUW�2:V't=Jm^�H�z�E�C�[��0#��̊��>b�R�ʪ����ەG/(�Ω����2_K�����Q%����tm���[�<����Z�9�N�����շ!�����'�[S��� |�m��l�)Gh���I6v}��F��f��\)z]�$>�{�MC���T��<��8-v�j���$j��ϝ�U7cv�(�`a���G�����D	�y�<0f�z:�����)}�X�ZSTd^�+�5c\�,�=���|����5e��a��%Q������������p�|���h���d������j!̾��ni3l��*X�2���ɶʪ����:�yw��*���k����o�{�t�z\��n�Mo�ʌ�#P�NO�������
���� �+y����Ո�E��1X��g�\f3,�Mј�V���O���vC�q,�=\�}�!F�hf���,�8c��ʸ&�ը%"��춪?^d��7�W\IJ���+*�eĨ��*��r`����1��!�	�"��9Ox
���3f'y�O�$!��B��Y����Yp�R��E��<r�����ʉ�0�L�v��� R��u_����}���i+NS%cn�%����Ce���g>�g$�Ya�����}&σ��}q@d�R���,��oVk����[]�D�Ƶ\A&r:qzsI�5�/]&�k�]p�)�L��<%k��s�D�"y#E��U��2n�;�@d₭K]n�|�y~�~��`��I�g���J�	I�R���|���D�|�1v�9U�l�\2S�eJ{���ߎ�3�L�I�����z�6?��H��@��Ͽw�)�8Jz�<�@��|&��I�$��:�{�4���y5�[�.�hƍ�{�%,�C���aIJ>�k��Ny>,w�,����K>��:��,y,
[/�4���Z,"(�����jM���0�ҹ'潿qP!b`׆�:	s���89i/ݳDո�1���,a͙���0:���������I0`c�����{m�������_�f5i_m�NZ����J!�:]˥s���8�_Ԍ��LY/�O�lg��������(,2Z�p���/#92�΃�������θ]اS���'�,8 �����D�k�<�K^�e?9��O(��8��m��.�W[�d䊥DI�v�u�>�)~�S��,Q9;Ȋ&�$�`=A�k(��|6�ا���[�Hɐ���c.;w�vf?dQ��g=��7_21�
���7����q��%3�v�y��S$��8-Q�rЬ)n����@u��E���"���;� �:�|�4��9GwK�+4�9n�a�WX� %-p}���Y��[���Z�Au�lԥy�@cy���ߦ��M�[��֜i:+�)��"�w�62ϧ�ekF��Q5b�:<̺�O��(��֓wno쵰�a�kdI��Ӈ�u�s�n��
$�����N �Q�޳	6zi�a��(CkS�K�r�~,���w�Wӧ[�F�b���cΛ��#u�d�-����z7�D̮�i�6���l4�<8j�����}3�K�C������Ӽ�/o ��}U�Wk�OQcΊ��>��տ�1� 8c�q><lƞ�-���X!��t4ǭ�����	���Y�m`��F( ���q,bgX��mٍC��7\^���Ž��\~�b�}U�Sl���	}*����{~TȚ������بᇊ��h�޸�(0w��avQ���7P>A�������ᆜ���\��J���ݲU�qe�ZBzp�_A`�
�!�a�A��c{���u���o4�h*�%���N����9P�N��Q�P�Y#*�ZIE6=0�h���q�	s���=|�F�ږ:��=�ݓ���Ɣ�j�T����X���}��YB��Rύ�)�n�l�~�,eLFY�}��tZ'�ǐ�1�����M;D!R9�S3��13�Y:n�$n�l4�FO`������.���#��,O�S�r�y��3����Zj�В���`��٪��kr�q#?��"��'���<����߬������H�����>����fk�F((M��Ί�A/x+W�l�O&P��̺1\��c������f���� Q֚��{;ÖvL-Ѧ���Gg4\a����B���W�i��7/;Q�"k.�����{�~�p$ �(�bf=x�_�&���+�-���9;˅��*����?=��~�H���e:gK�!�h�䭰ױ�!��H���ᰀ�Qג�e�?G>伳0Θ�L������P�@���3�O�D�E��cH�S��ߏ g��{g4�D���*�X�_��dˈ�vo4��,*h.߮�x���v�ʢ��m�����Ʀ�9 �|��P>��s͗O^�"��x��^��ә��ӝ�|($2�0�(ݴraS9�}��8r�|#�����'ڋOq����I�����\b�/jA����+�8�� ��Ƿ[F�c��<y�*��*i�J�]��he����rX~>,%���I�B�vu�T?�!ò��$ڥ�CQ���U���x��nu^�l��g�!�R�c��Kozz|lAn!VC�*/�>t�F�����3�i��#=�<���}��k��-��'�ҡ�;��dx�1�3�n=o0e֝�q�y���#�kH�0��1~|R�e��=M�$'v~'�Tb�^w���v<�;kƎ�澇;4��>Ʋ�����H�� �|��3&n�EaQ��L�c^�E��B�H�9���<[���kl�--	�(���7��2E?L���=5�~��<�5�%4	h4��z�4Ğz|}�IF�N��r3|��n"�"�7!`z� {e�<�0t��3p���a��������fr�:a����$u�C��� ��l	=����ւ��8*��w�����v2�]=	ڛ���f���&P
`<1/�?wd�W(=��+�~_�L����aN��r}��2�ߙ�r@P.t�e��y-L[D��h���>��.���NfDH^_j����D��AW�J�ˁ?gB�fόv��'���[�H����������#`�%��]+�+�c.eq��@�5�>�Bg:"���"��+Q|�응�60�
cK6(�Q��a� o�("��?%.��f8��t7����eLƲ�	��~&G��,�)L� �F��t̬x��q���7�x'5vřq���N@zj�KS�H�Z_�SϜ(1ύڥ�t��mӑ�En�KtR�6x@�þ�Zg"�xbT�~c.K�Y����ᡘ�F4�coi#�G1	M��r,ͅ�J�K*�#��m�A^If[��m6���lq�t��ef���8�h}�G��m8�i�T���GP1��Θ���%��z8^�TP͖\����(��UweCՌ����*E�;s�7�����`ib�I�U�d�w��u'�<t�L�++燱60Γ�J���Q��E�@�oYg�%��8ˆ���5�ʄCb�&��Wo�ߕ2E��&��0Y���3��5�Ю��=��Gv���
ȩu��x��#Zz`��=��X�(^��D����J�����݅����J��Fxh/BQ��\�<(���e�ܥ;��w�L�����L ��׭�ACռ���$|��d
߇��'�#v+������n��EG��+���)��N���
���u(o-����F:9s1;ó/T?|�z�^�Ux��e�
��4.� ��^�y�;?$	���e�B��y�����93g���@A �C���ҷ���"�42R�R`�x#����b�zV�����)t_��E3��W����%�����ߚ'�<�<SfN�f�� ���AX;�	��������V��X�ݧj�dѳ�7�K��q`UX�X���GT5鵎����� mP2I|v��ūR���k�d�H ��L0�p�g�gK���jѮܥV��Ds�9�fK+�ٱ��*C��"H�����_�r��6т�O�6�f�z�"5����Ǖ�����Ć��rP�_���.���7��FY��W(������	J�M��>Z������@���U6^&�}[Ey��|����zhKK��#��e8��.J`��n����=u�$*[y|��@���_Ȃj�΀�����:���>�y<��__V}�,��2�ܿ���Jy�DԺ~���������4���4z�6Og���O1<I�{�{���3���S��'.�-�P/����%�e5J��������D�x�{Y������(����N�d��=J��EDq�L�9�An·3���S
pW�0��
�-PXl��=�W�MQ͇SSQ�x�,:_�}�c�z "6.�!�\]�F��F�(�e�M��M sd�ޫn&"��?a�ު,ϐ���'l����i�*����{J��ׄ�dX�"��=�-�Q��vg�p�8��3[ZJ������]9��~���6����N����47:�	{\O�ղ`�/�3ۀm��f:}���apW]��k	���j��bQ�|��%]rqS���D��:qs�<rnv���\*_�l���@?b;;b��/w��V��A#�Z��>��{cMF��N��<`[.�'�rO7a�`Jԁk�	b �j`i#��O1�ʃ�$�j_7.ñm.�N�)ȭk:x)��MT���2
`ht��H^�I&�|�z[�s��.w�\V�C��H]y�@-���\�=�մ��n��U����R� gX��6͒��Ğ�s�Lʁl6�`Zh3n5���<�.i�#@�}p$�]�!�0EE�Lu�2w�	GG��ɏ���%a�VU��.zc�Ii���ʝ�.㒈P�j^C{'m��ۭm�~#ba&�
JII}D�< ~��Z @�O=��(�f)�Yc��A	{Z �֐�|Y%�NZ��hR_��$@!fZ�Qe�P�+�H�^�����?��i��=����yM�(���F�J�-�O����GR�dv�}�<�(;ffC=�6[q[/�.�Z��nl#�` l��Y��(ia��ߟBG��ok�m���n<�Gw�1�Y��6>�������B�f�Vs�p��h�yDV{�b�.�yl�8�J�=�h,�@�m��e6\��%I�<V��5F_PԟӛH��%�D
�e�D�o���(�[���D���4 D`�e���V�:�ޫ�W�D*P�A<~!y�Y*�7�4X%O�H9*�%�XHň�{��x���ϡ��E�J��s�P���`��M1w��D�,�jg�*��b�=������)w���A�&�	�����QM�F�~#s�ztn�osyڔw!�4���z6�N�?��}'r*����צFϣ��Ϫ'a�+>��G��w�"?^ta�Z���+'R���1Ի�`�&��@���Z��b
7�f���#�6�Ґ���Z ��2pG������5܏mTs׿�Y���l}CK�a3Z㹞�xT�Ҭ�]B9��5R��w��ؙ��f��#/���$�0�� �i$�F�Bi�P���Od�:
�2�cM���ŜVƍ�ƍճA��K\^������OeE��`�����R���L�9� ��KS�V�M�:�O7���Vٲ/_�i�Ig^!�����k������.^��S[1���1N[b��f~rݲo͈������B���c�M���A2G��aX�|�w�Z�Y��ҿ����Z����U�ب��X�A2z�2}�̣�_���z�l
���u��A��R�N��J{�I �F�� ���F|�D�:YrI��I����$7"�����ua��P���ҏk�M	�b��c�ז���u*��\��Kg�MiT?��M�n3֢!����Z�{��3
�8���4�=�e�<�v��ی�}ø��~v��h��JS���e�K1�[�qz"07�i��V9ȇ���ꃔ���و��`wuF8�o�w�Z5h??~�	'�UZԡݘ�A[�"z�y�P �v>�����\�ݠ$E���H�xӪ��HۗԿ^��s�]���I�*��a��w7���Լ�?�r���h�����YO|�qPC�h��)�]}�V/����?��k�ڒ��"��͋E0�A�����}�!J�2���I�8�ns!`��"��ǃ֥ 3,<���x��`�cT�T��í��ǊǱ�u��<��ヒ�$bo���a4�z���R��]6y�X ��;����5;�m|��b�J�/�T�*���=t��vM0��屯=F2�(��/]�;�>�v.9����V����9�k��Ds)b��-v}Nn�5�W��>YLg@4�x��o/c��P����)�u�9W{�7eLɺ-1�~rZ�R�;2`�t�eg�$	��f�9Z�i��$�((��h���O��
�t�������W��[��+)�i�����{�20���V`LJ҂Jz,��.�|n��G�BG����ۡ����ɛ�Lqߣ���-�o�����f,6XW���D��Q��6}q�'K�ւi�u���f�h���7s�p��7�I��x����҃���yķ��~G�d�6���Q�����r��ۺ�uR�Q��(A��q!��a��wrM�n�. � tv!5	�n������"�
W���Xw��:D|w��Q1r!�� s��>rn����\:S
�QC����]Gɋ1���/�wvn�ӵ�i�}>���+��*k�~}W�eK��C�\�Ǟ#���*�c��({�pe=�+��;.�����W��	�W�v���/�D����Ty��8�c�F�X������a,s���lԬ�`���H�ڬG��8lt��@+p�C:�H�k>��:u��%)%���*y�����h��6���(�9�=L�p%�-���+qB:zo'߉ٗ��{��;ݿ�R���y壟Q\2��_��v��X�Chv����?ى:gS2�� D̕�c!\/��wN�[���Ծ'/�x2���O+~��Cg�[*G�f�O�s�����H�	D�����W,�|k*�!�]�ZtT�������3��B��"~�*��>"vN`F�,J�i�z���D����/���Ǧ��x:7��qE�A�A�9�BH��@I����R��Jg�v&Wg����ݑ�,f��:	fj����ғa��0��L����(A؋m�pt;��jwr����lO�~RQҾ0h�gy�����K����
Q|ԉ
c���C� �f�bj��Y�^nz3teg���
��vS�,��Wˠ��'O� m�ŏ���6`^'"�`L�����v�2*��<xW�T���V�}���ԇ���U7���}��������_�L�=tax�n\4x�(�yL�2Q.�NV��X��pD=l\�̚��Wl,�V�:�����q�;��o,�[`F2�s!/����q#���<�ً��r��o�q��
6�?V�
���u
�v�������J�Ի�ɟ�ϔ��E^�K��t��T���;��br�̯84�y���MEh�jF9�<��bn���=���LM����ˏ�̝������'��8+ZT	]�k���������z�`�Ꚛ��V�]\��\_���KI���#�_C���Q}A��Q̹�r�I�l��^�d��]��eP���ȩv�Oy��zd˄��7X�t���������l^��s^���F�g~bH6�M�Hzi���3+���t�I�	�x�of�C(|݉����NF�%�L#�nt��M������
��B��-�{�i�Տ�7sX �sF����ďW�Zm��R(eN�{��|A,
E�iM8�[}b��'���K�b�UA3�KI���؃l�,B��\�z��)]����76��d}�^ZZgZ8��3������K�mW�����l^��G��}��_�������!�Q�G�����E�ϧ@��!!�	�K���Cs�~+�I!f���C�`
,j�-D�1��4�֙�u��x��|�m$�� �6�C]���̭�ƾ�"�k�����UR��s�����|�����~�	TS؜���9rk���m8k�����5�~l�M�j R���%�����=IX×���L���J����}�ɢ�ܵ�?�H���gk�;��|��� ��.�+�-�Ej�x���s�m�޾�4�YL�N*��sq9r����WD�w0>�=�Qw����\G����q�dׯ1�Ժ����^�S�5�����ޡe�j���P4�D:��٭�\�����y��jKcVb�[Ǹ��:U\r��A��_��Oo{`dp�f#�Eʛș��g��N���?�5-�2,���F�� �0{���O(y�|������d,��j����<�����f�}!�AIQ�)�Q������*Y
��ʗD���r�0fq�btR��TQ�ҩ>�����A�z}��g�{��b��9=�o���k�	nc�VZ�����ꜘ6��B�'�{V��7x7[�}��1�lY6���|��Q�q�H�z/��Q�����ܷ�������|w`�5���%{xQA�:šgf2�jэ3l��b̈́��s�y1�و�@��5?9�ZG��R������G��_��+䮬�K��֏����uI��fsO�pgM��*�f�)n��u���fĩ�LK��Y����'��w�H�(��q~"Q�b��/8m��:�/7�p��N�+%��&�b�xs�Ċa%ޱ��� )`©KJ��o�k�vb�Ø~��f�L��ֱpk���2�E��(!�1f� ��>(p�]$�0���h�(�w��=��n{`���!Խ���He��jŶ�"�i�Ұ����PEy�$��vs�-�V^3�����/]&��������7�Y̰*����W��B�Y3�������O<�AC��>TTA%.YN�e�ǲ��ap�ut�v�PK��S�d�C?�CG����r��4vY��I~��Ut�5�r=�tc�x��ݰ:
}|?�yҜ�v�q>�nm�7�i�K�0�k�ݯ����`�_���zmQS^{���"e�"��y7����GN���"�%��W�����6Ec���ڋ�����ĸ0��m��M����0�������\��Q3i�:4�7�;��fU��SH�9J�5�p�o������IzN'��Öz=fp�Q����N"=S	l��i�Zp��ٚ]s�MOZ���>z���^��b\�e+��*�H1zhu�?\d�|A���P���i�i_��F���1���b�9��0��د¡��K־�|A��R��c6��3�qi�S(�OT�Ah}R{�g��wʐZ�=�\��Y6���\�i��\�O�,��0o��/ɐR"�j��#�rD� ]B��~\V{�O���8w�)J���%�s�j�k<�
��,�_.9>0]*1���c ag�������I��_0�X+��+93��l9S�x��о�h�:�#�MccO ��3�E�<�L	���F [�'|�<�/�����zK.OKp�Xe����s%�ԭCY*�-n�,V|�<e&��N~Eȳ���TuU��!;0]ź��0�S�C�5��tլ����H$#�%Дrޞ�z,!!w`�5.IUd}*�TXi���K2Lu�zx5��y��e�8;|�wx��$�{���=���A�-D�g,���{��J��ٿ!\�xh��)۶|K�-[R�I0h&Aa���/�L�e%��{��tqs�r��,Z�|-$@�z.Y��?K� #�s2��ƀ|����黱o��A��`����w���0�5��3��f�s���󟺝vUH\sS/��yP��A�#'%�Կ\;e�#[
W��uQ���'w�\�㗍d�4̍Q�g���ce����CxY���PȘ��l�W�6�2���aߖ��5s$aq���Ƿ���?[�����׎�A[��RpO��Ϥ��\}�H��߆&��������{ޒ�`��٪\(�/�¾h��[E�#m��N٬C�s���{����-��G�@�Qp6Gf��\Ѹ�}�柢F�'AjuB�1j�0��!�~��j��&
�A�O�	<g�o{RmN@^;���[�fxh/�E�@���$�2�_���#i�?�4�hE7����4�ƐeS�	!�(�so�����;����P���'���qQ��^�$,��L�p�$��n��c�?�J�����v=)h���RI�4��e�c��o{�E���c0��o�9v �[1�֛�ʾ���*\����w���{�Z��g�Z4[�F���w�N�sq��p�(�YO�I���N�C�.����}���?����V�9Y�S���5+��!�K��5�\����j��؁|���ՠ7�>(�5��Ht��73�Ʉ��?W[�܃���z���ӓ�����{0����@ҜU#_��Ӭd���AN�U۟o�4������9�_r����;a����,	�%��KF�b^���F=j*.8 �Fȑ�h�Z�r� ������*�cc2..���~��M�ڬ�ʰϥ����]C�D���9ZOF,\�5�}#��x4%�%s�~A�4�T�������ݗ8����Q�x)Pz��ö�\�M`[<c��t�\6���^�vb�u`"/��o�?^�N�E����NP&c�:���'e��������L�:5���A������\�����.*��ws%1(��� 젢��/���V\����D�����B�
�LU�hc�Z����ƅ���wZ��Ղ�?,��"%$E��y��}P�m�ėul�2�`�� �q9L�|�wu_*L{�ج��xƤ�u���!�gP�lq?|�����/S;a&@٘��r�S� �Ի݋W�Vfִ�G<s�������#��S�\�Jr�ϥ� �%XVs�@d����c﹵��5#+՞��������6^�}FN�����z	��Ά)A��P������h���|Cl��?w���}DP2�^�?I��^���N����=,3q�Q�Q����օ���6^R���TJj��`]�ϟ��w��Q�۸�2�ɢ�ھ �Y
�ܬCߖ!շ��@.�/9�(
ro�S[le@t����>�"�ogSrs�w�� @���x�͵�MR$�#��dJ�*�����5R+�9��h�۰~L$kDH�݁�}�^�����f��lC��K1�}�5���'�ݾCL��̎�=��*[A���_M�{��IA��S��O�h��3�ŷس`7ށ���v�����T$��]��?ӫȜ�����{��F�R��;��4��cT�Qrm#�5���L$ |��|�A���E�_/_~j&xٔ�g�|sR��)7��X$f����'G�� e�Ae(uX2<�A7�Wz"*8%�~0�/M��VW"W0��߇�FO0�(�+��;��4�����.џ!�Q���}'^�)�T'�ք XdSM-W�Jhe�+��	�$J�y�GQJ*s�-��b�������@Nwp��]R���z���Atk��=��>�����m���6-��0�ʢM�w�t�O͖;1C�����FZ�A@���	H&�"9��{��3���Ҹ�����Cn�"'M=���e8�;�%��M�,�2��
u� '�k��b���op�S��ڑ���ڮ�V1�;o�88���/ݚ��#�%�� �l��!�
�;�؛U
HЛ�(Ieb$�r
6",8�aX��¤�:-s1���=	ٗ`ש3�ڡ�*v����j0�Y�����fG��g�,��';D���q��i\��y�,���Z|����3�{o��' �.T� ���S������b���2�te�gج'^*���fiD LLT�7Y�1G�:׭.����s�/�{.���=J�j��#�W_�������y�X��ӛ���K�	[��%7���B$�n��2<7��L�@�Ie�?{�#�*$T��_b/"���"�I�`��lń�H�s�Hz��S�~�.	����yN�ś���v�J K\�[��.��0ܰ��3av���U&o�PNƝJ��dk~I��]�*��7R{^�BR.�2���&l!���[~]e۶{9�0���ٳ�^h�?̴D(�1�&�"�W�{�m,��<�yް{ԁ%˪�dl^2�x
_�TN*JMk8�*����O��m��I�r2�`��y��Z������}��M;z�BJq�xGƈ����� �ث��ZO(��,�NPZ^� ��fi�˫w����ݿǈ�;�YT��C'���-��YIM��5�TPb�\�������~"�t1J���N�A�zEZ轆T��e��
���5�����`T0+3+�|:r����D�#]Lu*�ڳ�o��@sF.��
߭�P��F�xa�����c��No��01j~��k��6�#Xa�/� !1�;�w{1]I@�B�Nh����ްw�ڪ��r��>�g�k��MI6����)�k`�'���qu��^?*�����+���sR?:� ���x4:r4��>�������|���~���v1�2B]7�f�ۋs
ĕ�j�p���c�1��Z���$��]��w6[���q��{��L�2Y �)>7���2�h���m���]�\m�؂&��5ve �L���i�]����$��XS�w��O;BlLI�-7�D�8�s�fL��+  |��!q�KJ�����r��:�_�F{&�1�m���,���x*��ՂX1+�~]t�#���=SW���5�sUsT�Qn'������`�H�SBӌ�*�,N��o��#�6#��vfS��[h�!���f_�$៮ۘ��ʐp�"�7n]\p�)NI�����]�:�d��]�C����y:��L����i�sY���N�n,�S���޲w5;S]�"��1���V/�%���T���:�i���|K{go��|�G�$�E��]`�=DD ����m�5j����o�Z=�n�YF4��"��F߾1�����#s2�G6��Hl��c:���f�q��C�!f~u�1n�����PY.���b��[��(���A}��:?��BK�N^������*��*�u�K{���y��?����,�g�(+���`~��=�ݗ�B���d��if�5I�ɶ-�.=[b�E$J��}��	~U�}	/�����Mk�4G�K������/Φ٭-�(��-&x��b�F"���?"����)�4�QCK��O[~�jN1`d�I�z�m�Vk\b
�q�n�˸U����%���T�C��A���7'�������{���M���O�w�C���
�b�!�'_m��ա"" �
;k�>����J>�$k��1b/en��ղ���hE��B�lo¤��f��C�)��7Z6�A&%R.�?c��;�f�����m#G�*:Ѫ�4�+;9e?�O������$�&a�)-��Xz0OL�5MMrf�mwa��Owq=�a?Ir�69�
�>���
}
E8Я#���bg��C�..�t�cdz���tؾ�]C�Rr������\�h������?S�ǉaӧ!��[�>:>�`�x�%��Tm�����U�\�
��ެ�ŋ�}����%�v���.D����pV��ы@d��ۣ�L�G�p"���E�&�cb�DVv·O�j�6���6�F���z���]��W��_ˬ�?0'Д�e���,�ϑ�B�������4X�a]�Yh6l(��ݝ�j��y[����q�Aa<\YlZ���[��,UX��V^� 9�����"�u���z������7W����+��t�^䍱���n�	�F��/��� L@7�Y�t�W<J��HV�JC����?^&拺j"9H0�^�E�Tip�;P�Ӄ�TY ���qu~�~P�Q.r��n�� ���#0P��|�
���m��]ܧ�=�,�:�*�E���T7��xhn�'[�\{w�2y?\�"��*}�E�5����Hܒ��>[��`��1������ �ۇ ����� h#.:\�I�K姓���o� r���|C�zd,+lb�_"L,[���Zlo�mT$k���R�\y��	\ܢ1�~��E}�����^�]2��O�k�e�[�B"�5��]�,�K��`����b��$��r�a���%N��T������[#A0=>n;x���jֱ��5#w}k"X����SK������˵�P�[1y{����"�4zǷ�y"�K��"�"���#�^b�-w:-��&N�)U��q���\�I��IY�FV��� ����4n����*�C��O�<��g�;d�=KӉ�_'v	T���^:U�2�`�nuF�s`��g���%�%J5�Q�
ŵ~���_{���)y)�rQ]6 ���#Kg��Y���)]mv�<����f��/����]�F�X֣����g���u�A�E�2�4��?C'�vL����p��ݫ�˃,��w(v�R� Vf1J��W���q�=֤��Z�bc,Kly������{�1{g�K�:�#�;-1d$�-[�����_D��×V��U-�HC.ǏJ"����p2kl�*����w�������I�T �,�oR�I�.��� �]^^�tuqi}�t����Ԙf ^e�*�d�rξ>k:p��BK�����w�S�bS�D��'��-L q��m	LC��)����t
@�<��^E�� u�+p������m����iJ%����D�/0����-��8\�()�fv3?^�����u)�<L��{�.�lv&��a��Za��`�+Gm�irKw���I�Zm�7�z�D����s�)J;����|��
�m!�	Y�yd�Z���/�{���R3� H^'�A~��>�3'����M�8���W�b�U�B�����ҁrz9;���.�N��{���c�iA���B���~�DF����`7X��em��~��6�l?Ť�
�P����=��[�@u+���7o�o��OZO�i��}Z�~,jj����������Bv�a�g7 �UM~?R��Í��+3�I�x-V��^ߓ����N�zw�?0)�/�
p�>y+��*�J:Y��m���'ԙ4B�#;~o\�
��'��t.�ɋ�G-�*�GG�4�SƩߙ��f��ԌZ��m�[��we�׾�N� ���sD�rt��u��5:�A	H�d4Z�Y����^Wꯔ���g�W����OG)�rڟZ:���K��؛�|X�a� b>���a���]O�Zݡ��3E4��%R�<x	m8����jǘBh[�g�F�ܘ�(����JO�UKjQ��[�
9ٕc�����̢HB`��G� ���(�\1�����S�+�p��R�(���[�ꗫ�]Zb�;WM�>�+y,��F��PXNO&��j51��TG��m�d;vF͝�W|gx�j�#��Ĭ�����*��ض(�����[)�ݽhq��-�(��ݭP�i��A�p�}|I���3���k�5s���940���:�A=�
�LPh��!��4~�־������f�D��}CQr����Ɖ��������5�spSLDPS��׍�Q���vg!N�D��w�E�br��9J��̜����FW��U-�f�����:�c���SR%�hh��}�ǵi�Y���vΐȻ3������؝��_J�=��J��X��,/��qo��X�4��_O���0u9���4����!��X��%�������]�$����&�>~y�g �v��a��o �3]�~Ϡ��0G��鿄�f��lf�솼O�[����>�o����*NӇ|ѳ���oXN{�H8Ѭ�����;��p)*aE�_f��|��0Pw7���.2��VC�Ӿp@�A����y��M_���!̓��}���\�6nC�(�
s6l��3����&~���Z���]�[�k���!s�f������%���..��9�9��P�%$%���C���~<�N�kwU��꿥�����O���bJ%]!�
�S>3mZͿ�w%�!�m�v���D�5rz��?�����%��h�*"���Eu�����X��ܼ��Pj�w�v���B�`R1ymIg6R�U���g�]ۋ��*�'�"���PƷI��h��cK���+CIݵa ���'N$�ؐ��|���l{�������eI�@G'm\���p�~	2c^{x���m��W�4-���^��I�s�+@4**ʘ�ߟ���,�����ܜ��+'P[Ӭ����M%4���k8+���6�����5�7�M�i�X���T�ϓ9�p����P�:��4y�!��/v׵����]-6~!��S��eN!0-
F��M�F|.Qs�d����HSW��~���#�n� ���7�����ȑ���$�ϲ����`��=�G�O�y��������l/
���9'{`�;�$=�sHyۆ<so$;Է���uo�x��6���pL�FX155\gg��!J�aZ�,�D�/�XI))<>8h�k�ݎ���K��p �)5��������N7���q�OOI`B{����~=��xPPh�b>��,5�'��*����W(A�����>vU�w�}I�7s��c�:8��E:��I�1���(��'d\�?`n.,��sd<���t���+#��E$�6�e}��U/Ǐ�n�݆�XN��L7͍%��>rmb���C�h q*#��� 2��7;>��c�姰1V���eҾ�n	�Y7��G�먥�ȟ��H�Tl�gY�_�ʽe�d�F���L?�"\,��}�fܒ2t��$�hzm馂iu.�����17�΅����2<β�(��P
�S�ݯBg�?�cR���:�O�ܪ��G��0F��l9�Q�q����	��,`����)ן���3_��M��1�
�`����`О/����B��2e�!@Ƃ�f���Wv�*�*s?zA�/z��d�ؑ�ZI����OS�v�NY��9��ӆ~�*�ܒI[(����*6���W�X][���#_����|xv�:��A��
YWn�.A:9"zl�^l���w� ����|d��>�Sx(�0�ԇ���xޖ�~3`o���\l�u=�+F��O�㛇�)�b�Np�.h�s���8��e�I�Y������!ܛ=���S5�����e�J�fo�|��R�a��������#jz����dj��X�f�E2 D�lٶʤ����	!x��8�����ܓl��!��,vCYR� �%�B<�b����?z �IU&��sӞ=�{�k)m����6v*t�rA,cg����2	�����Y���r!THC�!;�ndG����
(4����;U�@��~v-���
��dÃ��#}��Zg��e�봷��I���]��O�!��=��L���<Ep'�T���>��Sꘚ�����3cK;�d�۱OO�>w�	J����~YA���'D c�xS���9&��b�t|sS'�W-������
�9^i����8Z���q�b��[�o$����w�WL�p����}SN$^55������9lc�>ļ��444h7�+�ܛ��aߺ�H7�Ub�Y�|}��VPW���.g-[J�ccR��$fs�W�i$��>7Wp	=w,(�~� �󖥹2��v8��^������O�}`r�f}����㬆���$$I_��F����>knZ��@~��J�h�e�K�Q�������++sv?{�@S�Wn�P�bQ��u��e"�5��'r5�x���\kC���U���d^�c\��v�j�_-L�3�'��yF��N�/���@!r�2�5��̕�N��fQG���C����#&H�"xL3�xW�Nq�FqNy�l�
m��Q�i���h�jɧ��I�B>�sG��x�$0�H���=�X��=�U�'��|ۃNW�n��R5Bũ��i���uj�J��k"<��r��}���"=����J2�xo��V��%?�Q�Y`�Ղ�����Y���X��O�u��)�
���%�G�����vu{k6�#��a$�V�����~ Wih�w�z j�z!Ǿ��ewp)���~���ɛ=�X�����	�����2��"�����W00�w!�w^�
�ܖJ=��q�ïŝu(�܈�S������ˊv��l0����6�;��u���n��H�!�3ؔ���6k�WD�����Q�É�[ �/T-�#���G�[�&����v�����(s����bGs:.�����u��%4�������=��.ˆA�o��6[������8ʜ��6��o��r��\�cZ#�';Eǔc�9���?��EVPp�h?�������',O!�Od0��o�GjL�v>�Tr�����Nvm�:��:�g���n+-*��v{�X��߇��,�1�pn:3�?��ؗ��A2,�Ԥ}h���Ex�;�q�U�er��j���0��)��$�r2z�$�Y����(1a�R���d�T���D&o�a���L��������G�I.������򪢧,���Zܒ~���zQ�����x���ϙ�8���,Ƅ!W�Hx����ń(dY�}8�Ј��JP�D�D1�<�a�yp�	��2dx!j��.�w�p�,�י�l����x�FSK5,��9	O��'��#�I��_/���e��Wg�ßףD�~�=S���Ɠ�@?��X=j���y��bũG����O�5�eM�O��9�q_c�͚+N�G]�ok��p�����2�-�`���^���<���m�B�"�8�u���B��naNE�D?g��1�K	䗿�[}c#�=�(.���TӞ x��O�g�B�h���4��8�x� I,�	pr	�uK��@c�ȟa����0�u�B��"�u7Q�
qִ�VC6��)����w��y����4��}������w�������V�"���Y�G�G�<Ȅ,�=��g�/�HJ�K�/�WT9�d�9yVm?12��6�'�Ԩ���[p<ck���4���(ҭ��M�w�͔�
H�#F�nH���	u�-\�RLɐow[�: mI��P�}�z���m��I����d�ĵ�i�_���\¦sF��-D�	ܚ��c!��rv��4�IYV6]�����sFQ�"�(ᔒT�V�<kOo(��_W�1>>~�neĀ)Ь 9e`<��|�W�D	v���2�h���p��v%�wU���`DUk�M�D�h<�M�ӳ�PQ�͠㚁��o�����M�=����Ίܡ��@�xX�Ιȩ�)M�.���n�IK�-TP9�o- F|N��@�)"��C7ۯq��:X^���E2�� ~�����M�����]|/"?/����Ɂh� ���v��`iͶ��&~�Q�=�u�&�:RMu�WT9v/hll<�i�+�?us?�����H��|�4�8����Ը�cW��U���a�[���e:�j kdD�?stA"��/B��i=u�m-Α/��=ߑ�_i�J�8_KI<����n?���]��J�㬁��F�T��K�Cֶ�ML=�&��,z��|�2瑫|�B�0�[��Z�5	�D�E���6̅�O�~���y��3U�}Y�޲V��A��	2�t�ʼ�1��5Y��d��������M��[&`��y���հ�ϱ2�Dx{�JTA���B�hY�<�D��J�D�w�W�����Ǹ��ٸUePd�0�Cw	U\��!�̉�bI��qK)�R�N�Tߩ�t&�O�9��a��^�N��QA�
�����D���B��R�g���mk�Kv�����*�	�٠�8�����a��8�BF��J5`oId�Ro]ƲF;Hd�m"���x�`=�[1_Й�q:ݧ�KDSo�E��.����?BZ����R�6���ޥ�^OS��}� ?�y��40W��4���3�R ��ο���y��:G�&6ÉJ'��ے1���<(<�l�H��5x!=�جqj[�|�DD`�j55�U;{�>|��\IJ�삼��f6 �V�%M��Ĥsj/x,�.A���@y%%LD�7ce��[��]&�Ͼ����)�@�D�~��3�˦wx�{4�d5o<l`:M]a��ïy'�4�rH_}�̶�w{:���T�^���뱗q�FE���ƞ�����7���r�+�k|7���WB=,���3��VkQ-~����XP`D�hx�5A��p�д+�B�z���p��~�m<���ؾ�+<^�%���A1f��`����1�N�Ԫ�+n)���bKI%1ײ��`'p]��V��	� ����%tzv� P�����akP;��Z��@�0����iIT��dV]®O���{��1 K�S���K��\@0rH�>_�io,�lz6a#)#���.ک#�������[��.7�(d��s�u6�N��f�Ղ���oм��4`q�]�@�L@�l+��q�M���[��}�����F 2�v�]C\l�i7C�?3'���8�9yn�iW_�@6�̺=1Ep���+S����;���y8��%�jZ�n�t&t���� �Z^�A4�J�%�&R���,��N$\k[�� $����'�q!ۺ�Y߁��¾t[�N��4e0�S�*�W���*��DO�c�����������]2�&?��&�=��|q������/�� ��E^*"o��3@PO˙�3�U����ΚٙmH��
��S	��a���nN�i��_>9�ȃ`��H��{ȱc����bn�ۦgjq�&]4���z�n���)C3s�ҏ�o3D��'�%���ץ��4���<��+�V�{
��@��U��Ox2���^<�YQ`�[�#���B��W��c�*NgEu2.���[ƀv�竌�X+���񷑴���p��6��)>A�1+зc�Z	Ҽ��w>8�Mfn���~J|��A?k�y�����!�r�|wOl�H�{�Lziƭ�f�hd㋾'�9�e镜F�W��6����c�f9���U=5�!p����뙿mB��$9���Hӿ[e����� /��kh�瞫�9Άb��4)��w�E��>��4������KN=x��o?St���PB�H��n��dNP�\�z�������:B����NvJ���6��Z��];А��9I����W�yh(l?k]h�ܩk*���W���uoU��T�AK�]*�����rbo�J�DZ�:�)���|� �0xl	�t�e-q��B����9>�D�h���b���.�v�p������Z�9�ie��Xg(����:��̛�����u��>%����e.�xW���ʱ�8$m���ĭ�S�`����[J�U�3@^�*�=Lݼ{4��Q�6��pӄ__��P퀆82U�3Vg2�Rާ�����U|IUf�vYu
5�kYFzIEN܇fʵc���̏׫���D&^�B�6k�Us����m:�.�����	!�>g�R���B.�� ��8 @j3C����7r��w�ǣ�fM�3/H�|��W]�����U$����x-�a�7lC��{1=��U�^�҅�H�^� T��[T)�a1|G��d|j����6?������T�畴��n�rԜ`mn�-3��*��rN��I���$珌Y-?l�3�_������C�d��M�7�i�]g6nȨ�������ؚbvqU��Q�W�"��/6��*M�8��OPD������/�v`O\`)��d�0��b\Z�������_��$@D�S��PC�
�U����&	�1&��	���8t=�	j^4k�4�*�,�����45z�ۊ�+�'~|L�Js��V�J�,\�?��U.�ci(�+ntUlf����U�n��U����;v����v��'j(��O�x��,�w���&ӵ���l��e	%8�uۋ�3�D�M]}�Ǭ_#".�c�i:FkѪP54��iya(��~�)T��n�ϣ0��_J�6�c���oL��eك�}��ڋ|�q$�>�b)��i�_M/��"�yP�๦��b���<s{來�T5�΅*����dt���w.��8\�������^��[O�S�IݿB��h2������m|����꿕 (]��w�K+1q)�^eR*!,c�+Hs��ѩY1C��>˩��<yjV���aK��YC46��>�׾-��K�\� **"4�_M~\���1>�ӥ�<�d\�Y�x���z��T����9�v���|"
�Eu�;mU�}�������T�a[Ð���S��}7e�W������L�#��Ⱥ�����	gX�0�� ��k=@����[�T��vj'�����m��jFZ�w�T��0���!n�Ő|nݑ��AP:) k��T6ߠa>?��>�B�����׎^���هaa��K�HIJ�E�RڼM�@�i�#]�2C�6�
�����S�|��btP�sh�O<�
�8QO��G)`G����Ap2w���P���eC����կr��v���H7;���X/�Q�$<>��,c�W@O�2=F��^���>�1��L�Ls�O�s���� �s{���-,����J��i��D�O����X���F}+6.������	�mNqم��\˘�����u�Qvȩ�J�R�$צ����5�������y� �grY�H����EQ嘑#  r��#���<��w�̊y�=1xi������o��
NB�5�mZ�f��vs3T9�ol,�t�n� ��{ό�i��엨��7ֶLd3ut���~�t9=#��N(o�,_TF��/���|*�v��d��r"_>��[۝�|��
���x��)�r�Se�8Q�ܓt�~o8t���Z)��t�o���m�lX�n��N? Νk���-~+�]��^F�N:e��OR;�nPQ� C���o����TO�F
4)<�&�(D#T�Z��R>������+�Jx�ss1�}K;�bx�R�ش8�0�)�3ᇇ6�B���y��yC�f����;�u7 d��C@ݑAey�^�0Y�)̱�鼕��+�����>���d����n�a�3���G�k)�ʒp_ӧ��܏~땲N$x�]vm;�]�	.0�T���}�ׂ�&�ei'�<<u�yI�������	����v��c��h�=	�-6��@��y{@�j���y'a�x�E��	�9Za%�v�
ڊ�O^�1�8<zNyu�2�u@�Y�C�=d{���d-Z��ۂ�p=�L@#�ʛ�����9
���X24�|�:��T<��1�4W,�D�6�Z�"�u������s��_5�8����@���?�etи}1[�l�Nؓ�E�I��m�;��}���F�}k�&=�8{z�ѺR��V�ك	!d�0B�C�n��+B����Ĩ�x��*iGn0NԜ���Y��3ES��h��e5F�#'E�p[���<ա����= ��9+󱼘h�TY��:Z�}ˡ��<䠴�D�-��b����0��v�ߣw����T���K�����Kr�P�T��3�����[�k��I�n>� 	����z\�(enPPb]}��os���8#%"d-�'A�s��k`�F}��j��7�o�.��n[ww��,,B�tØ������z��9�MZU/I����1�[�,O�ٙZXtNűs-�,����(-@'�I��ۭ��e����&�럩�i�cu�T8���,�R�&�vRˀ�|S2���߂p�ˤ0�I���h�4������a9���/HB���2��'9�����Ī٘�@� ��[�j��>9�M�f��F����	���0���-��e�2�5ڛ����i�R@��.B��b��7���-Ž�#��~�rwPG��X;������&�^�]�x����#oB�No�·E��`d4<�m�2!u�JFqG����[^�߃��^��1�>���Cz?J��'n6wjb����
�{��\o���f��9?����+��/`�#���܉���,��	�d�"�ڍ�ZKIq�M�4�>��%`�� ~��#/ext:%�k�K;=9tB�i�Z2���u���=�75(W=-�C���^�hE�<���G�������i�= xz�vVgO(���&ld���mr5s@
��h�F}��u�noi�������[����g�"�|f�)>�j��`�� ��͠}��qC�r���L��I_aSgڥ�7�N����iE��� � ��ĕ���zنuT�k�yzsgO��ÿ�0�j�xuF ���ZE`���jQSHL����Qu���e=�zب�p��h휋��*x(���:�>*�����صT�
��|�2v�[�q�&L�p����PdF�$�*F+�,x��뺃��1C_/���\Ќ�.J:G���!N�{�Cl���VIE���M�����
����L'�H��M�>�/��N�y5������+ݝ �˷��,P�6��{�z1)4o0]��>(H	]��cM�%8�{�|$������v�����*�ȇ$�Պ����`��6MK���OOC�|�4Y��Y���E���&O)R
�AT����S�g)�c�H�!џ�䶇R>:�vz|�o��y�9���|�4�})�4��ɢ�e�Ҙu*�	��<�3��u���9:},"]À�]���i#p�����0	j3֕��P5�MT�r's�rx�\I����UWb�oƽQ����"���I�dm�"q���hm��C(љ 0��fw� �R��'�ţ�ʛ9�Ѯ`�mʵrt����p�N���k�Y�$�]P�P4����4`��j�6m��L�� �ʭ�C��]j�y!�ԃ`1��E��Hy~0�g&IX�9�l�e��L� �\��56��rz�+�#�ޟ~���،I|��B)�(��&,Z�3i*�_'�dldKTu|�W��\�b?Ύ���ŉ��C��Q�'Ʋ8cu� ��c ,p�,^q ~XI!�z����m����{�����t9�^��X�t_Jk�ժ�kJ��e�����1[�p!�|'!������1�d tZZZ��3[{?�����i��۱�L�33�Pj�k������4�w1.�б�|d�o����	K�OVZ�Ԣ��ϻG�%�
Nײ�+��y;b�d'8���t�8�_�i��`���I$�5�̞��IWv�1�c�w��(��ӈ!P˵{r���^�ɳZln %mr�\9q�1����ˎ��& ��.XZ��]'�|���Wˁ��"�-W��
=/��u�D�O�� ���Z~��I�?h��ZB�7W�5aFя�E�~71��`PD��n�w��L[�+��FoAYu��u#�xmM�����=����n���pxo�'�G���wŊ3"L׻�,J�E�$��H1nnn@kj�㞵��g�;�O�/�ɷ���=�.f���+5�mřL���8<di����j�A�,���Ma�G�R�!X�����T���8�F���x21�޹�v�i!�R�e�Վ�GԠeZ�ԩ��:�tR�uWAX�|���Eķ֫��[�'+�l`��$Q6�/݁Д��&�Y�`ba��pe��I�G�Z��{)�>��{_�!"hHJ����\E�鱤�T~��r|#?ʬ0�����*�?�4O�����V�>�_��ފ\uD�S���E>���MB:��^Ao1��X;¡����ᓌ�;;�.�_QC��
F��7�����c'��z��(�XG���7�����h6��PƑ���`
=�?�;=�.N��Y�����M_t}�Y�җ���jlWv�mv�ﾝ��$���)d�+s�T�Ƶ�����-W�ȯB��2�}�����i�a�8�z��Zi췕�ܽяM,�8��ɼ��$��36Յ���e���� ߊ����Q��<��|�y	�n��;��lx�,��C�%@�ҁQ�B�o�~yUn؋�-2&����%��4�w�����9�F�6��o���'ϊ�|�D �,�=�M�SD<��'l�m��3�ޑ� EW��a�����߰��Iw�|�����6���Y�_2�Fm�ssm��q}��N��i�D�6��{9���=��A�wa�gK/k��Kі1��Sa���{�;�kx,ʡ��6���%���z8ijK�-~izK�Z����\b�?� �����稠��S�QXx�FN��~��OoKFS����HMG
�ֵ��OWI� S9��6��qL8�f�� D 9N�}��t-�Z���
��+ʧ�Ss�E?��{Eu�ҟ��¢Kqr��`�xG�i��	�6p;�rq|]�\�H�.V��������6Ez�)��˧�o�O��)U75ʊ��7�8Ԥ�HP���^��ik�b��;�ô����Ϻ�E�h�J�]K��I��Z���nV�op�r
R��X
�Xu����i�$�ơ5�s�t�V"�e���A�q'6|��Xʏ�G~��� [<�������iq����%C��ˆx^)��r�{��<�L\�Z�:��ysD���i��ew.��(^��0.��<h6�[M�w�}�6�K@�xx�J������<u�m�~���ژ9�zA���Eojz�q2e���P���Q�i��\
����r�q�;�����f���wZ� p�޺I$2!#�@\I��|Q����Ox6�/�Ѳ�TPi����JX� $l��|�a&���PTD)�iT�I9�	�@/+�Y>�!ٵ��]�vk���=IBC�	D��r�&���X�t��?^�/���z$�N8��MW�8"�E�.-A�X �-a�9��1�X�m���blY��k\|��������c�8�0k�#��b��׸v��^<�פ�����.{)����e��f�LHz~�i������M-kq�fʂy�)|iHAQ{�-���~����vRc"�r>�T� �6�����N��Iл7���\�:_���&rcph�-xq� �x���I�w2��訔īx�F��y�X���ɲ�H��e�]�Ʃ� 1��XWc����ʿ
V�hQ`R>}?_� �k�|����̃ē��l�M�Š��$��ް=o��KY����C�h�NJMM�v�5j�L�>�)h���=_�B�K������2V~`��5$q�8ē��7�>���ټ>ё��������M���(UH�0}^<�]04a��''�'wkV�]B9�f3I6Г���G҉U�WTOO��ʣ��o,�����#�v�;4;�:�����\�w�tE���a'_M�-������f,���;6:����F�(�2��4K��`��-Q6������P���-G4[����Lw&X)t|D�s~��4Ϋ��D��e�&�������,A��0��"�*�̽�� �~++{^N����qOFYIi�:����,$��=fNq�s�K�*���`#�t�̫$1�}��p�9��O.v�$�pȇ���a�^'r�{=�uH��I���髩C�w����6��$4�>����]W�����մ̞ +!��j������"w?�xĖ����z;��O�mXB��{�:;;M(��Չԑ�U�J��#V�j��Fٓ[�V��g�O�$=8��pϏ�H`�UT��j�Te�p�U���^쏆B7D�(E��i��m�H��Y���-�t��H�|�i�P�)ڌ]����^WM�չ��lS�L�wq�#""*���s31�5���'-���U>`5h걕|�$o �����OĽ�JRꆿ� �I�콄p5��p��\(��sگ�+���&�9� �a���T^i�0נ�B����Y!���͗��ݾ5O� �V�:@�J�@��s �U�����ag8�&q�mC[�R��8r��Wb))�g�)o+\~Q���@����},Q��)�"%9U�/&��_�B	 6cI�2�oL$�(n�/X��"5cE�o�:k�'r���U���H$i�5⪀Z㌞/RK**�j��'HK�������O���x�R��S�OB�^!���/(&�IW��r,�b�c��o�P�!��$�,��Fد,/̝,��=Ŀɶ�>��Ѹ���N=�
������:���J��>NħR�����b�kD�4�;�a(E�1ε�F̷��{ԩ�IEk&>� �\�`� �d��E/�ݾn����(
Ev!P���}J�/B��x&/�l��������r������&0.�#�2��	�?�rE4�_sA���e�1�Q����}>ǵ�ɶƟ���x��۪~ݶ��gv����Zm���d$H�LZ�������?�= ��?�i����������Qh�����;�ͫ��?;2^f �%f���M�G e�9��y>����\r����|ҕ�h��~�j4��I��á��U�K�:.P
�|qoL|C��8h�M�O�ni�r��[����ZT����^�i��IA#yZ�Ah�4��<��}ު��?E�_a���<DD0���K3*��%p$5��-�9EF�j��V2�� �+�����˽9w��F����ԣ��X|���V���Π���zm�AR e��D\���
T�$�|K�?~�:�}���u�?�@=��}���<7��:�Αn�i�o���O�Q���(��\+��0��g��`W��VF˥����^�UνFr�s�y[�A�r����@�W��)��Q���ܜ�`x����hKN˥:CYJ���pL��D=~y����O,�[�����$��90�%9Z�T������L�*���"�
����Qt�kW�t�8��;e�� n����{��n�J,�u�����h�|*IK�; ��)K&����ە����V��H�g
�B�]�����8����O�C&[S�2�C8Y���Ǳ³ l洣���K���w�1��kIwhjh�8D�D����*P���\｡�ݭfR�T�o��ӌ��S<���{���zZ[��A�X� ����+�f1͜�����t��$��K����5}7��sA�g
6�Yv~�g�#=�3P�&Ww����ܱ��d^}nj�X��mM�-fT�L ��f?m��-���3�.q��we�ߩ^wʙ�����s�7%`�7Z���?�̩�������=����h}7G@Z��T����i�.���������H���aH���u�g/z_N��zd�����Ȣ� p��B�x��TisDEK���d��c���P���F�ˊ���Z(E��ר���hR��V��L��-�MR�	��@��\_�B}�TX��JW��ޖB#����<�aGY�!��'D��Di������'�6}��D���1��˃	�dW�y�<츅�U�)V�_���+v�.9$����]�K_-�N�3�wfW�1|d �� ~mG�)��%y�#���9���֧�$�_#:�_׎�_�*9��	�c��L=9_��=����M�c��<蕺TKt��NכA<Y
9�
�n�2�m��/HQQ����_���.X�4��
���4�c�֡�T�c��D��gW�TTh�D�q��z�`�CaE[ΩZ7�!]g�m%��a?��&��i͜������w�1��ӮR��+ވ��W�6{��ET��M���?�ʠ_�b808�~vP��ʮ	�g��RYV��)D����>�O�VQ�pP���k�w_�S���V�=����]�(���0���+�
�*�;7�$7��)�cjIU�T�L�f���Ax>������i����V���/��]e�Wý����35J�Ϗĳ���T��{����|����=M�V$#������!4��hP�Kc�^喑��3?GG>P'��_�Q�*��&��T���.t�h8�~�H���<Z��98���ƾ!�m��7V\���V\��*xڕvjhPO�.��E�H��_d�lk�s�������CؑR�k�h�<�0���s��~l&�ػ�{����,q3�>�%GJ鞩9ic��p`eC��IgB���xû?{���J�\7�8l�����hj"��f�3��ʩ_ADDt�g��~H��� ��/rB���d4�y�tk͍!�8�u�`^�6�s]��wW�����A~�_�d�R��َ|d:���*̌��y@��54�P��A`���E����@�B?�����R�:˅������a2����G�n	�̟�؋'�O��4�u�=kzz�fEh����^AT�E�a=.9-6�L�4T�W�ױl�L��J�d��i�D�:0 kH|���y$!�����ǵZ�		J�{1��3�����_]����9R���)|��,N����;�\�6K�n�[�΀'���r�m�w��pX�t��#�!m���Н��X�}ڟ���|<���f����u���Y��sX�1D}�KB�Oj;�6�?����9UwQd��ԍ<m���H��ͥneJ��^�輙_���*�6���U��δw��JD@J�L��gs� F7.=���8n^���4A��~��o������Xg[�DM���3�X
iPc����8���!}6�3�Z>2)��&+�?��KP!��3w:������	��Im��?8.���r�������Ģ۷{BH�}�N��V�}�3���T��SW:�<.�⣖���h%�_����lh�pp���� �s�L?]N���u������2�-ŝ�R_F�ze~�g@���
�����
���
����(�C���M������?�$x|�
s��#D�G�h�}[���b��:"F���\%$���0�]��o��R)��2-3�D�Qu)�ӑ��]�xL���i���|��O{ 	�B�_-3����H�iAۯ{��^�9	�c[Oct�o��0[O�]�
���UUɚ� $f��1*ȊK�[^X�G��͛T����9O�}��W�ࠋ�^�4h�.D��7uZ=�#���L�����r�V�t�H'%�,tdy��!�k`�R������'���Ug����vpl��
1�Vq8
AcW�JB��g�~��Gr�	!�hq���Q��w+U[��f'`�Qϫ]|���:�,Y��R�|��A
�7j棈��CI~
��w���յ#t�w�L����/���(+�fѤųZ�����Dr	�n<�x!��3ß��!k�sqk��ww��v�p��+gǳF�:j���6p��u����A��dR]�y� ��:a�R�))93Ix���v�0���&�YV�*a!�:��y�v���-�ŎZĽ3~c�+)H"{�+��NU#������ֿ}[��l}ĴFL%	F�L�Gp��}������5����3���SOI(�^'{ꐃ�Dh��%ߋ�f�A��մ,F���կT� hD��{���J[U���9��.���_%P�:>>�����
خ��8e��1�mx�R��F��#��o��N�X��Y���_�����d,�7��EEt���dw��$������ڎ��k3�UK�V��*U&;'8�RqG*�]3�8_u��O���ھ�X��̅���>����E��y�SkV��1����G0���JSc7�j�7�JK{�o���b@!�i�{g�L�u�6���f5ڛ��j�����|�����#w�e�d�r� * µB/�_S����[���?��z}����5���q;ޝ����цbH��b�p��actbQ�6������cI��>�4w��)d�m}H7����2zd�r�����(�L���-c���R�s��Eo�0�=U4G�~��|Vtz'!W(�:�ޚR,[*���n��̨l~|%��rh���-�]7�}������Ur��7'�o��!*��珯�T0��?\iO�S;����K�\�6����T-�u��FWWw2��R�/��Y������i�Sc��OM�Y���)Q��F鳔�~��$U#"A{�<$�û��5��*�o��G�3:��m��{)�OQo�(q�Lj�GA�{	�<,���3�J�P�R�P
��+�a��"g�t�R�9F3�k`o���Ʀ�f���{[����P�����L%g�%�<�\����ׯֳ{�s����bTP:)j��))�8�ڕ�2��hY��yʣ7y�j@sW�\y���]���Q1i:н&��S���� �'��zu ��]�1��a�c�I:_�b�ϔAd���|-e�����6��@���@D73X77�b�x3�t~���L�[瞊#��g�ˇ��)ңuc��³oZ��@9�,_]�_ͬ]��ߜ����5U�`�O9��@��X\ӊ���o_R	VN�6ct���khDuy�H�[B��~� ��#v�����%�z������?��2��&��E�Kqk���n�+�^�H� Ńw����@���!@)�~��zY7k�#�{�̙}��3���ܜ������-999vY���Ո �!�܅S�,����խ�j���+��&�9>��%���>ˆtU���Иz̊��O%e�A���G��u��qr��q����Ą��YǀͿJ�L��N�I��P��Yo��!4p �V7>O�0Y����L����G�T�/B�ut��>��x����T12j��S}�_���v#���CQ+?�o�jis��xq��"��5�ٲ"*�y��~_���8J��P�l{}j�F܋����7  ��"��H���,ѫ��U�1L0�h�,���s�_���}h4�|��,�'�z�4�1���������]�x�o�@��n`i
�z$����tE���9�8GFP�a6�H�#�!k�ȍ��&��U�Q��-#�|;���c�'zL$���H[�ӡ�z d��r���0K�Z6����L�^f�FX!��6�5�,yqm�m�Pk��b�RL3�*bex88:N;K��}�%��f��A* 9R��;z0؊�^J~藇�
�b)!ԇH���)�<t�w��c��s$��X]-��q�Ҳ]�2w�B�&�7�=.i���|7a+=`�w�����s]��N�~��Z��C�"cN���,��\��0�}���"g*T��~�
zL�U��5[���ݦ�A"�Ɏ�1�J{q���ط�e`h�������I5)���A�iӭ�慵2K����t.׉$c�Gٻo�.rL}EM�����5�Q�g}>)��.���>�i��I�L�m�e�0O���^o���p�X�c��m1J���=�� �t����kl׵��r�n���1�k߃H:sz���)�(O]Vb��2�=H���)��Lyy�S�q��4������%�嬣�`��47ِl��8�Bos��l��+�l��3&wY ���0�]���;��ۻ/}Wÿ�S}�U�V��o��`WH�~�^a斏�r�^�9�f��U>LH\�>=7��k�N)V�YO�_|��C*"n�tp��z��P���S��/}�Kڰ�9�)8Tv��!̛EI��3b��~�j9�����R��/>
.6��
�y9�U�'�}���Zs�=\r8�������� 8�?_��į��hX����Flẟ]�n-��!��^)��UL���^��;q\#��p������ɒ������>�z�Pz4A�*�ʋ,�"̇'f�)�E\I���L�%+Y��唆�Q������KY����B�/ك{i����� ^�q���%m ��i��2#�+���� ��jԇ_[�����~(=|۱��|�Ic�T��yG�]�w�:������J��,�13�aD��=�W���R��O�bE^�<O«�7�[Q��9����}�����PϮ�8���^���k-����ãg�5��}�����"�蒙y(<	� �}�G�>�0��5�0WzM�p�'y�ϙ����h�%�J	hO��&��#V����f�d��������iI�	S�^�y'Z�����?+��4�����_6ś/5��7=�u_�krSt��Z��gp�����U9'��ؘV��R����jm��!v�Oq���?��n%�9�O=��*K����W���d����u:�>��8�m"E�p.�|���>/^L�륥�)ˋ��:J��Wj0��������i�_B�Jb+�ⷳz+F�H��C�h�-�qL�Д�����pz����=�/2usB%X�N�W�<��7 ����3o}�ɶ���˖����J���&�|N� �7����^ҞM�(c�@�7���
+ xJvv4����KI�}��BD�7'��1�����t� I�1�z�>7B�yZ�5�]�M=��k%i)F������{� ���xg�u�%��$���'�'�]���Gd��:����'�[/��ŷ~U��k:C�^f!3+/���:U�Ҕ�J�H-���t�
��ܙ8
x�phZam�Fn�����@*@�C` �ڑ������N�3�������If �V8wՆs��:��Qѝ���s�K)^����EE'~���l
��M%˯r�ح3T�*y�fڀ�%�g}�6>\kv���:JT��"�Vat��	���՜��8Q$b���6�K�M��^�vv��ZYE�4�s-,�s-3=�.W�p��	�����z�A���B\[��yGŉ0��==���	�X��AC~Ok��lx��}��"��[=�n�^�H��k)w#G$��#�V2:'`zn��맕h��r8�:j)��s<�4�E�M��:E��B��k��=��s�t��8�&T�ڌ{3�QCC;6�):nO<(XJ��L�S����>T&J�z���&=��c����	r��D�_��sg�zdܽ�b�s�����B%�d5�������ׯ�(�\�yo8-���j���C��.�2�73��י��\�~/r��EG�ՄY��p���{ E�ؾ�&K$����S�&m0-r�d`�(�~��]���=�|�ڭ�X2���:�y��T-���HXs���E��Y�>:7X���1	��#-=yE�ַb?
�oy�g��Á���]��G�Bƿͅ��Zs��r�/�o�tK��P���3'�=Wa){��6l�?����%6�#�Xρ���8)�9�zL/LV��:�� nkkK��`�ѫE�{�ǘgA+�vK�����$�����՝I<+�:Du�a�N��xRŀ�����bX��-���;=������L�����n6RN��p�K0T�ya����}�B��P:}��L��t��ai}?�`��	_�o�����ʛ���,���ǿ�!m\nK?��Ű����eT�mo�OX���m�u�sC�+!��K�˚&&�M�z	�۳S�z�=���ѽ��H�UF�f��*���x�Gc�����+�u��su�kݬ}^�	`�@�tf͓�����J����(m���M!X	�X�6f�冏����7H���R��$��4<�[B��^j-���<��s�-7gu�e���ٌ����0;WDM�ʥm���x����͒,I������;��l8�9�jcX�}��dz=��L�?�<uې�F�&W�n7��u�UB]:Ơ_���<:�Megfe���kF��2	j/+sɁ��p��O����A����z5ۊ�A1��1�n`'U�\^wX��Mka��G�=R+W���s,��	=
���F�*�����A*���6��� ����Ւ:��$��E|d?�aB{�@V�v��
$��l����$����:���+]�u��=df$%���ʭآ�uJ��� @�O68�Rʴx���`Nxꄾ�Ί|mgh�qW��	�/��z���urr*))�)xCY��K���A~1�HR�r��Q�&=��ʶu>K&"۽
��6�\�]���U�u�����������e��	���C��M4��bś���1�1��7%��Kz��	�Dy7k�"ZϞ���NW�=�V��䒳���)>�Ӊ,���a���F�O!��=#�IK������%�r=��W)�����w��r�KsQ�����	@�>Gs�5<_5�!�D�
��	���}z1F����uH�RPOW�b��P)E�\iҤ{�e�#YTN�A��w���?�b���ج�I�m񜽁�Oq��~Ͽ��.H���э�ǥiMR��էRV�4	RH���ħ1�n��I���J-��JN�kv�ǶvgZPӼⳍ�VJR*0&�'~bO���1�~�f�����%p�ӷy��䤯;��?�.�7�=%@�Z���N�	������� ӌ�F��,�%8��PE��r@��>y0o�����;��S�n��`���^�7�=��h�����ǿ�eCH�b��d�iʏ/�3���՗k?Z����$����Ж�&*M�.&~�ޟY+{EO��O4��β����G��$�jocђ����z���/]{.a�]AUS����|�o���q1���p&@����y��e!������q�u@�R֣$�ii��_|8���"F�|�7���C������<'�L���-`�x�I�����x�E�a2�	�6�G]��'3}15�U�c5���1y��ȏ���A�6���D�~�l"^��wQ+<�7����۠�؁�eu`��O(q9�������c��wr��.�:[�L��[�f�Z ��KܝG����\G�KN&<|�ByM�H�c˷m�x;��뭩M2]qn�Y��������z�U�Χ�o-@�b�f�(2IJ�T&��l�ʘL�ǋT'���U��ә��-Ԝ�̷���gG7�*��,3Q0-:3ۀ�D8��j��~�"�~��Ւq����>���֋F�i�6����Z����6��;�c�+�>�ؖ��ן��|a<��kL�61,}�]bo6�A?�J�_�wwQ%u_P�9v��=Ν�mn�];���X����/{���5���r6�2W~��e� p}y�1&�����8�$/��*O���
��A��C-K��q��_��.B����fصˀ�@��{�.5{������:{�Dy/\�p �0z�U~FYۅ_6@�"#O�S���������εQ��ǽ�0��֚iս8Yz>Nx�}Y�b7��w��KБ-��%��`pH�:kT���-*��T�����FJ/�)�_�4����h�$Ķ<����aI�������C�h@�h��a��������kM��F*%j`�[^�TR�j]P^��N'^�/`�ꓻ��eޟ�'Ut/�ۈ���iҬKh�B��:��~��6���P��w:ӘnG�ge�b^t	���J��縒	h��kv�%;�x���r}�G����g��W�8��M�Y�Ҟ�
��f�j_=x���C��T�L;ֵ�T�2�����Ĕ�Z�Y"�E�v���+5����v>̬�6*�Gގ��Ș��Lg��[Yh_ &դmU��D��ƼK�/���U���"�z��[1e% ��~F�U4.�}ꉼ��]���lI�����{��#q���I_�ɒH��������4$h���#�{/�N����D����aΫu8s[��
��D$����q����᛿&|�9����h^�X�jQ_���D��a��0础�����o����V5LɎ��� 
���ޝ��wAG�7��M�ȥ���C��X,�.����#?���Xݲp$q��n��ͧq�����C4��e�!�[�]�������?<P!-7?<�J]��.�ǖ�ݐ�G�X��N���G$�i�����(�,y�k8��YQQ,�۷|?Jk+���<��ֱ��U�W�
����z�τ��cî7���~ �5IS�����ፎ�ވ�б�y 
��,�	5�Q4�4uuÝ*_S�Z}"�/�e58���ǲ�l1�_�s i%�2^ಋR��P��	��[>]_����bd�W_4�F��܀��������P�6�ǆv �� ��\�=!�R�����1�c�8�Z�R�(prWj����r|�@�v,�}Q�,B:�����܂�'�5LFd]qq >>��fZz���>	}B�{"t�x��P�943��i7�($, ���c�ET*�f��lAo"���+�8|��dan����w41���{��?��,7�֋vL��$۱��ٮ`�Z�!����_D��|�|^�����wHƲ���#&�5n�|.D��:Q궷$tt�Q�9��H
���E�_'�:�T^SFi�;�/�h]���P��X:7�M�dA�Rz�w�9o�(�������cf��B ��!��N�M--d���;p�ɭJ��h?�:����|Jªy;�(3G������Ǉ�S9k&��:�F��/�j�{&k{�.q�O]�� �׶e�D��=}xS��{v����A*C�"�>
T.LE:�,=�����m��_�0�ߎ%f�^���(w�i����d�>��JxǠ�^w&�38��k��7DY��j����GS�����P�<���׬ ���(�n4�Ø���хt�~j������)�9���#A�}_� ��/..6�%'K�ɯ\��J8��%���t�<�CJq�
��g���	z@e���ëG�'��a��D��T
�ɷ��c0܁�"��3z�O��]��8�1�|�jvr����F.R��^Z��W�*+)�u~?�HMNc�T�֕���z�o�pU'��cT:�-.�U���,�t���DC��S��u� ���D��DK��く?��ȍ���sXLxxI�j�NZ�8�'uv1kq��SQ��-���s�ZL2m����G��tJ_H�0Yϝa�{��?G���j�R�J�e�L��U���/������!Kp�o�G޹��qR+�M�i�����#���8V<�A��}�=�n���i�9==y��|��4-:Rߦ�{�v�TT��jj �3q"��6�?jd�<yoG��d�z��&=��$��<��*�;�c'�!:�-
V��0�El)%��Q*@�W���5L�2�6̷�D��g�<��,��ń��H�T({Wy�{�BWT��`̒���Sk8��������t��a�˪���0u#s��i�a�N��Yr�Rb�=�>3����E�����c�~3G�U!���Q�zq�g}� ������_^�p�6Y��r�@6Q��d�q�:��D��l�Ǐ1�uB�Cl�	5@+_x��Ϻ�⬖��o�Z!���9����,�a-;�`9U��� �|�V'�Ӈ�.d:v���H�*)�J�\���`$ �f�~��B���>	�h0�Yc�S!J?ճ�U/�$��C���%q���ܷ}^S/��-����4'�=�����w��SM�VRH��F� V��wU�*ӹ7!C�f�Eyyy���R[ �o�dh}�\��(O���d���JFEE2M��u��x�W��ӡ���|�{�ulB9j-FU�	1k5a4�x�C�s����]���ķ��W�0M�l�G�.x�'�o@q�g�o�D�X+ y�i8�E�:��G�����Lׯ��jO&c*xM� �3�[���~"k�d�	W�mU�\��ŋ�]�i�}�}ݶ�t��9~��%�/G��o��c�����q����)SӮ�=&�P`�H{��H�`Z��v����魯L�ws�;���bU�e���I����x����I�\NK|����*�`�D�L��5t����~�ƈ���{fz�( ;�Z�r�R�(H��yρ���h���N^f�u[��'��)��.U�wW'����[�]�[�����S�]�;mgH��F,��(~]H�����ń�F>������A8.� N�#3t����(d�z�E쇶�M�N/�z[�W�tY�����U\��pv6ݐ�M6��Qt6��2�tUڏ��F{��e@*-:\}h�x�@��0�� Kj��1�0���ڑ��v].�cȫ�@@������<^�m����痗�$��jm~�k��YnD~�9��7[�}�ϡ� �-����k���@Bu`R,s�F�]�~����5��uG�[���4��c�c8I[=�rA�r��M(��=����b�E/[N����������z��z=S�S�����,Α�7�a4!>�#��]LC�Vq+z�ϵ#���_��L�֖IDDd��.�$n����>�zD�?~oױ��#��L��B�Mv�իv���ko���#�r&郈���	P6GZ��|	�!1��߬Ow������FCS�" ^�ffB_���7�<�ɕB�D�#���O�h0��&��vVjX�ێbG����]���x����	;����KnES�	�$��ǽ`T�:��S���O[��dO��p6ǻ]z\�"yI�z������z�Ĳֵg'��$�w-�V�v���@ƣq�f�נݑV���<>:���Z���PE0�L�=OS(��98N�ˁP�xQ�f$??���R�����D��T��dɠ��!5�]N8�8��򀇿ry�LO%������`9wr����\�zh����d _Ӥ�+᭕F/���ё���D��v"y��3�,�f58�W��N���;�h�����+��旌U:F��t~YYd��7�-�{�l� �,8�	W0���'��.ٺ�4B�����ao`�I�#�$N襉�����������Q�$�w����2�]��UG�����J���ߙ,_Hză܄(ŷ��8[U�a�]�F�*�#T���f�S_	�\i�2K������_ބ�j����L��֭�,`Awaaa-���5��2�s��ß�iwצ���l�Ƽ��\�͍{�0�Xj�{�;�0]P�|N-�>���q����f�Tx_5T�X=�41�JN5(	�^yQ��hִ��V2�w�d<*5����M�xC�'�Bx�ĩǲZ@�e&����~G���8�p`T;��3G;��9/���0�d��nZL�9G�V��ʓ�J�A��D$ͅYj�E������X��>�=2��u�������eRwZp]��3R_�)�}RoIp\�����cC�"���0s�9\����%�L�����^ù�S`����c�����^Eѫ�_j�˓�R�|������LNM!����afnn�ҲQ��"�$�����:�#�eI6�"�����$C;O��?;#����vf��S a��cN�bcȩ��<���g}v� ��e���H�-���i��o�RP?: ��cuՄ�T��P�&7�I�_����;��w�������_�����QAAw��"|nVA���_z�O�m��}�MX~b��?��Xlm�3�Q��f��@�f�����ڙ�C�Y.�&��ϙ	}�뚘_[#�Kn�Cv./���]��!�^.���@��{�T���	C�n%�@~��!��,#����7�^�+y�y�A���$��سâ�KL{������vw�i�5{c���8A��������6��i��n�Qd)��ׯ��
igg'%+��ٟ�9[�vB�n�I@��k�TS�}����!/_��e�K������������K�<i��<��ކ��ۧ�^N�͑�d�,������S�l&�^���UY����IG�'΀������᭻�8قrX��Ͻ�a��3��v���zJ#h���Y
 o��ۇ���S&�'7�'�#I����8�
m�fQ{���ur(��8=Y{0���}���U�x�W)����f�e�T�)���מ�'��.O�O��A���x�<Zt�������*L���I9�_��v/�l�PKk"-��k��2�PH�4�����)lJ�.�!�����#ѳ{���D�+Rxlc����Cw�W7.K�������j�P�?���Q�O]�O���.+>�
:�9Pmy���TЛ�����Qҋ+�a�mIV��Nz�;�X�M؝���;��g�Q��(�5�e+�'7���N��W�k�D�=��Ֆ�Ӆ ~��L?��Z�Ԝh��b�w�!+����yM)�^IM���h�P��G�o��Ũ��"H	�O��ʊ�-ӊ�%�v+�ı��m��T'��\1����"�m����.T��ښ���������e]��"Ae.lq�g���5��0���)�o[��Ë.�f߽NzΣ��!��.G	��%�D{��,;�u}:�^�V|�F�g#�(����֓u�#�Nx���	1������jo;sԤ��K�}dI�i�G�������9Ȱfw�4�V�Y��~O�	b��F�_����\oy��j���G���E������F����+�����Y
C���	F5�����8�џ��Q3 KTIc{4b��c�F��Qp&���?��M� ��=���*��b!�\���H6�n�ֱh��`jU���j�s��j {Nx��`7ٍ��v�̜ڸ-�:[�O+�3�W�F�<zQ��`�����M8�l�!��F�/�"�U�3Ѻ�'�n��DFGg�m�H����h���@P(B�d�s^h�xI�������k��t�m'�p@�d�>��y�細���a(��o�Y�IP����5�2�@�ݡ%�����]���Ã��in��G����+�iՕ���s��͔t�b�Fk����L7�ˀ�Ņ��\�;38vn2u�.�g���䱝::�:n���P���mM�.E�L�T�2F�ؼ;M�G�����E�7u�:�K���[?퀜o�aO��R@�%�gDoB����fdﹺ���fu5����xh���h�'^�9懶o6%Ya	Rrr�v�B�q��/Dۏ9�,̘���kĪ��/U���\ۚ;�z��Gh�[-���j��i����N]	�`�d���`!0���̮��<�`"U��))���)W�|X�`�꣐K6j�*��'�
�߆�a�Xb��Ҕ����hf�\!Gp����{:_\�wϏ��6ٔ�
*(���s���l�}b�GGG�6c�n�c�y����~>?���A��C��a����Im��s����`����'���|wp�a�p�`�8F��/Mḭ�w귏����0�揪���>����ĥk�7vZL��ƞ=N�cU�Z��s����& 'fU�M�;�q
Vx]'��>z�r]�M�g�u��;��LkgH/�pUz����1�,�D)��3wK ��D!i��^=�B����6�ۨ4��P{��Aā����n+��!s��	�y��!���mn\G���Ö���ˎ���rT,o��$,�O��h�u��s[W���((8�0��5���M�,�������;-��1
ʀKvI�^Q�i;�j!7�� �`R�����r���w����	Uɳ���di���1���-�(2���,�[�Ӹ�a�帷Ʌ�`��6R��?���DƸt�K��v��;�$q�]w[��wS�O�#�D��fA~���N~��8
b{׻�,��}�O֋NW����W�t��)���SI����r^���3�s@����^-l�ʠ*k���m����g��E�<=Gq�Ns�_�w�JB��N���n��Q\��Q���DHI�U�椽r��<��2xm#����W7rZaOq���c��,d��zP�Z؉o͠�t�Sm�$mT��QQֶJ3w����T�CO߽���
̮�\�Y|�U������X��L���e+�rE�[�K��ct���;IUPB�%x�je�p���KA#�|��+S(?������@�&*�v��'4<���s�/�֓x\��!�r�����Q{�g۫��������n�����΁���)���¨�4k���+�\ÕP�nmP��WTL���82.̉5L��y9�g;�F+������y��P�O�LZ��>w���4�-~�+�pT��vV���#p|��gMO�	�F{�
��ee`�B#�T�Pϗ�C]�Ly��KX�������>|�T���竩�U��N��f�$�h�\�A��WS��g�=�cZ�?ʜL�Gi��!�����k
�,쇛����~������)2���t�l`si.�D3b��&�_#ƛ[2��OE=N���{c��oh�wr4�zq���k �>��c��q%�����p��w�vz3�����t��~w��zdŁR�T ?���{pg�>�)�+X�c"��fX��k��j�z��k�
�ƶ`аQ�u��6��`滜���Q����r|��>CSQ���O��U4PՁ�0��k�����*&�*ƒ"
sTߤ�h�Q+!���̌�4�ݚ8�*Uqi
Yj�R�ʁvJ(A[	� v��X�`M���rd��+���2J�E���/�X��'9�o}�3$Mj
��Z��բb�<��T����uX�o{D�a�r���n�w��![#I]6��x]T�k����	���u��*����>��v��t��p1�+V_�a���4��:[Zx�ʫ��U�
���>5wע��+������/9Y� ,roN�-��4��A���p	m�FC��}w�q��	5�m�.�i���J����.�����D��<*�}yAy�[qc'��%3mc*�Ab�d��2�`;�}�x�z�
�^+r�\|�������	��He�4߯�YTK0Ӈ�ʚ���A���ѺD�6��n~�����n�宝b,n�Ӥۇs��E2�h��\(�OXU�!$|�-��S���o-D�
	�U4&4&�r�u��wI^n,"΢,ᭉ��~�1�@�B=�*�|�Nf����n�yT*��N��8w�[s���7��J�uT�&"�z�Uv�ڟ7ב�������"y���)��o- �i� ���ea�������zN�N�h��
i� �$1���[C�R�!o��4Vҳ?�E
�c�(3�Vf����	;]��0A���&�9s'4O�!�����rv�|kJ�C]�#y���bɛ(�TQ��d�l1w��x�CwC��=��O�U5��el}~7�Ғ���O��X�#qw�I�Q~��"��ԗ���F��3>�_lt��a��7��[(�C�<������9E���;�I�5���+R}A�eܑ��7Dz����0�o}�Ő<�2Ö�.NӔW��L)Тkʱ6�����	\���)��T*g+N���$ +E���g��y�~8���۩������\u9ט�"�M�29��f�����#�1����u�Q��4u������]�։�5��7GL��O%��{��i�yȹު�n�b5�x>?�~f2�Zx`��ɠVA���p��ޅ��ǿ�2�J_Km�T`��@`�f�ME%v�� q*�o��&o�i�5cG����~J�  dB��l��yιێ�C< %�,:�5}E���Y��=ӬI��8}���l�;�l��ÊP�J9u���^�u����[�X#�C�%�E����1��%�u���L����{�~���S" �?��}W����~�&:���G^Ib:՝G꫍EU³��B81}��l?E�T�\�qj|�E��y�Yˏ�u٥R���	��y̞��V�r�m��}.#x���u9�]���i\�Mr���=��r�y�c��iF��.� �.S���?-���^���՜���<�Q�\ÙPR��^��Q��_�p�?�P�IɆ'P��/��赱(�
>y���[T'VNK�7&����	?����J�0:~Y�����*t�@=�V*պ�3��
2�/��%�1�P���[����oZ|��%�M��xh�̫��uhW��'��8��//ӄ��=��"K@�Q�u�1h%b"���m+Qlh�~n�����tӊ]��׵�>���&�Q�>|�z��6�=�c��C�F��ݻ�,�F�R��:"�-<Lw�,����T����7nf���������1Hi1�H.o#���8p�):>�~%lK��~�o�Ĵ;���S7g�g���Q�m|���HDDT�0���D��(���Q��۴��zp�˳��OwZDˠv��<�����+����r��ܼ����o�K��'ojۉ�]�F�	<�v>�r�&��t��4��,5
%�2nk���ދY�ap̤�鑑Ǘ�3Uغt������_/��~lک	��9)�ʟO�`=Ƕ��؞�T���Ĺf�:}�i�˔���̮}�lrl�$[�K�Žj� [�_�����>I�ژw�1�X����j ~�M�B��*����F��2�sF��;�,��/�E�5ń��\�h҉3 ��;������ U7�gp.�#���mM��s�v�>��@���rt㚡��B��Şm@V`��T	%�� �&6	��Vc8����ԕ\ߕ�@��ӎ0��M>m��eeJ�lQs�ݹP�S:��2?�s���9SY�ֱ*h)�Z��'B��ǳutZV���[ӥwVR�Ԓ��+T��ߵ;-vS���2M3���~IΫ�-�a�/�N�����W0DX����6�y�3�obs -
���/l�2?Ф��j/�0�<��fx�MYW8��@V���D陵�h��I�{����4��_֙&� @�,���f������?���3z�	{92������#+s^���hl�;�s%�)k$�6GV�t(0��H��;p�����t%۬�<]�c��t��a&E��FNx�L���S�l�@倽3B�jln^�ꢏ�x�~�p]�&����LV�X��$*Ѕ"D�*'\QݠY�����|��.<��^r�O-³� A���
g���o�ӛkN[gH�5׍��z�b��'C���+��>��Rw6��	��o��`�6G=���Bq;����m�W����M��g[E�$�3[-r�6�j��1�R����c\��bV��HVo|��� �(�3_���|<	�'�O���0sln/�w����RA6�r���"q4����'r�K���`Bg�H0�{�yW���~��T�	�[�c����U\����̯1�g;�1X+A+X��)̯S=��pg��eb�ڭȮ��	�#v ��i���c��$v,�3Y�u�u<E�ӡ���ɢI�9��௪����K�_�Qb��G�5V��=[#d�K8������4-BS����=Р�E=�Y��kQ^�]v{K Cx����ڊR��ƴ��Wr��XZ#Knr?��*V�O���C�Cg+w>,iG7:s�{̆�c���{���N��h�l${�0"C�z�PBU1zK�+qH�� ǚ'f��E_�6V}�Ǵe�B��Ԓs�Es��H����l�9?O.���s\��	ݩ�^n�������� k9UO��a=�+���<�r�F�~��!�:����BT���۰=���ڢ�O����)�ʖ[{�L�&��h�f�e�"��l����XZm�����G�Ɵ�I.�j�JV�}\@�W��+u��"YU�pp����$�'\*4��D���ǀ8�X��~x�P�/}��\��ULh���!��v�A���U��:��+�ov=�>4�7`2$Mԟ�@]���Ixf��H{'3S&�r��&��`D�D!9�\�?��iFEwzya��#�գ�0Y�gr�>���1�0�'P�Jp{;�����HE�gz趍��"n������|��������I��^v�����7^����`ƛ��jnTH�r=��ҿ؞�Rmm�ɛ%*�����1،+��$
bw�U��F���5�� c���:��lP�L�k�4�6�jY����)7�e�?�M���\����lh�n���%~�rDY�{6Ѱ�aӓǺЍZ�iD"�WϬ��rC���K��0Y)Hʠ�	I['��v�(�h�������W�Nc�LuQ��KCN������Wa��?���W@"×����c�qt��C8���<�/ҾMW�~3��?UȆ����$�|6�<x>m��Ԕ�œֶ��R2��`H���?7+����4���Ͼa7���=7|ʻf��tD����?�g��[!�i��+���GK�}U��2������EN ��}_�mq�x$�3)N�쫶�4�Wp�Ԕ��|�8����s��_\V������Mh��:7��e�i���R��]a���p?� ��٨n�%�-��r�uF��UҸ����*�a/����	�����6�$�_vKM��+��Hq)t���-VwX�X&k�%y�%ʶ@Q���)�>�Ģ���O�Qo�8�k�{�Eг��#�Rl��ʞn����eK�-5<G*��,%��'ߎ|�G�k�_��=6 ��mOP��gs��wӡ�d���Ȱ�Q�#X���Er�I��:���u1+�p��)��틝�����Yq�m��?8���STm����L�ǰZ��0�	as�-��:�*��wl"#���`�������7��u��a�,��0�*��h�1JA��b/V]�z�y��?,n�-��T	{��
4�+/j�s�3����c���w=�jc�ܥ�!�paH������3���ؾ��g��bUKY"#������!iA�	W�T�����z�Uu��^6��GZ�Ť"���.��������;�qT�(Q��g[���3E�ɱ���*���H@�*#E��UhF�/��R�A�5���s��Y ��(��ٰ2����/�w��͟�Z���� >�x������\�	/��ã	�/pR-C:��[�~|HsZq��Q��׽;��+�f��4���C����ړc`����Ǽ��� .<�h�kI"ܢ%1�����{*<\�ň~ �ӑ��\�����\��X������륙;�1���0�ls2q�c�E)�E�����-���5w%`٘�?@�7A�MEP���z� ����m�s�S�W��	o����p�Tk"HM^�=5�o����c�}�iS;6<3��j"_e{�I'���p�H����"�@�k��>���ګ����7M a�;��?�u�PC�QBzc(�K�"�(�eo򋦓؍dPӂ1�����q���Wժ�gn9A�j7�~��8:��Ӏ���A��w~1��ׁ�4���7�ՂE�B�#>��C��MZhf>��,��td]]]n9(����o����3����#M�F9���˃e���gx8�D�aH@���\�kjhk�σ&\0�%�X*i�h��5��Î���3Î�!�)��U�A�؏&�dea�zxT�pL吻\�vw��S����:]�5s]��R��;����x�T<�F��ٺ���aM8�20�$�|_M������
�8���E��;�{p�A����/n���w��%����;o���_�7��U;�3����sϹ��>���e4�j����'~�B���Fn�J;���~��7~~x��1_��)ݿ�,���u� ��9DY��z�o�/W ���ǘ=����X�{��J�]V��zm1�&9c�����q�2���6���hu�'���5�H�4�D�A���S����pm����k�\˺22�67ۙ9���ދg�,�ȕ0�ׯ���Zkh��P3�a/����[����Ɯ�6��bR  #�U�.C#hJ��>>��<=��Mq����a��CY����2��`��d287u�WZ��`��M�z������B��I��kX5ECW"Yl�
T>�c�=�}3�'(0���sy�����:r�9���
�w��g@�p|5��r�@B��c�ۉ��|1[鿍�O)�Ϻ���(����ۿ�S���L����KF#G�Y�����߿�jY�ۀզY���m��yC�I�~����\�^J��_��|�f+P�k�|���0b����n)"��Л���g���{ܧ�����%Iu��vY$�b5��,i+='	��ɞ�	�3`id��To$9^�y��W��ŕ��تx_Ay463��V���G����Ҥ5j]W)���o"IL�RQ��}p0��Z��*�;oZ�FNMF3�\.�b�0��WM��,$���]̧��ƝVL������&AEl���1��b)���h�/���7t�N�H�xq��B���tt�>-�wL� ���">�l�׆�į�L ��E�!>��8�^�0)y٭O���[\��n+ТЛ�{i~����n���=%���+�4�EQ���q�"����x4�r�g�	걽��2��,D��q�W7�x���>�r���w���z���ytYNIp�i�M\6�k��m{��CY%X����4 �K�!'n[�=�dYS7�j�@��G��.)����hc׺ ��狙�H��,������(�����8a��tSǉa�ђ��8�'�|�� ;vX�8�&2"fѿ�7�Nj���ҙ�cc
Q�����tH2�Ш܈��W�:��O];?���j\�$��v�pʅ^�0KX��&�o��X#�z�1Y?����z�un~^9tۜ;l��s�}�7~6�%�j#���U ���QN+d!akQL�1Yߺ����Re�?;����<�tsV��LC������+���f��4ٕ�kq��3X*;���0;/�]H;c'�������5�:�X\`�r�4�x�5�TuøWd?�����ĕ^��ej�L�i�������v���>op���Pb[��e�U�dw�2uZ�;�ڨ�վ��v4��,��IGt$�\.�8	e��W�[�Ⱥ�J��1?����5���G2f4��Fnh
��k���M�x�2���6Vu���S�����E;v��+�Y���T��/}���P�Ucś��8�ɣ�������v����>��X��񬢛?\嘬�:6�7�ٟr�����~Ը<צ8�`��X�E�_Ȉ#�Ky��9_�,�`!���RQ`%q%��f��s�Im#Ik�_�k��ǘxـ쎂��R�J����_Ж�f�N#k����Zh�#�m�,a8RTۢԛ������&3���T��̈́���&.$���֖e���x����x���r�xU�#�l٪-��V�� |�v��g(��e����0 ��,����2D�Pv�L�F�őO�z+��p��7�K+X�}�/�� XJ+wZP�)1������д �*�Y�&�q��v�|���yz�4qb�k�N�@��H�F�ef��<�,���ϲ��R�:���K��zH����x!Ki����'�T���&�y9%��;/7 �;`\���k���TAณF�B��L�v1����_�ZT���7��F#Ӌ5>��R�P�}L!������c�>(�[|�Րq����t��a���G�Y��e��?9À�؛�n����Fc��#����ɛ+����A�B�!a�墺�?�OY�&��b�66�i��4�����pV��Oz(e�Ao��\�՗�=��o�+�໘\���5��0��n�"Qwr��&�y��e�/�x-1��6���j°`v��n����ﻐ�8k*=]�v"rmV����ur��4����O�����<[����;+����"�f�x0�jq	���!�H�d��7�
�O��Oo`�x ,S���9؅w���.�G yP�UK�(�x-˹��x�!���]�ʚ8���#����6_�r
J�Y프�g���Ąs��Za�.���A��sZ �-Yڼ�X�ЈKj��3zݯ���EY�[K���[��v��B1�w�-����f���X�9��3�z�}�YW���3�ե{�U[Ic�����Pzh�)�K�ˎ�8��t��U�a���Y���B��*��m�����Y�qAR�:����a�����#���H.5�ZY��4�����ب���l��6�`#�)af��[��$�-�M���x]���ŹX�A��#�ۍ�����������h^b?>ְ�&l��a�?&_ ����b��AC�oR�F�M���'�o��+�}O�;O��llrWI��J݋�#~P�Vn����i*=�n�2���Hɷ�� �_U�Q#��s�s�W��Q�F9C_Oa��m��eط�@�� ������MCCWi0m +�M�T��3��ʔ"�Z!���Ә2�P��|bj��qk�F�oRҍ�	��á�sХ"��V5V*������
���eo}��<矂vOu���
�ݣ�R�ڕ8�9���a�,�T��N��	E;f)D$�}� ���,^�ڹH�yW�w����^�����#2�V^I��Su��� ZD�仒f�e�xh-��+r���!_6;���C���6�DfYl��h�~=���z��1��m��$'ٷ̓G~� �sBr��yc��4�
�K/|��Y���h-��h�5�#;�����|y���^� ꪘ>���=�-��`}�	/E�i0��}!�8�֥�u�)^�Y�snsq?��"�5�s�W6!�Z����G�G�b�M�ٔ)*r,�6v�tsb$ڴm����<��zo����r�J�\+TZ���[�Lj+�EU�0��ښ�CZ������*&:����Vt�F4�
�4lx ��U�t�@��ݿۤȫ�I���*a[�{2�`F�m��E����<@5�Ρ��GH��u��|�A:4���֡�a���&g��һa��qe��D\p���� ����r,�=ޮy��� �����+�z[���~����(��#b�xd� A�\F�^Iɺ@�H[%\+&F$+]'�#��SYu�����������zS��,w��W6�b衟)�����Aky݋A�xDI��ze�Y�獁G��쾣�}x��=N[=�����	�Ċ�ew�\�+?��[�z��.l��1�G9E��j��}�L�ۼT��y�VmK�����S�{zB��vFN��U�i�O��T����	S�q������t�^*�H����R�@HQ�)����HL?Mn)�g�@�<�2��o[x'L�C���4\�A�L3*3�ڽ���	���b�h���J�~�GA�/�jk��Er>��4�B������0��)Nޡ���N�#��o��r��<�R��rZjB�7�^�^�PI�?i���t���w�8jH��Ѐ���Z�����Y���f�$��y�)�������	H٧N=�d����5XL�[[v	���I�������a��� h\�Rn'�m��zi@qV�-`#w\ܫo�O���� ��'L(����w�!h=R�Q��7�1�J{����=G��Zn~Tow0j79�Gl�WH�A$����t��#?��"��^���9�|FrE�L���0_$c�_�+P�D�܍ �m&v;�S�P���W�>� y:k)��̭�é�z�\��L\��0$�.-X�+�Fr��7�QQ�\on�<|���6[��nI\D��J+��9��O�C���(�	�{���%�ҵ��+�LqcM|��T��`$�1��4���ǹ���x�t.�}�<�I�~��
 z�k�Á�x����G~�R�ݐv���wذ�L��B
���a$շ\|?�T��F'��S�X����Ӱ��4���7����;|�84��X�l��"��p�S�u{��&������]��Db:+�}�GI�v ߋ��LW�Z��N} �k�^!�Nr|SA�+T��i�DJ���N*ح�9��"��G-a���&�N����SU��PTmF��E�n<UP��b�`\6P\��ov/>|[\��Y���%6� �$r{Ki)+�ia_e����C�R@:�������F���;�n4�ԉ��4�N}�5�	S��'AOgV=�aU/�9F�����O�37�k�n��l�:��ךa8t���h�g�A��;QJ��<���� b��A.���H�_=�n�S�4������\5nq	r��#'D('�q�Vq�Y�f�x��8��pkR��������2��l�T:L�C,z��Ɔ�.���i�!�&쀳	YG~sl�KÒ����P6��c��^��1�/�Var�E1��� (N�t`����'�����g�F������ �ZT8}�1��p5���#���K����v���3Y		�.[�.:���8D]�h��iXSEV��,���ZY^1h]�7� ����v2(���i�-�HZ!�!��J9��ޘ�k�/�Z<�Kq�~��H�#Y� R&B{ӮNO�:�����gݔ5��A~'�:�>7��t� �9�i��J�p��[��vg��-�FX��D12+���l�%�n�$=-�/�ɿ���0Lp��w8������n����/�P�Xg��2��*d����} *�%�D�]��Lf{��,�X4�����D��z�j�:�����_�����	#Z�6/5_�(#�
lF"�ٴ���fc? �]V�P2��é�mJ��l�ŷ��ڞ��6�.�?���zǽ��|��j~�i��tX�62�×0�=�ϝB�ę����V �q4���=�fV�Zh.3b��`�%�ʦ���.�۵<�i���q-%��/
�* p��u�
�}%�9"'b:[���7:���z����<^2$`h%����O�28�k6�P���R��4[�+|y%�W�yl�o�M�o�X��Jj.��u�xЕ�+����G��7�{� @k�q��/ټ��ي�� �P�j��ۄ���E��>��3��Ḵ���Kx� ����ϗ`�5�:�af�����[��
*�5��Oc�k��o/��� P�#}�h{���������_�i�w�
�
?���F��>�5�\�/��jR0��p�̖7��7�S_�D���L谠��=>v��᭞��]#��S�գ�~͒��h�VD�}�g�Y�����Ɋ��M���Y�[���	���cJ�'�V����a�� J�٨t��Hh��K��CV����T&��[�Xb+�vcv�xM�J�Q$p�~X�-���.T�6��V:F����K�׾C;��&=&?Éd�<��tJ���C�`���h�T3ߵW��U]C�<9�r�L����g7aޚM6`�4��C֔,)n�c�z�Лr�1z��B`�7�zH�ڎ�6E���8����w�l47>X�>�����?l.6��'�z@,����EicM؜�5#:��W~ EM�5djS�N6~��$9Y0i�9B���$�~�����cέ���.�['K=!���p������ƜM�ۍ�_y>��i�<�&��v�U߳�NV������v��7�^�ħ3��j��	]�UX��d�)�����o��A�Ě�\��� g���/�H%M��)��*��ɀz5���3Ӧ�Ë5��ኞ�ONω4X7�Ip�OSZ��|`k�� G.ر�q���c�����-%��p��G��
.Z�QT~���9���fj��*#���f�%�Cg��i�l��,T�`����)D�7N�K��-�~��&��R/����;�9n�I���S��0�׉�iO|`ui��Q���b�n�D&'w�꺺z�
�͵��|���]�YJq����G�e$8��	?��O�F�|�Zi��mr}�ӧ��MM����3_�t�Jۯ�	y�d2L�,�.�A�E)�����q�b��^t���{2ޛ%mqbG�V:��=Iu��]{���c��!��_u���>F��T툠�5�2��VQR\g��:��8N�s'Q1}ӏ�w�YZ�?�>3jVAk'��B)a�#�������ƍ4���l�� k��^�H��DW�NѭIz�����=,Y]�o�8�m3��m2O5W*�1�I,��uv�����:&֎��;F*��]A�kD�>���4[��FDG?�Ā��ܒ��U���-�2M�<�~��z��� %@��}�@TO<��ky0ua�A�@_��	�cD�]��At;�ߦ���U6� �q\O�ON�֟}v�	N�.�O��_�f?U/�ʣ�t����/G��"���> -Cl��(ǆy���-F�β��w�3[�\����]�Y��3Ϛ���.o�3OT�w�y�9��f���Eq3��ۘh��m�^�u��9���;ݪ�clL"E�3h������X{\M3c���]�t�9�n�Bd�t����ovs��P��J`�D��<��ÀY������Ǿ�{\-%�'R^�b닕�`�.A�&��MR�ȅ�m���D�_��.��G�U��An7� �jˠ: ����B^�q�t��s+��s/S�˘e� �s�OE<�'l���7w�J���Qb{�Ok>q��jZ�N=�>��x�'���D�X���nV�?>�ʍ^؎$C�	�)l?�U!w��J�a��-{�"jC?#�G�B}����Y�i���������RbL��v_�]�)G�l�w	�g\�_����(�B�z��Q��G�k=�:�6ˌ���_)Q�]��I�q�2x��w����h�R�I����� '����55��A�0�o���~v��@�;�ɨ~lH�Zu�.�8��]t��ńr���k~ݾ	� �R̫yN�M����q�Vuu-R�;.�p���lKW3j����U���'�?N�N ؆&��jxA���֮�my([�`>/����Ga'S(/iJB^�UN���E�4���p1S��^m���V�B`�iѥj[����=h}9�^����V�r�EKf����^i��WH��s�ж�/6O�k5%��2WIP�}�oAIT�
���4	u-6�C-�?��2�^�.,�0�4�0�8^T�95tR�n��H�������Zf����	�g�˿�5t��P��AL�Ő]�Ɇ,kC���}��2�N-d�,��ԶS�j�[EY�Y��0[Nk!��x��F�v�%P,��;Q��e�@H��Xg?���j���g��4��+�,'��[ӆ�R�T��*i*_�>r��kv��@��T�Aoܽp�4m�N�$��q1�q��=�)�Ieo|r��S@l|��a���܍�⪜k�'~���� ��!�����gI�]�lP^�©[1l���U��&�c���D���_��+_7����4�6��{{��#��.��IJ������
�V����寁=���f7v�[�h���F�;�q -/^���W~������1
4(�,#0a+�?ɮ*�/�|_�%��֋�n1���??�hD��L�{��R<�]ɱf88����Lm0��~ǁ((��q��u��7ҔO[���g׭�n�<�Q��z�-��ܓ�n���
����fm�7z"��~�@U��H<�b�ٺ���^�Y�U^�����ѭ�P����m�O4���d秼��Z��&����m���m��w�z�:��f�	N������<E��rm$��_�����~ù=�^�1_�p�,�*ҿ�tD��j��ܖ���1��L�;�:���>ӥ8�n�a'�_���F)Ǥ���G�>J�/�3����1�:_�<���
`�;F�d_>E�&`K�$6�T�k�ѕh_�"^j�Y�a���|Y�X�t<��3a�8�D@�x0.����|�u�#�t{t�b&	NXy�]
����U>2����H�������bқ����h(I�h� ""bho<�ݿ���\v�̈Dz��M[��5���	�3�"L�eDoa/Tac��[t��qA{��p���cu�1ݱ/�6u��
�Y��e�m�_nQ���^3�����Ń�A��0�d�\��k����R�L&*U�O��A��伅_��b�P��(D�D���X��Gc�OGX��Vc��<�?��W_7�e\�����]�zv�����ީ��]�u��!V?T�͟W^,���!���^������`Ro��k���������'�K����)E
s���G�z±�fR�>��?�����dB�$��	<�Ti�|f�\~p�S6]�Rx��m�@�)pu�JeT�3� J�W�.�ף^��dFB~��+l�Y�NUErl����[����FFB�5f�I�=�8����J����y�q��Ug�9�� u���!j�x�y�SW�����Ft:*3�x�ļ��8Ӄw5p�!���-�;��/5�~���]kI�B~������T\����k��J�2�����7^�sl����`��aa�����خ9K�*��b�V�ٯ��jf�|;��{qn+��,)9��j����N���@���S��GE#�6���y�i��g��#�1b�C��:�Y _�C*��b�6�Iy��m��65O������z���c�m�P�N���&R�����#_
���s0��<�������z�s���(&�˴f�C�ܰ"��[��¦d�|�q[z0qw��WK6�gE��3LeB1�$l�(�H�\�������>��m�׵Dgljt~d����g]ۚ�~aIe[ &�D�>Χɼk����*���^җO�T��"���`��ڒC�#x@#s~��"��_��q�}�߽���+2��|��L����������W���L��?����P��/�7�X�{��\_��`ȑl�ˆTIr�+O8n.7}�J�f��W7������j\F��M������|��@�3�jH}H�x{�#)��T�uw����0Y����X���kX��Ec싾j]��?���������h��@�W���0c��^���Zb3��,�qZ�����!L8E��v��&ؿ�r��1-��y6�]���ȭ��W9,����o�Մ�ф
1Rw�����w�DD9pܜ�VT�+@���؁
�ه��Fe�M�w:�g�����9�/��F�C	���+��z���p(>�?���U0�N�s�)(��Fe�w����[_K�U���?g��z�V7��>�̘�	��_�3��+�D�J<��O���om�H������vc�!s�����ږO��h#��kxywM�z��ĲXX���,���@C�5w��brnW�g��Iρf�*�Jl�¥�P:�sdkv8yo�~Ei�U ���	[fը}��U)�oR�#�� �gD�υ,2�X���:+���[).���Ӂ����ȧz��\u�Q�� �b��τT��a.��i�y�]��_R'�����g��^&(������x������dh�;�&�;���\KN���{۵�Ǧό��v��s�h@/����ǣ�N�ѥ߿>�!Eb3a�:"���͜����y=�z�O�aj�� Ԑ�z��Ӻˆ����T�x\	R���?��2D��_�?����b�Ԑ|��^��G�		�717���2α��k������®*ʈɄ��m��vQ攳(�hM�&*2o�]�2yʂtq�"���>��66}�+��"�EQёS���,La�;-���-1Z��s�i���o-�^>t��*�U.��A0�M�΄|)��{����8||�ݑS����G�l��x�8&yU�>#(��ԺQ{��`<�Қ������Q*��f�S�2�E��c�U�C�A�t?)������XG�c��=�J1
S�k��P��O��0B|j�[�B��P�ѳ?�6DBT������pnu�U�V��`|��������s��S9[4�L�_A>�5D�R�:�;�,6��B��Mn�)�����Y���}�ͩ��Y���|�r�1N8\B�L�?-Z�������b���F�RJ���C2��b{����	�S]�z�c�i$���;�hT.�
�	n�ew���j��n���Y��"Lf��� �?�P5/[��␲�"��Z	Ĥ���n��rm}9���؊	P�Ш�>{"����K�ݬh�;�(�1)S�&N{�k���TJED��ɮK-2��@��3�J�0��V�xK�����J$�$VzQ��[^[q
M�1~�,�����y8����d�1>�5	\�;0��4.�F_b;Qd�9�b>�񰤳\�S[�A�hE����˩�
ד��I/���d����F��į��q��m��|^P�'c�Pm_\)l���0=X�?��X�F��U� ����&��Vʖ!rc��P�^#�@tי��:�~���ݾ��Sz����w&����Ҧ����I3��FnC���
���Y? &<l��Bڳi�0�8Һ�<$
!{�!C]���$�a��$��A[aP�9d���ӌ�8�JN�f�H����A	�`&\k�4����{���*Pl�*�ckQ���B#�'�Q{U�,�$Ig��4��~;��������\IL��y:_\773]æG��ҭ�����v�E߼���r�E�ιg���+��r�7F�y@w(���zA���kҔ�o�WO�ɉM���N`f�m�]�s��׶�J���
�i��H�("�;ܫW�Hl�Z�	�'D�M� ���q5`�S��k�O�n��� �������'g3��H�+Xd6�Xz����x�%�?�MR�@H;��J`�:!�Jo(m��K{]����J�-4-��e�g���2��fE�D\�<s�k�'�oѫ��g�=E��B�*��K{i@�����RKs=����|ً���yz+�Oc-N^�P x4*»����}I�aײ��l�KUl�Mv�պs�EL� ��D.Ă�<ThR���D�z��|E�MN]�"��h�	5�Ap�|���`G������G{�m�o�ƾX���+����A
�^.b_�������7�/R?v�ݸ�o�2���1�v�`(!�p�gY"�U|���k�TPT���@W�	ƻ��m>gL]av}�ml9+Z�0��W�\~��4ů�ߕNb���~���mW�*�j�YF}��W���^���]��Kkzj~w$=?�)�<_f�
�c{�v#�H�H�9���grZx��t;�f��}���H��Z�Z�n0��.��f����<���&��f*�V�_����/6y�* `�~8fK�j����?]�ĳ�1�z�{��{h����<��=XUȗ����%�_� ��� �G�s
�1�\����:y3��������B*���G,�7q^E��	 S�j��c����������>F��#ר
e�F����sC��Z��ѳ��7h���ʃv�O�"Xs=�sT��F+{#3T����@�?O����B���u>7����±K��Bt_��N����O%و�t�JSNT�E��h�1����Qhq�B��A��8ot����&G~;�g(k�k��Z�wt��oL��)ј��"B'�9�gY�w{�����Ye��UV�����W�O�W�bL�ͫ8�����~� ���'
�Cy�`�{��Ʌ����l�;ޗ)�+�����B��q�&��W�k��臌���W!Þe�Z�.w�K�Z���3��P����B�� okQ}��W�U�F+���ʨo�FN�q>��?�5��c��X��i���6�/��.��Xe��#,�O?z�o�C�o�����uVqk��\�V�;�Ade4�#\�&;z����� xX�E��\̭�ҲY{*������ -\=�3���Ɂ���z��,t���}c��1\�qQ;�s���c�K�(��Z-������SIQ�օ����#����3�b�F�j^�z����\��7�6�=3fZ~����6��|`g�h#����������'q��/���n��^�r{�>*W��>h�ښR�D�o�t6$@���6!�a�l?{�'h��,p��{d���SN�4�[)h&P����q�a�)LJ#��q���b�w��&�#���ګ�7�	���8��
���ܒu�V�s4�!m�G�\Xm�{(;���=��{�w�V�'
KZOBt{��0����Aq�D]��՝��4%X����� ���qv�/���c�1�/#t03Vum0�^o���/����gYi|�M�����
�$���k�kGU� ��OιI�_R�iU������������qg,'sr4]|�����ޫjA(���B���.,�� �>;@j�:�+��qjw�V�����¤���-�5�05>���9�\��`f��k��b L�}�gn4�ًm�D�pV^��5�Tc�}pfD�,�%��D��4���d-q��ќ$�LL#黨tz'SU��	��V���:v�#e딕��H��w�?:3ڰ��C�@߷�B�..��v���D�+��}�c��e˓�5��N��^~����O�et�5�.�8o�PtjC<l��>'B����~�0Ō95��`ɰV3!�ڽ�?�M�RR��j�qz��Tb#A�)���闀~��
 ��2f�	�?�w���@LaĞ�!�S��Ѿ��6w\>6�{��f#0=k��!���rqSLy�"��n&��d0 i]ٵ�揄,����Y�п9�/�g��'կR:܇3~<"]��Jf��L.>�t˒�˒h�;�~:��
��E!�!�<ze4l��W�?�$}��k=C��kd���I:���ZEpy��p��^���G~h(�I�2xH
����Qj��f�K�n��v)S��:� x~mr���bS}r� Hb%m&h���Hm]���օeJ/�,h��.�kZ���d������4�96����2�A��ά��(�M��V�ⅱP�l0Lhac���4$��C�q�u��-�����@�;/tXd_�9N�o*���3����;Z��\)X�x���>�,����D��0	����Π�x��}�E�.�l�度5Ү��A#�����˃C��=@�`�nM�5��ku�Mk��9��W]"#�����H��r�;�xΛ��Ƒ4��]�4�}|>���~��#�a��떶��]/���TFȗ��0�2�?�wg�$�Խ�f���� �" �;
����o�9H�ࡑ�qwX�6�1Q�`��uM]�����|��6E9�we3�:��$��,g���<I��ԅ�]T�}��g�8i���߾>���op�e��t,#��E���8ITZ��UD�f&��]zdޔ��t^-��oZ�z��p��X6��z��P���K.6�����x�e�c��m���} ���U7�w~ܝ;�ꞧ���e����3�-y��4~�6D��U�a?��%�$�a�3�8d�a�%8�ӫ9�7������zk�I]��6�cL�c�P�P�󟕂�����sfP,w��"�4�U�J���|��'�!��F�P���g���R�F��G�m)� �ʳ��}�}3>��i? o�p������&�Gwଭ���Rm'�.�����f�2�ux�Q�0��x������~ӋG��4hx`���`� 7�'�q����|����|{F�����%��߹2�Pz�;?+d�e���� ����_ô#'5檗�6�_ǖ	�Zr�F��Ơ�gLq2i.�i�C�HJ�&��ǿ��e�}>�lv��X!����~���^����.�/��u�M�(ş�F�FDH�����v�%���|�y�N��v��g[0=v�I1�-9������Z��nt�=���܃��W7�CH��M�)Fgx��8*U�_�Qr'���_(RĽ�ԋ������,��YOq��h���c7p����uCybO��ӬH�lC޸���L��K�1G������j>!4�	��n���!�z��AuL��xt	6�(a�B
���f���*����\��}Ow�+"5?�2�}~{e�k>J5���~J���_ZO;r�X�K#�'2����߼2	ظ��I_�U�9:�����������ߟ'��˭���`|x%(��Jѯ�R�����q��z<u�>��M���~���{��"/KsA�����u�A�A��:#
*�˾f��!���7�1#����+"�K/V�4��=����CX�TR� �8���b��Mwy�|{����o/)���I�xx�<�٨�g��>koӶ�K���pɆ�Ek�@�����=8��V�5�2�~&�>wc�%Y�����V[�#}��z�<�ቌ%%��"���$�����F��]��M=(Ȓ3j�Yp���
�!(�6ւ>㋝ϯ��GIS$���ED7Eätr�{N^H�"�����Z�?X��6��Uy"D\q�g�I��K�����}����9�T���쐑���9������9�V�`���*!�l�Kn�3��4C��;4��$~i�����[/���(��&�EA.������FiZ㚣'���e52a'i?��%@�b��l"�s����q���6��Rs�DmzA�ڃ�q"ky�&��B��Ƶ9m�Im2x�y�z�js:���dS�:;Q�'�N΢2������C�����A���ݺ3	���#l��)�-W��zw�>% �~�՗�I+��xT�1���x>0���sRK��J%#	�"l�����*Ɏ�GX�①�g>}�N;���k�~�9�xH'E}��c~?�{|�/����~���
�9���Jƭ��#6��*��׊�
�o�/<�S"]υ���ܳ����g����z_VZ��l�_/;"�K*�G
+��d���a���ӫ+�~d��.a���������h%K�ֹ`�C�O����6m����ض�:`Tfaφ�j���*RIC�K�O��A��p���E/�+��f�=`j8��`X���sA2�Os������iM[Q����<��'�y�Xۦ�Kk.@����E��UF*��4�b��xkl�fN,���Ҵ'>��F�^��f�[:'7A�ھn���q.���6#����8�XI�{+���v�.���]5�ڊW��Rv��]��eD���u>�dË������S��&£fsc;J���k�w?� ��[�}r`����+����w+'do�c!	p|j�~w=�H�u�I7������:�E"Ƃ�Q��wJz���(}�ֶ��B�Z����7���e�a��#�χYy�U�m��i����n��L4�����SPGx3�u����˖�c��d���VD�9+��T|�l�O���'�G���yٝD��J�xq�<��5\}�`��{ף��5ER�#A���`�U���nTc�%�c���}�v�rLW�����´{[y`0B�w~�u�e���yo�`�IZ�םG�	�x�3~0�]σ ��81�%ĄU����ޤ��z"?ڌ�Gn�ɋTP�so�3�|�j9�f�i_��ns������<��HB� ��zb�M���LЭcn����T|C���|�1�J5ۙ������!�z����oѢwY��>z��H˧�el��@W6�Pm�\��X�vX�O���ï!��ue�.�.���z|�\������yث��cuD�'����n]��f�D�)����%$|�c�
C@:,�-i�#�d�
ӥ^&��T��p��:�M_�����W>w�`SNѠZ|~���X�٭!ռA~��F	J�' V����؉o�
' A��*�2=+,��$v�Li�O����.u֞�̧�A��7<��-hֳB���T�&�
�:��p,/	V�s��c��3CCn����y�mh&y����ꭟ;��$n-?m���n?fԱ4������T5m.뚞ꅾ�?A���_���1+zE��/�	(�]������:����z�<�r-;V�/�.�Xh�:��n�xl��b;�`s���?��(�����b��
~�w���9�W�G�3|��a�;�H0�	}���uj!�K��?V�@�N:�)�E�O��q9��F4Wy2R�6�1��d��\9,�������
��m>�,d\�& ���hغ:ѿܮ/0��X-�^+��S���I���EV��pC�w�l���J{ʣ��vv:{v@(�-��'�)@�(Ki ��z���ӎ���)��.?<f��Ŋ#J�&\�Q��uiO��e���+��3���c	,vo}���<;�[��!��T��Q-�ڂ�ځ��ȫ�Q^������V�9�>
o�#�*��8���~%%�ѝE{��7"���WS�@�����o����϶mײ�l�l{ٶ���2��e�jiq�>a��S{~�����s��q������;�r��v�\��=o����TF����p>�!�-�6�1�d����n��j�N�hW:��A�V`�:k�)k������۞�[��Xً�ݷ�Y�xV��-��#%��P���{-�������L�p��2Ϟ�钚 `y��܆ԑq�4|�iCA<�6VEv�E���d�J������d|R�5i	��$�Tj�z<{�$��Z#cԺs�('��%m�V^\�������=����a	saJqe�?�s���������G$��6my�3ԛ��OnT��k�at��'ǽ�V��WIu+�+��-����$}8|��i�o/_��j}���ٚ��gP2�q8��r_N@�(,������>,"�SR���5��sk֪2.��%�w�gƣ_�<���lr��pD�`'J��+�;�^	�Û%�zk��&����g��F�#O�L��o�FC�[ Q�ocgQM�"e9�>�[!�*��i�i=z~� �=$���4����Fe����<O�,ÈD��𵺗&P�w1�����w~��$g+T����M�R��� ^hD�ċ?�X6_���ހL�l����	��/Ω��0_U6H������/"?;��0�n��A,��ç�ߧKQ�F9[M�������DңĄuW����+?�Q%54���|���T-ƒ�:�&Pr��0{�y(u����9�)�%��y����JEDn��~ٯB6���m/�Р���'nP��`����_��WlQ�k,�0���@����⧳��~U�0v~��*8�-|Cx��O��Y��걖�
�Ld
�����Z��\��D��ps5��Y�����_�eK*�UN���������#~l�ȣ�U��|���2�>!d_~n�0����i��4���(�a���qWŉ��q�wN�Ȉ�9)���7�Ǚ��׾{Xl�Ai�(\ߐ���X"�����]-q�9�L=*�ΰx�7��qSB3@�0v�[��m���"?�d�h��!c�3$ q�vh�N;a�x|�.��%�Y7���n�&�*|((#�\r�kzi�rk�˴Ye����~��={��J�Ʀ��a�x����N�W�@l�T8�z��6�'�ٚ҅=����+�*�c�w�wM�$g$'��}��߆Y����/���]h/<�e�gU_x4��1�\��4Y)�7�j���Q`H�Pƺ�}�˗�-g�Η/�[~�����?���\Mo9.�R|GW�ew���5���dX�`O�O��G�o�&]�ή��p����Y�oh}5-��z��h�z=��F�8N~�ԋ����{6�@	f�~�{
3�VNjҙD���UG��LJ�]�1�7A���G_(���`���<w�ا`.��������=}��b��_�@r�������j�f��]Hj��8y{��3D�H��]樜�'Z�C7$s����ߵ|^�k*��>�G��5�P���9��5�U#QZC�R�\
��b���B&Cj��yy����uI�OOv˃x���պ�\m���&�/��m�:r�ܴۤ5��o�W�rW{�UP�/�Պ)�G�n�b[#��6a߳��E'��:D~�7���)����}R!�S%���Sf��S�|Ժ�6��$g�EHK���hms�<Q�v���-Ħ�"
�r��ׄ1���wq��t����,$2v��8�8���w�
ߵ���qM ��ׄ:��AA�PF�X���m�`���������w�j���b�/q�A�RĐ�G��}��mm^^g��v���5TS�(���Vw��#3�_�	�Z�7��0�CU��r���;�$��xu,����3�͐��K���_���XZ`�#N����kv��y���m��j�&5ko�(��ߐ�,�����[?Q��7-�b Pkk���o)ba��?"��l���o�Ll�lW�9K���K�MAd�·"����[L]�M�.d��(�g�v�5��rw��t6���ӱ<�yC.Zc{�w���@�6M��Xe�b+̾Cjx�p��T���7�w���ϕ�����a�J�*���3�T~�ɂY
�u�^珺Yf\xI�R�T�w'�ۛ�'�-��]��<�ɩ�~Q�U�}�ːOf�ԆzF�V�ЖS�^@K�ߦ퓖�(�Tڗ�F��t�]��wV)�'���� m��c4�,}~wF!�[�:4��++{�ZL'6(F�B���>���H�<�Y���aE����*Ċ�oz�����t����EC�����K�p��8�AW�đڲ}m.��>��C7M��
/̷��A�y����*�౥��y(�`r	�?*����-Ō����;�����|-@�N����Dt���-��!�v�hB�~s�O�mJ%���Ԟ���'8�<��Kjg�Xb�k��X��} CĐz�i&���eó&��I{.�ѷc��1�^�̂���|��e�8IU�t9D����P%#8�()��Z�z�Q��f��OP�~jI��r#�xo��.6�j����b��S�ܢ�f��FM���3�tTIU'<��	�lĳ����A�2����8x�C�u8hR��Љg�����:
��x��"^p� �`p}w�=�l>��Z����f����s����'u��9</C��a���8<}vւ��Oe-���AJ�]7��j��_�~��b�M�����b2�����?��ky���cխv�$A�
���f�b�V��} �`�M}(";%�ei��{��?Xbſ����%�c��Q�����Ll����D��lL�gt��f�����R�n1��}J�Z����[}���u��Q�����42�+�J�K&��B䏑z�.���5EwG�F(� u�&�~�kH.r��	���b��?����_X�8��������d��A��
�X�q�׷�A�?4��꠭݋���"i�V``��p��T�����Ĳ���~�9@� ��(���4wP��#4D��V�& I���u!ڷDn�N���9U��[��no�IzHc�X�"p�S�V�X*��Mݤ���FH�AY.���e�bY��kU-�KD�l��#��� ������w-y�OE$��ƳN�پ��C���+o9�����)#y�ͯ]��n}-�ƒah.�n�i��)��r�F�P9���Ab�*� ��r-����,�6o��?��5+XC���4s�{\�bë�=�ӆZ	2����Qf"I����:�Q��L�V�Jo-�3�4�E��&����5#�G��%IF�����vM����[��\��B��a�$���_߻t�ιE��)�:~���#4oO��J<����6ل���ng����Xm�oI�iK�!2�B��W_��:��Ü�g��ȏtx���&���44(�j@��7��0EZ������e�l�gҚ�R2 ��Tv�]TO�v'�n#��A4v�W���z_�"��R4H���@F-9��
�%�a_�)fN�|���U�_L�����a�Z�� ��=�����%�E陈S�^]G<�4�x�O�QcwP$�>\Ap:�8��g�1��.�uF��܆F�%u�Ԗ �
e�����V	����] ����*H^��of����0p��[�臠VGT0f'�b�S�X�T���
�~�X��m�/��6옸��v���hPo��@�I���:]��6U���O�S��SSI���o:�cI��ӻ�=��;�^iӸ�j)�b�/�d@��:����p U#>�N顳r��\/ގ,��yY�\�����K�/ t�?:�������&M��(Dt�[ǫ�`��MjZ���y�D� Wo����V��(��)���[���`������:����cj��y�7�}3*�,��I�v��Og�2��e=�^]|�b����;�(�Y�\����b2�(-P���q	,�V���]%�0��?Ѭ%Wբube�!G�"P��N���ǃ_~:�MLr�'�8��a�{��/g��N��m��ɩrv�a����4����#u���p¶%��S<�./�4]-���G�q� �$���8�)�4�-�'�|�)&Sj�g��!dR�中��H��j̩	�זC� M)8�xE�
����G(���P����^����$aɛ[�U���x��B~��ʷC7[T���]�#�����'#�=<�G��b~--$�8������!uc�R�4���kۜ;fQJV��i���/��,X��c{;g�W��aa�i���511���(��3#���燁L�\�gA^���)�{�1.���<�ň~�|Ue!���w�P�P��G��6�&I�`�(�Ul�TQ��g��FW��ayt*�Z`.��o��y����X[�Us����3���5��a@�=��/;#`�G��Y��
�D>nd��Ϥ�b��N�(�?w1�Gz��� !6�Ь��Ɛ0˭4�.I�>zU�-��M*��	�-Ħ�pex��ϝZ�]
-D�7]x��ep�7#�G�t� 8:�f2sB8�w�i177����nǄ{p6GL�W[[t��Eo�G %��aN%R$ =?8�����7PXݴ�=
�ZZ��������J\7N��ϾB;A�8���a�Hڝ��<0�7j}|�=��E����A�,ҍ�ȹ&H]����*Yc�MJ�Gى��e+�����_��ٞY�b�w�htx�����Z)J���09�`���c�m��n������`�M5��VL��(ٞ��`�Ċ_[��Yt��C��o��R8�X&9M����ڬ8E[���"��wN�����t�n����k�����߆� T���Vy*���-C~�X2gJ.� ��V\#�[��/u�ձ��!�C&U�	�{ �$�7�5h���آ��8�2%�T�%�eU-E����6�P�ܦG87�qߚ��&�pW��	�
�-��@OX$�<�"��菫����$SbXF���_�1^,$���1��;���`8{��c���'�/5��< c�E%��~;�~R�����ឞ��E7���i����VMJ|]X�hG��N�Ű��i�V�������ʚj`E��h���|L��WV��/��Ш�12���ˎg3d�����+LzX�_񘰛��Kd�Wl˯�D9����W���=0������tC[	�͟��2�A�t�Z� ��(	Ÿ����DV~Y�1���� �����ݎ�`v œBΊ��F���.�
\%���@�~S�b� �)��_��x��r-=��d���9���;��6�}�0�� �˼"���+�lɞ�q��]T���R+��ԍ�$����"UG���X�;���nW�3����׏/80���kJ���B)#]�7Sm9���<?�4��̈́Wń�����H�8:D�~�1{�^_�&y?XX�����o��x��:���#�v���è"�lcF(��L�yk��#��W+� ��a�J{Fy�@�߈w��� c��W�����Z�)��&I��[l:�~$Y��f���h�36xk[��r5+5�h�)`t�n��2n���X bG�t�.	�0Da�o���]c6�1D'�*FS��"�m0Q�r���!Zk���`�+Κ�:�N�"�4��;I�2��NV��@�o��������h��G
ݏ�Y|B\7�w��J'��Q����n�~��}���A��D���H�\��5���r������{��]&̿.��AB���onNߘQ�}��6�"T�\�-n%����lֈ�+a����p�,�9���U`�v��b��rJ�GiA}��D\��.n��e�}UM�	U���#�D����J�DB�_��P��y�}��	j��{^��AT�3:q���������[�������͊ػRTIMh��s_34�b�7�e���y���O�))A�(�ќd��?��5�S�#�*pC>��:�����o�s	S�C�'�2K�uCjp�V>X���.�"���{/N�����+!y�}-�[�>1�������~��ʠx7M~����D����̄�̈����>�ݿ���g��:�l��X?@ؚm(I|�*A?�ŧ��ǒj���m0���6N�������.�Edt^źTĕu���B���4Jnk;}r���4J����$]�&14X�_^.L��0�_ڗ�Y�H�����}2�j#:9C���+vK5���z����+
N0������S7J���[J,������)��7�/�}��IBB��';�=ɐq����J��v��Q�EM��˞ۊ��, �������}�u2;�\�߃�`b�k����#�]��(W��6/�L��\��/˦1�އ�'wǲ%������<��#�_��x d5U�g��x^_�,@/�רa�o��5	�M��DR�x��H�o㖋��D���g<<���	�����9�[U9E�:�ߓ9k��^g��\ݼn�J� �`o��1aMR"��!��I��7�R��v��a�h���DP�� c=�:KX�cJO��ǌ�x��^V u�5�{VwS�,����9�T�ʛT�ܮ����4���"Ҩ�I1��O��������6��`��@�i���q+��-U�}���P����7�����<5U��H�H:��Ud��-�s�M&�{	�x)�Oh��V��kxH�H1X�L��to�O\v��Υh�Z*aa��l�ķ?��m�\�XK��z(v.a�o��̾��3�MX�(��糖>>�Q�g�w�w�����>��!6�0g�����},�.5���>ƐD׵�"�g��N�qz;����V�4÷ t�Y�no��3�S��S��pE�3�~���Uf %W��wؚ�Ϸ�s��iwk:聚�$�[<���3� @sʶ���N�I�M�BY��|R��m�:��a��ɀg���hĩ9�{@�~�K!��� x��b]o��]W�<�o����2��,���-�T8C<�ZP�X&J�h׭�z�x���]����c�໘$l�X��y�.Vi}�J�*���ߝy�៊�kj�/�R�( �4��5��l9o���_��IE���-d��O��R� p����q�������^�a��cm��M�uԎ�HV���2�=h����8>�V�U�L�h�6�6��'�[d���,3�E6W?�[UF�d��`�)k���cX�y� V���VI�M��'��	oX��K6���}������H�X��X,��X.y������Җ��I���N�A�/��v����T��O�w���̡ �2*0rm%0��S9�&�čs��!����~�/�֮��~��%z�[�G4�|�I��)�Ϸ`x����:'��-$=a)�~���H����}�3�:�K]�o+)�$�w��B��dha)Y-�ϯ�ߏ��1�	n b��o���/f�7��C�O5�8�Ѹ�����M�v�(H�q3�?x�	�[Ͼ��]���^y�:-[��� ��4N(�}���oX��׻D#"6�d�H�(ۉ����)���:{����u�R�Sw�S�wk)�֞�
�&Y��n��Vm߁
tv�+�T��2�iƮ�x��VJ�i��K4b}� �χ���_]���b�l&�&�p�r�4�Wƃ�,�g��4�"LF�V=�,s�s��Yo��&�LEץ�tƓu�6C��at-32���6����s5�\��lS�PX4���/G���|l�K���JnC��]����~���N@�q�OV�{f!Ú����[�r�'z�h���n8��[/M�s��V��ޤ0K>ƞj��rO���RL;�+��t���T�_S�d4E.�T ���Os�W3􎣒D<���F��m���儋Snԧ�B�G�Ȑ��h�8�	�%��0iR�Zx�9gkib�$/o�5���d��;�ݟJ=�e�=u�OH�	�L�e�KҺq�Jg�"����P4c��k�W���ñ��
���[4��������8����,�x�L B���$!1��������	S�7ӳ����{`29ݓS�yiFM��$o�����"j`KD�yF���*̉��ۗ��z��������h���0��^���t��|/��QtB�1��A"�V��9jS�ۗ�K�FZS��J�6u��dO>ʶ'i��TQ�g�"5Їk׉}�n'LJ93�(��B5:�c�ݎF}@K@!�|�Hm'�j��'�*7�����7�(\a��z�`ɨZz�'p�}��3{E������L\H?������h����k�]�k�aHS�c1<�Ae�6�}����j�D����ޚ}�T��?Ѹ�m_�L|/ɯ�% '���f�v%!^�B�`i"/6v�6o����'���%f
��N5���;'/lL):ק��Ƭ��՝���]k���f�7El@�z<疨,"X�}���/���s̔e�:k���5KH�|ϖ�B����k�+�*=�j�*X��ќQ[]�|����5%��lP�V���;�˓(iPa���$QZc�bY {D�{��;D{�O�϶&��V�P9�AR
�J����B�R}���P;�+s�9#9��~���c0�ʮ�x��Am &�7ټ8
�".VӲSi��
��U�6ƅ�z_�Y��ۗ�h��F�Ӳ�b�C_�^,: }�7g}���oR �E9���3���]S0 ��8�]�f��+1�Q������Bv	W[m���[�^&����B�<���l�V9�Ѡ��ٯ,!���\�g"�m�~���j3��J�X�5�Èǫ$x��"R�g=����w��AbY����N���y��B�nT�=y����@��4ƀWF�?9�s8ut�ѿ���χN��s��Ώ����Yx���dا��sn����}�Х�ↈ?��}�1:M�������c��4�.�ɍ��'rF�nt��t�c8�
������/��v?`�h8�����_�3G{���0�^����a���n�� ;�)�^60�%]��'�[*��t��������`������cz� ��Z��%j�<��w]�o�=��J�A_Xӕ�,s�~C�sN!ת�z��?}.;sd��k����Ϫ��e'���}�l�\3���~� ۊ��Mc%_����'M���/���c�\����d�ο�����TDG���V������g=�%����(���a��R���g�Y���(�?����(�U�7��5��7ɿ#p��G� �՗E�m�я�N��=����m]��d��g��V~��C>�d��@=�p�R�dg;ȝ���3���s
�PaY�����~y)�?�UkO�x���d;�$����ߡ�C�{K5U���G��}5��˧HP?�5<�v���5W^Ŝ��@n��#˽�g�֖2t7=x�7�W���� e��Y�t��:i�٦%k4��~����cŗ��U��! �l��Q�� UA�C�^�	� rJ�ڱ�z���(�����_�8������ؚ�Ft�[�v��ܜљ�����Sw	�ѡ��(F�׌�|����X����}�/Oq��P�O;�܂ωs��v�7�G����7��|4;�������j����H�j��1+�r��ᨻ�rG3��D�Pk.�A$n��]�� ���nѠ8.X[ +�֪2�O���z��QG�H&1�O��]��No�[�Z2�v�B�F��OA�|L����
/�b��Uթ��ko�����*[�ECO%�j�%�yԨ2y&}xN.犓�������vgM�6��+�L�P�����}za�{>ag����0n��4,�r��pW�,�:r����5;ل���@�c.C�o��/iL:F�Q��"(�5nR�N)����Dtucے��/3�T��?�a��b#�e�Ӆ�W�n����'�H�R���_}�+�'4`q���H��ĈpnX�r��g�1�h��]0���=�Q��/��K��Eq�+i�~�ψ��&8�G��-F��=�WsZ��yV�ƨ���Yx���ԗP%|�4�V�����B&� |N�7�CQ*����^'�Q��+�ݩ���Pa�h�30�G��e��_����gUV䥿���V�<�*#Y_go젧��'����ߣ�����u���io�d�.D8���a��L9��q.��xu�,����Z}5$���nڕ7a��&ӽ�D�՜�������Z��Ob]S�E�}U����ͯ�����H�u� V�5��;������D=�W�cq����}>���/�;�Uګ�����a-�2	�����|�~�l5S�����A�^�O�fTߋõ�<λ�:T����-K�2�	}�>�,�0�����kϙ��=�y��aj�d`Z9���K7���o�L^ן�zĎ�]���*������O�(�(\���w����Z`,���gFk���T��%5�'}ݹ������r��lVC���`��
<���aqS��
�˵�}UE̦�sM �	4���r��AY���Z��c���Hy��ef�e_N�p���/;G�ZC0��9�A���q>+����}(A�ĚB�A4�T_3T����C,*$h=�s�'�
y!+�������d��Ŀ�{@JS�|���i�۞����i�ɲ�Q�BB�\�x&@A��w@�׮��Y6���=����O��VF@����$��4�~Bu�{�|�A�'���kTSJ��zY�*[��aa�����÷��&��-X�����*��������� ��5X�(�-�6l����M��q�<���Xҵ����w�s�4�	��[�������~�{��k��[Wv�Jی1���Z�F>(id�SV��NG��[���7�L{Hb�;�n��1�1u\��ɩ�T���NZym)�s��]|Q�k���9E<>�-��0�+!������
�3��BV~H7��Vt <rYV1v��~K)Mb�BB�� �F��F������I-��Cz�Xܮ�1b��E�A�ޖ�?�N��N��� 4�O����>����(�	Ɩ��]�^��^����nb�^N]!{xP��5\�h�N�4{|͚W�CD�W8��Ϧ�ϱ/��Nb4�՟��e\ʯ����Za��Ó�z�X�l-�i�k���_����6��������l�.g-�����\� � �-K;�r����im[������"��5�(�Ԧq]�9?���i,;��T2;��N]���Zq��N�#͘�k'����v~+l�B��|i<!5��k�7���,9Fp�J��?��AfnX&��
�f�j'͙�p�y��Q�i� _;>��Ѷ��OǞ�j��5 �QԢri��Ю�k<���	��ާ�yl�i���l[�S�� 1>o�(�hk��ا�tA�l�!���4�TF�\���G��t�Wjja�.�_����+� �HW3�e�>���Y�VZ+��<�S��E����WQR9t�Y>�Q��'�*���fs��!b^�A®R��k;>� ���ͳ�"����&��2�S���<V}5�]�	�Yu����m�J�����/��4�ԺC�zĐE硋~�Hyb#�ڋ�Y�G���S���E w{VODB��6�SK(�I�.�j��g��A� ұY��M��Ӎ.��tu�b��ыɌv�ё��l�%�^�t��>���ފ����'i�~�S,R�[��i����/z�S�3;&DU��a�v�rͶ�Z6�bI-����B$��/�JD����^�.5^^�.G��~U�{K��;���X��A,ഓ��l�_�N�]�U^ �o�l�;�aI�t|��{���KJ$�`��-H�����Nbu8k�$��6�4��������M���4��B�~cFQ��8L)���SYɣ�<�f_�����_�#�նX����i�H��w�ɖ��*N&�R�콞�^�Y�؅K�LH�K�QXb�Ψ�93`�j�2���衵Ei6����0�^8s��jG�I�0)���yц@��O�ES�i� �	�r�1�g��>����&n�X9|�rI4N���x�龜�MCu���r�����I�o)G��{A](�W(�c���p~ag�����u q�h`�����ɭ7��΃�IW"��ԉ'���J{�Q��
��m��ʇMVTA�x*�i����3��u7DN�C�T�P���%יF]tג/�c���n�_(�vt��_�AZh�S�����E�d�;9��������ͯڞ\a���c�����>����͐-�J��@��<C1N"���K�.�\s�1l�q�7��I���<,�c	ոo�j[}}�!6�)g+����?[Q<鸷�3���=��0�syH��I"���J,Kў_�b'�PQBy���؞&-}c~�)�usC�rF%L�@H�&α��4�|�X2�jDm6�V
����S��T*;��I���p��t�y^�gLH?���1�	�T|�0)��I%F��U`�S0�>�(���p��nmUq�
U����;́B2Y�1���7A3<]EE��Jw����'í�"�$N^6$)I����{�*��f���#ƀ(�4�����Y*�޹����ҭ��&��	��`'KO�����j*���
rəO��z	��x�̒�I�a7����Pk�g�#��<+��W�H�.�.���h��5��k+�����>R���ϙ��euIg��m71ݟ��\��y�_�Em���j��"Z�D�ze?pY�h2��2NN�
OT���ō�OE��ӛ��;�(	UA�0!�n�ۦ���t����vf�Z�4�fR�4���C%�X�D���u�G����T{��D�N��_>_�0�Op�ObJ K ����,��*hU{?~�K�u �5������CXeG���m�5���ͭkuJ[*F�	��f��$b�T��q��$�_�S�A�8b��^TIٶ̰
�Hcl}p;��'�/efT
�3�j��~gC3��de!����k�XO��S ����@���~��L���!Hp����(���?-!�Ta�?B����=ݯ��Us�'����Gy���,B�}�,��z*L��K �Lsڦ�b=�m|.�B�֜���Q
W���?���W�Б��3'Ԑͫ�:N���9�)�+m��a��6�������FH�2��K�����C�:c@Awk_����A1�~?���8�K{��Q0������Y-=�^��l�}�:H���fm@�+FY��[=`����Hpq�U .[�Wz��wwaL����q;D�����$3}��3�,�bwu!�S��V{界�r����Wv1��_�GQКy��T�i��Z���L���c9n�؝��6�x��Ȗ`�EA���"�D4n6�Ҹ�R��qC��q���Q�����I�\2�i$j��n�o:ֿ�3����
|�8��iT���	C��ƳV7򟭧�;-�x�L�y�����.�x�~���7������=�fGC>��c�I���b�����$|bΣ^��(.�쓍��<�6��
@@���,���ē��bM�ï\������;1�G1����}c�vKtҡZV)�̷�Xy@eS.Z������}��\&�(�ZR���ܢ�p��C~^T4�y���ڦca���HY��a�[&��N�0��}�����	J�W�D�gm�5TK�_� ɲ���b��i[I�&mW$:���J��{��~�@�iB�T4)�rC��㉧b��Sn�F�����Cȏ��2��9Y��%���Q�"���f�7[j<h�@��Ś!��
�`�.��͉4T �����b�9�n��t�� ag3�_~�9�=��n���u2��Ld�e�)�	;<A���)���FN��L����"T^��V��뱠��+��N��ֻk�8F�N�d�I�v�W�lB	�V���I"A9��5qKof���ЎTИ�n�t�s[0gT�ym�&���tT/H��D'Ͻ����c?��9ő=3KG��_7�ߕ���b�pu�XL�z��%��_��'� ���`=��Q���كنp�=��exb�@�͚�k'�ש������� �"��>��6���Md2�8��P�7*���P�Z�����H�]��}ʫ�&*�us����`�����F�i(Ym�g咹�����{KH���v���]Z�)��@�}=����~���Ȑ�)�E.B]���@���k�,�1Y�]���i"L8�B�p�1(����W�[����	
�o���ƬQ//��^�$w~�w�Po�P��l2�a�Wp�f�Gnm�"\ȍ�~Yr(�`�����甔Е�����M�;&�b~�dVVV��edЪY��H�z��wr�ַɊ%\@.�J�B�c�
ֳ�zQ�o���b�}�}5��5'W�yA�p�3�����O�By�����sm*o����3�-������6��O�ښa�>�E|.N,x���O'	J$$4443���	yLL���L�M���ߊL8➞��.��<>����>�t���LX�/�dh``W���w| Bm���
JK����C'�t?�},0�P^r���)����>��� EژR����M����Skk	��	?�(�?}"ԢˑI�1g5^�ế�-U����[ZZ��ztlV� :�w�خ��<b_�ׯ8WWW
�ډ����/КZY�k%�s��.-/���f``���VbZ,��؜x���A�b�e����R't5�ă_�s
�j�@M��(xd�N�XZ�]�W��ψ۴c캺�N=�D�N`��ğ-t��C�X&�/ϋ݁"`�$�pq��QԾ+��h�HZ�A�����N�D��L9�����{�+f�����VWK��i�W'�q�:�ꃊ�y�<|	�ciW���}1ջ���$0z�P���h���°�#��-�1X���n��{��|oNz��A���V c_Z^�IU�	$㦦�Қ����o��IQ֟�@�WSü.GVWW�'�v�'Iqrs��Aaac�؛)Q�����Ui�(h�yvI��h��V�o�L��ٍ�PoOm�>6"b��^ ��Y�����vM���^�yf��$��T���d�$��>�����������&��*%�2rrH޾�xt��o���S��Ѐ�����������r"+:"&5-�Ï� ��/��Q�ܛ���Z�~	~����nMX�FF��8h}�t��c
�׻��-o��EZ6�jXN��1،*ZZ�Ј8y]]9���Y�۽�Uzu�����.�j�}*��I����<��&sQ+��=l$���j���
i
���i�A��`Z�Ѓ�P��&Bm����&�NC��f�Ln��e�f{V*�,FFF���,T�\�'L�$��k�sR���ll�.vxsx��e{<�S�����U�Y����o������n��@z�i)�Ty�K�l�/q!��W๛�c9�#��GG�&QJ�:���i���{��X8\j�tq1Ljv4[ƻǡ��S�#�:$���l�'��x����@Id�������e%91ሸ}Ƭ� �����{��Ƿ��ɯj���RqE�w:�T@�饥���'��.������L��?��z��4�v��H����x�������d�dI�ǺkT�	ݸClW�R�tMpּ�&z>7]�D��z333����F�K e�w����e�q��5�����ro\�;��^�
&q8���V(�p������a�+5��~��Sw�*PBV��t�����`��,|r%�
)���
�(Q[ L�n���ξ@�K��Q:%��/vEYMu�j�M_����SX�n��m^�6$�Vz�پ?�4 �5Z4H�u�J�댏����a��E�a'����4V�S}�3	N���x�O�� W��X)����*�4$I��:^�.���s���r�^u�jg�а��P:��M���>��<
r��J2�� �`X�'kT?N|e����"��1@����y�A�m� �=�u'vu�"�����u��V�ώr�$ K��17�J6j�4J���	%��%�P"�ؑ��Ά+j�b@oT6L��߁9M���=���]ӥ
�G�C�J���_�u
�?V̡�,��2�}��9�q�x��I I�E৔ AA�S����n�[�㤧R�����>�WI嗹�vEҞ�'H n�֪=��w�v�ӫ<�SѦ�����oU�_��}(���8������+q�����d�\���(f�>��&�,��׷;E�AdJ⻿8��$V���4�GV<	24�h�5�����������f8nAW�!09JF�I��E�C=�4A)�pګϵ��&q�>]��N�d&�+TD��AA�>a�Dj�nQ��5�/׺�+1鷢���2�I�s�S�i�`s�Q��2 �vx�M�D�4�SS�#�n���m�D��/�����I_U:�ն�.��"���O��L��:S��bj�����Z�*�#%e�*M��Pq"H��a��'Lқgk�����㽇?;?��,�,**�����o�3���^�ϵ��s�<�N�1�&]��?��߶�-��B�
��
��:::z��eA��\8&�3�<*��]�5�lv\O���,���}v��K�DYI��*�M���9Ւ��݃^;��WMx��nQn��B��FșE"�v���Ȉ�2�&T�n6Sɞ{	:�����X����Y
^M�k�:�w=�44$�!r��l[֥��'Ä׍Y�xxp=ډ5+�gQ.Ջ���A�4�#���6
ZF,+>=�jFP�0=��j�ۊe�M-2̕A�!n�_�y���\E�c����PUtm�H#�t7�4Hw�Hww#�Jw
H?� ݝ��[�������f�E����=����y_�9�����(���'��C^	7�,�9�
*�#�}�����=A�~)f�~wo	��� xFcd��1i4X�{���Bҹ���aE���>;+**0���#�������ۯ�Á�-���<Ċ�L@}x��d�[�d�kv�x�+�0���ξe�ìL���ӋJ��h�o��љk��.$U2M)$D���n$�]�]�%g. ���^0���w���o���OφYL�cH4�]vg�0�;��x��!�I�|\vv,��C�lel�����P�T����
��)(�%����u|��R�T�2��_!e�L�ld���w9?z(�J��!6W��P@&@�^5:8��i�YYS3̒3��]�E3z͜i,6��?l���qg �G��w@�g��Nk������^$M��+� &r0��V��{Q�GG����A��H���������
�˒VY:��\!����uubA�>5b/��_o���M5U؟6��)LG�B�/�s
խ��G���=���A�㴟+|-�{���r��f���"R�|���}�Ղ"| )]����GM�Vw`��3�e������j����O��[�c�r��z'թb�U�)�Q�A&y򩓣���yf.�����⊆y?2����.�5_��E�[R� ��v�%��怆�4�L1�&#.�T��r��FZ��������G�H�4�^%j�N �$3�˧v?����R�<d�GK~�B��Ġ�d2�rh���f
���|�gh��R�%�����y?�/_��s��e%tGG]j�e�@+$j�c������	�G�T�^�p7O\Y��OPVN��]��IKNzQ�r���!�jl����Ͱ�S@o$�F2�Ȝ�m8���7��ϩhBt�y[I''�E:���^c__�����SS��I����@,w���&$$��kUs96XJ�����[@N�1��I"��X-�UX���e��a_��@����o���oወ���뉹�u�$& |���"��K�<]p,�����`9���;ݖC��x�[Q��Ui, ��r,mA��Y���		Xn��q���b��� �������$�+���Z�7x��W����p��_[2��]c�������}3x9==�⼀� ��<fɇ,���
��17�"�2��߆'Ѐn'��/ވ�ȣ�Ҳ��^������{��϶���f$�>U�_2%h^}[���g�]4ay鳂��XG����f�Q�W*�١On���U'2K��d��2�����r�����
��� D����zܬ�:��������h�.�4��8�$Z�ϖ+����V�-S�0��q��g���ߘ���n���/b2����
﷏���u(K�S��)�)�6K�g���-���2�c��!�1��>`MY�QԤ~A���
n[NNnIj��я���TYBr�������כ���ll��b	�%�;��k:�:��It�1��G�J�z�q���#��4��'0]Weap�����q!d��=f�P_
�jI��26PA�����d>_��B��޽.����� �ƕ�
� 2w�ن��L��V�CnE:��f7?%@ƵT�,��4��S9�����?��Sh��&%%���w�Bfg�f�����C���;n�qq�.���{�m �����HD��{������4`RD+��� e����+��)�(Z@I�c�*A�[b4��e���Y���
t u�xL�C	K(��z-��qhA�}v~������V�b6�����ύ���'?)��N^�Q�>+`�����F�T�hbuw
Y�Q-����B�Ȋ5���i���_̆�31�#s��ΜGR9B���0$0�^���_�x1�����_�R���{l�Z(".2�"����f9��2�zq��_;����Ԍ��'>:eʢ���0���]�7Ԯ����OM��@��5*e�y����u�'3����� �ykDxLY~�ɛ�K/�t.T�����d���\�Ws&'�>� ��uN���>���%

����<-|
8���GKM "? m	خ�~��13�^��:!��������>4�k"%d��:���Mw�d|�����'7�y%%ȿ 
���֬�w.c��P�g�#""�pm4�֊,�sR��f��7ݡ��\T|zz$p&=����L�H��b�E�����;K��HRXٗOp*k�,��N%r_陇�^��f�J�Դl���&��y޶��c({U:�T�B�NC���VVVVcFlX�6�1��^�}QNzE�{�y��sX��.�p���5�Jr�#Snes���}��j�Zޢ��ꏮ����������r8-.g0)p�i��p�Y]EW�V��
'�0�)ۈ��l�|���2p���f@9} S�B���-�7`����~ʒ���B���wɼ��L��XBwL�����O�)�zĉ9n�<�VH>>�/���}W&d���-�[*�2,��9�l�w���c�7����C�Q[{HNK���B�UaQQ����P�,h��zo_��7;y���C�Ð��_U�Z/��b<d�:z�V����3Z�m���@�~�z�3]��/q�7G!���z��`"�G�x�J��B��v&;>Vt *%80�>����l�JlU�" I�6eW���_s�R��&`���ײN���ж�J3C��yY�ۘ�0���4��3s���M�ߠѮb�G;r���|2�|V�M��PKC˾�{/��?"��=o��m~]�f�o7e�-&
���D�\ a���@	Bi�*�]��ӎ���Le�ˌM�!+~�PXu��h���19�Kf�]hh�D0�ܵx�8������*�_�+l��ݬ�����v��@o����{gf�9���cS��1hニ^���ie��=��u�G��Q�빤�cE�O[r~�#dx����
@���lIF�HW�T��ǗODD� rB��'�V���)�L��6 &�kAA��$燽�4Iq�U��(�%85SaC����Y�hP^�ǃ�U���	�+>o�G�>I��_�^)0/o������]��낡bG9X�Ty������ub�rsº.�f4���0��5m ��a�����6xݑ������)xд�����������uy��^zom^M�������F6��Y�6}��N֛��ik
Dhqeb��X��j��P~�PQ
���Z{s�TyKK�_+m�tuR!����)� K@0��`E��؜��ny��l���tg�<�%��s��@tm�/-�M0��A�M&�~d"f+^RÖ�����Dվ��)Ē�D�BRN�%AJ4�T�zI𴵄�"#.�<�T�i����V�Я�,�w!�����	 wy���9�������cM@Q�7N�^Ă���LL�������A���(zm���1a��o�6i�7I2��bw��dMX�~��q�k���C*nn�h��E[5��a��VH��3�R~��& 껂X�uSH;����/�<	�ga��LI�L��BY���f{��$��?��[�zQ�Z�N�S���F`���� �I�� s���
S���L�G�9^f�8��H��u���߹�K�d�AW�=�300(bY�G�B�v]ZZ�5���0��#�)0�Û�d�\n�`�����2d�/?߬k�ԫ��j��i����������0u^r/�/O�卙"Fd�����YQ*4T׫K"�Bs��8ڋ�͘A�Y�_ ��Qy��仺�����+[ȧ����͸8XĂ}�	6��w%���w�K�Ag���z��dq�x� �d]4(���˂��ȫ���^z��y��� 8�D�LE��SH?��5�S�����d�vd�����Q��y�6��:zW��`S1ZLt��!�S9b"�5J)!%@�(�z�(���m�1������?��1I�2��ǟx_�|9_��w�O���s�%Ip��b�XU]���>;j��ʹ5�899�형�k�׺��q�&
謥����}�D�}���ெ�Y��	��|�3�ǳ���0h N"!�@.�����3�-|鞔�\Ǭ���kE�E�Y�s�yPnx*�a�:_��!�?Ԭ�Fv#��ܳ����bїU�i�X��%�))�=i�նM	LqL�)�No?z��-�p\�f�����ZH������ΙĪ��(o�tg�I�)����U�oF�Y�	��kΏ��;���>|T��q3Q���Vay�k��؜�ĕ:ڥ/���q�R��KBM���f#�Ac͑�����&]�[�����OcЭ�FٌÕ���̤Ze��w��kMM������d6����q*�H�}F��_���t�Y�&uankk˰��C�+��'*99��!�-��Mg�<��:�¡�V7�E
�j�6}�Q'��+(�z�LN���=f��}Ԅ �|�֣�]�{��8/�8�嚣�-.��H��'	��O�Q��h/�m�S�=���0����$��e���㎈��C��UIs�hV3?19��ӺIiO����x��^]��Ҁf��ܡ�f�LD�UuNQ�|���%�Mڒj#CC(**�0ɼ�;�f�������֭�j�R�dNyƲlvJ`�Bi����3�ŋ�|tQ3�	XԾ��L[����WLn/ﺼ0y�8tbb�����3<�܃�:d���������-��X�����t��-���$�>]F�mq��ò֏�*;���^����D*4"�v0��ȕ���9n���:9W����X�ۣ�c��t��<m�){�*�ڥH�.s(�T��_�t¿>����a������1�B��S��Q�`���S�`���_�'��1����miii^sQTSCAG�w�V���H߽����Q�!I��"m|xz���¤�^c�Z>�k=f<�Ϫ��0Dٴ���h�ҫ����ˡd�4��iV�}��؛L�,�<�ﯴ�jh����SQA�6�d�ȖS$R�S��A5��������޵+������3�m�������!;^���� %A@y��L���[U	$����nll���MN&�s<!C'R���~�>8(���H�8��p��:�.��m���:�%���1��T��r�a8����5,K&!hk��`��}��;�㯡����欂�1����j���M��l�ܡUUl###���8�]}%�����#��$�p�H�� =�Z���q�#��������Ϸ!��љ������"�۹��$�~rQu�� >�K�s��ߪ��2}���ȶaQ����߶��FF���<����AC#�W/��̔�']����$)	G^I���~�p���m����^������=sckkT�q{�PQ؅����X����7���.������������L�1f*X1��!3G�n��vq}�����CC��È��mR��8�V��o0w�y�6��㱝�=���ᮿ�?�_I�����1-� ��ùi%�c�z2X4:��9��o��mk�Yi }����l)�ig����� �m ��|yEEc{��[`~���]\]w˷k�e������ԝ^�b&�ڦ���
=�I2��]Z-��}h���=v%HDx8�������{�8'aoO,.�p���>!a�jEG��Waò�Y�M�K��z!�4���$�������^'m��B�{���rM��ni���rxSO���-��!E9�c�b\;EL3���z�'��Z�]xy������x�������pw6nzzZy���PX�=��S��sm����{06�r���T�N���~�-!:�".mr)�e���� !������h� �����_2d��xz ���9_��z���"w&sќ���響�T������i�ׯe���K�Da=�1�fER�E�t�>K���&�0�N�$��=���u������J�a�[�}Kcd�ٮ��ba�P�
������|���@43�l��N Qg>-.n\Fn��ȑ���U@@��bǭ�������[}D@NN�]��45���u�A �d�45+;;%��tB�ؘbm}}��+�o%��������j��z���60�U���#Zɐ�����e���֢�?��^w"�-]̉'M�D���򵷔2�-�b�c��g��D�ށ)/�s~���ˍ�/&B���,�Bq"�c�}mm�^5�cRY�oZ�����no�݃Q�xK��	B	r���`L��!��1�����	F�ƌ��ܖ�-_n�������������>����d
�.�2�bK� �����аbaa���y���]III�>�2>�9�HOO�L#Ď:ex���ki<�B����0�fB�z�:�?t�籷 U(k��l���F��ua�����k"��M3��O�x�sһ�bo��<Vx�`�7��F�F��
�����������B��V)��pǣT����w�2_���=���]���:��m���R__�����*��pK��@���	�s2l,N�	��Bg���AX ����V�t���%�A��U�{ֳ�r}vD�JQ�����;�x�8MGD�չen�W�C9V���J���)�P_"�Mw��h���z���1"?ޱ�]$y!@���0j����{F�*�_��b��_&uڐ��2QY�`Q�ں:��s �;y�3���@�m�g��1�j�,C��`2���\��#mԜd���댜����fZ}`zK�����W��߫F�N�\�}�]x��{z\��#�U|L��|���X�7�cT�o�T7�%�V���L���g��M��[�b`-ǟ5��(����Ę�p�3t9K��Gv�[ۜ�E�k$�:��� ��u��,��&'�� �-�:��J��X:jۡ���qj<?�.�rbo���p�.���Fʏ���/�����]�c(m>kx#Z���n0�"l��m>|ʔa@��o~Jed��o͗4�z��tԸCX@U�n��8�n�^��d"��MD$�F�x���i2�����(���[*!������� �ҫ�>�ը��ץ�|����j3��b���Է���K<6�\�8,��sIB�ׅ54f��o}H�����ծ ��#=�V�lVM|<��{5���#����ds)��%�U_���U�n��7���q9���.m���h�1ޗ�rE���R4��ei �\vm����w��)f���^	(MH�=�V9�4PR�x�RY{��h�'�~��@�ÅT7����δz��9�38��i,/m�^�G��*��XK�R����γD�u�'���N�[�4P���ҰHL�A/JI!d��c�,�}�ik�/���.�T���W�mʦ׸����q��e�H��An����_A2�$g�b �`�ڞ��� ]h��+)���1��J���`���iќ/�X�Ä���l�����e��&�flԠ���	�-�س�t}���{����[�e`�����d\M%F�4�m���|O���ս�wKt`�3����g�s���?Nz������|��gU�9�h���+a��j��x�||�����*S��]����98(���3�ӎ\�a35���'%%�)8���[XX�Q�ݕ00XM���sGKa1(W�d7�����4N�R��9�[�v�vΗ�@�����7�^�B-ˋ�m�42!��.4'J����`�u��t�k�vrr:�8����F [���W�Xʏ)���(�8��r��tk!�4�z�A�ǧ�1���)��$R#������2��hO���i��˻�&&�f�߫���Ĉ������;/�_pyA��İi7ope\�鮦TP�2�P丶�}��:z�9��0;^p�M�f1`���9���`33@�;��26�{�v�t�'`�B�WU$��75}0e'���Z�q�򎃡^�����B�*��(�*My�(dXh�2����x����'nԉ�u�ެ�K�D)�-��@���|��,B>��'� �:�mғ(+m��Wr��3���$�����E��uR���X:�a��f��:f��p%����>���U�k��]��N����v��G4Ğ�y��J�����ˌP1�����f�t���
���III�oa�\Q'|ޮ��f/��462F5�
B�kB""�*Mq)�I�jG�z��?z2� �y��� �á�f�r�疸������y~�J�!<���N=*xKDbY��-�0i�\-8	�t�m��iG�	-mھ�Gt#�R|_���9���hN��w��EEV�C6L�(�M�0���Y��~�	���T����L�%�7����6e8�E�`�K���GGG;%�E�t��)9'3�o�f2���.���f5���e��U_���C�����ϝ���<�b����I�`��?u��n�B\���6(8��VZU�ɕ�
��F�C]�9E�7 /1.�E&`z&Tب�h#[�Ґ��~�{4�;┘����i xI��B��6w۩IWǞ���f�QS_���xN�&���!%.U�7���8S �ì�TP�=Mv�אoidN�ت �|�Y��h��h`r^������"��w�e�1��B��p
�6Z�c��d���[�ܮl�|1sK՗��	�OU������&���g��K���������ˋ���70�a�P���[e���*���ҝ�+��~�2`���1��Fuw7*��s�Z���4����>W*�\�<���\���A���̞�32�
�u����ť�2@�H�����K��5�e|0	�"1��ćM2#Xwį�Di�8]!�6������a�,�z��J�ͷ����kˡX:��SB��B�^B�z�^3��`[�h�D��{� S�f�����H[�w�v�O��� b�_.�����c��u��"��HoV�����E/`������x'  �9�b]R<�mW�7����o ���5	n��xS�p��������v���B�g���S1��khP��Mz.��*��]��
.Q͛�*kj�Г� ����e#����xKL��%�t9w�a�-~�u�E�}}���GW��� ��������#nx3nв��A�ǧ��ůc�kn;	ku���>�������,a	JQb^�UT�	�&�wp��:�L�=��j�U�D��X��m$���8~��3��P__��i��L�Ï��q��-g�yQ|�T���<��<9�*&]�[��$��A��9}�;h�K_ۃ\����XZ[��/��wQM_=�?;���i�����513�^V=;	t��O�YL���o�:�꣟�&�M��rSu�/�j�n�,�<�4�5a���n�v�A3x���e�R����RQ=�W��f��2ee�6ېX�������q&��̞��g�8p ļ���V2��8��Ҵa��`�6�$$$8d���~H�..
����'�FpO�!irs�
���.x�~�AX7����O/!%�I����Q�7ȶ��D�ԅ�75����6
;Ǩ����:#C��^ ��e�[�S���w�6ݙ�o5��	0R�I�{��G����;�^6=KPc}]<,ߙ��b�W�����X �q�S"g͢�:7ED.h'�y���(	=��N�A�֞��i�=y݌�`�dg��� �*��:yH�O��Y������	1^��h��ݽE�d�W=x�����u�6T�z�1�H��s�J�~C����F7��N�)��w@^�� �
n��8��ISC��A�,Ƴ6��|�����(���s��]��H�x�yC(��(_Gd��j���Lj���h�u��2��X(+��tL�����؍V6�ޫ04���4�=�Q����A���B��h�U3�=ˢ	�Ѓ�4{/�A�!;��J*b���5�6J�Al���P�~Vo8ߥh�'��O顄Nky�J^%jo�L�*}��6�EFF"�D58����ǻ���%--�Ν��)�>���m���ЃBDs"D�N|!�<3�pvK��9May�	�k�-yG����Z�a����(���
�I���="w�Nt���M6Yˑ�]�HJ�����lo�09TvEu��J��N��������$z�,��?ZZ1=3�qzYL�����ܽ.�PK:!Rz`t����f͎�I&�laC	X�vh����h�In~���U��2%ު�8�������YWW���rKX��:p�(�ޖߎ�Vv=��q�ˊ ��P�n������J��0w�<��	�&��ÏNg�L�r��ݿh��������;��W��bE���5#��z[QUuIKO��|�jGT���6����C�c"b�HI˝��)�=�n�����I�H�}�n��
��~G)��P��8���e��T~OPTiRU�0.�P����T��1�-d�A-��y�	�SX���ˏ7�s�<V��%�[��}R�%�M�S��)�_ȌP��aLg��_9%IG;�H�W8�c.���Y���
ΥRE��SA���**l�\(�$F��Pl�׫���u��ܯ@[mw�*���s�n R���<��[j�Z���3�:�w����<j�-�r�\h��_�
��`LNI��/$�g��I��-�0��w�`���A���oHr��rNl�/�Z����9��arj�J��@v}o;"X��s��6i��7����;6����z�;�.�o�~?�������*K.�RoD�\�?�P?뾯O �O���ZTT��E���DPA���Ȓ�,�m���V�ۯ��T|���w_�&��S���ӑx8<cGڬjM��3~R�m��I��2D9��]R����kf��Qx�	ǐ����qqs�n��;��� C�����H<0F�4XHԉ2���wJ�**Sp׽�/����o����(�_%7!��ج^�!f^Y����!o�� ����+��'6<l-R.�쯘,D�\]��Uc�j���Ք��0X����*��5�l��U�̆�m޺7�:�,��r�������,�z��C�4�XX�d��}o��<������]|k�É��3���kLL��x@��@�m��������a��###s�0� ss��l����v��'�%���,蠑�t.6�ֶɞhL���9S^��<��:i�`SRRs�� XJ#BBB.s��ῃ�Q\ݙ�����m`1h/UN[��yCz��-�԰^Y�%���x�xc�q
�����t���v���̕�[o-��&���g�!��vxC��`�8�'1a�+ܖW������Ҍʊ*}����7pDF�+*�x�2�!����}m�R�:����c�M8"� ��Ɲ��Gٍ�*��cO����-��)&s3���X`�۵b'����;�!Wt����Л��X�2����:]-Qn����������"����Ů��ON��9��i8t(�;z��+.���&��PR�vd9��4�B<C�-���y���Q�j��F�'�8�{=dy7��V��?xuܣ������w8����>�h5 �S�F�Q� 3 �+١W5k�E+2=���-�L�l�1ev5��GkӇ�Z�����/�Ԋ�����{]�C���]U��z�٥[�/���+�h1J^���9-��GFPT�̪9;E>���"J(Ǎo�r��]g8�������-��M@OT�]�7�4��Tc��y�mw����s��YA�鸚�+ҹ��͒�6�ڲ��O�&	/�%M�[��c��Ԥ:��k�6��o�Ȕ��!��!k�'$���;]�¤L@�e�d+���L�	F�F~K�������1e��Ъ�&�7j�ٗb�đ'
9ˏ��/,�+T�x-'�o#��f৑��s77�n�?Z�8��Ԅ�2h��j4�t��Z(��l_�#_��FUa��ᗯ�:jq?x���7�w�5>.��d�1���-�fe��%"����2 kj+�F�z��G�Ј
�`2�������Ă��ׄ�-�v�'P!CFFUK'�+���GR�T	��5A�<#��j�#�%���WPߕ>8�v�j"��uI��j8�`u�^���	A���cK��|@ j�3�q�W��Iv3Y��
z�>����>�Cgv��zM�*��'b�P7������Qj�9��d�wrʺ�'�c�ٿ�m�ͷ���I�H�c�ծ	rr�0�d�RSP
���0�k3m���ќ����fщ�s�]v��e��MQx&F��AD����B�5
y�uǆr}��a29�|x���٢;�i[��@M(��/�H�ZwkE2�;-����ٯ�e��p�3�\�f�!�ݭ���q"ɦ);�n�	�>�5l��-�G�?3�p�������#,�����2C�_����l�QL���Ti>ɣI &b�(!]	n����a#�t篳�m~��/:ٳA���o��3�ō�T2��q�	Z�_��P�Kt�����%�~�k��5ǯ.<~r~����o@^�o"Y��|�մP�v����Ӗ.T��$+*&&d�驝���x����\���=��mF�ںu�����"���Ðik����]�tYO��/���+���p��
�:�z���d{�?���	1�I��?�Z*��c��q0���NK��A�7�T8����q綁wgF/��qz3�XO'%e���=/�#B���e��çnw��S���Iq�X_Q�[s��`"s7vH#��5�`;V�h��PVЩz�Ҿic�@�m�y� �P1���~l]����%���z��ʺ�����t��]�i�����	���.���8���}}p^���W��҂7wv�i����p���J����H�����+�^��L���
��k�!?��.*�<�2����M5柹�A.��UfV��S� æ2��[V�Eǔ��H�=ќ�¼v����CH��f�G�6�+5Qng2]��sS�t��l�L��u�X���?|�ן���@{:��wԴ�_��RZ����!�{׶���|�j5_��Ӊ��C$��*�[�$G�d��@�PP�14}��L�X��1|��d�z5�Rz,dU�fC	��_�}�I�D��0oN��LL�p�Rt�\�c��Ƣ���~�~3���xI�=��{�4[K\����y��y���J��e�H�ԛ��N��6<ȁ���˲���TRar�>8o`^V����9�`��6'���>��&]����g�q�7k���K�X�Ǜ��D0�.rC�ʹ�����1��_k���u�=,��ύR�~�J��J�4�YHS��Ap!��a�h��[�����"�{y	q��&�gv?�F�Gݯu$E��@��U-V.�i�U�)���I�"_�7�+w��=�
���j�F���;���8���V���Q�06��rxZf]q�E�����^�	�8D޸~�%~�]��Q�e���݋�A�>|�Gcu�c�˜���8��b�u�v��ޯ���c�8�~���y��D� n�u�1�+����u��Y�1Q���Mn�Z�6���BX�B��������˱J�k�~���c�>�����ƙ8��&������TXƈ ���'
��u��$�h럵0O�fRl�f�?L��QQR.dPy�-®|�@C� {G�O��'�oǙ��KR�^?%<t,}D��ߣ/Y�`��쟍��^d����seDL�Y�
]�!���y�n�D�p	��ԏ
�Yqs��j�����)o0�w=��� xk�Z�	��5���\4ܵ?�?�%���&4,�U�ʳ���8#y_ȋ&�����:�:�w@�ԅd(R7;��ߜ3.`N'�޴=�'r�``�f
<�;ޒi�V�㺅�|��4CF�P���aW��oh��Q\�,D�:�Ŀ2��|7*Ե7�Ã���IEk�v�t����$8�+�����*�MwsX���8m�h������=��hx�	�F�0;1��`lU�Xݷ�SטB��k�r�� @|Ο�pS���xe%P�L��yF�X���P����x�#���y�s���HxX�SO��a�/ޘ o��k8f���K�OF���\���H�;�jx� �i���{R�"����� >�uv��%�Sj���'E��5�X�?}��4�h���s��onf4�1��}�ip��e�i,�|��5͝�P��<dl�����9����g�R�]w�n�6}�?��nH����~���'�y�.J���e⼱���~��Y͕�����DZ�	��c��}��?h/7�$"2��I�f�����u�w�~>�S�g�R�8Ͱ�u>'��u�O��dVd��(��x�ܷ�z���k����}��Q�x� �@�~�Þ�^t��a|�"u=3����W����c�<����Zg&3͹mc�=��X@KL�
Rk�)E�aw"�B�6�Y��O)G/	��˚����ݏ&��+����lŕ��@]��K��i��A���ë����R�ׯo֞O�n:-����Ou�{V�Nq%G��W@��+�T�0�x3��;�ӈ\Di1qq�м�����`lg'�Z۞v�m<�^R0�'fC#F0��]�[�%��O5o�p�X����:s,y�����b^��VK�i����)�?�	:�.d��B��#{Ir�dq�o���zD>��,ɕIR�66�b�-��z@25�_"g����n\�j,�oTH�~��a�2�`��3�N�q[����*���=3�������)0[�ŧ>
$��3?b�VO����B�3"�[�úp���`L�e4"�б��co&�����B,&vd�:�ZR�72|d���$�H�C���-�l����1ÿg.wW��<L|޹(���J`�7��L's�Cn�
��>��S�9=��T�]����K�zMن�" C��ޮ;������H�F9m�V�nQ�=�jZ��)��1y#9�P�V�0IH�n��ν�D��z�G��fhoF���z�T��0����z�RS�Tj2ƙ�� {����h_��������������_d-�j:��CeX�.%^��� �"1F���N��kժԼ�����>iĭ�p����|#��D�Ƴ�]Ei�����Z<��J��Q���V\�x(M��rw�D�U��?�?p�ƯJ�,�����'jwMr�'T���r��[Y�K����@;�x!C%���3��,<H�/t�H��F�DX'����wx� ۪�%˙3��k:�1��#���|hE�kE�F��XU�};����%*H�K
��l�BV���b������������z3�C�g�q��"=o��a���:�� �o9Zrl$��8^ߎ�Y�c�>�z<2\��?����g�r%b��<�������nm��yI�dU�g;cn�j�vC>m^��MH�����F�9�az�тH�~s��ȝ��kF@m�d�GR1���nA����9
��|�\������}:^R����t1��kg�A[�J��P��+M�4y����q�|gF�:�Y@���Bv��M��q�^�xU��H|���5��F��|�c���j��ֻd�󴌎�ΐ'����t�^m��;�.�D�2e�B&ZKLu�R�v��I�H���Yn�Dd�y
�TW.�]l���&P�T�q��������Ǥ��;�(X�L�tR�7�g�y|�_x��jk.���s�X�v!h3���?��`�m���ܵ5W�*I�a��� �X�� ��┺o���Z$�ȋ����-~�r�5#�"�ᑊ0������#9�x!���VI�ww{A@���?ګ�+���70��:�{���Ur'��~��MM����|$�YT�|�L##�3��YL�q�s$���H����)��J-�b�u�����?�<f�:�u�ל�y�K�.t��"8�����ƭ-*|o�&��C�D͐p�ja�Y���`�a��&����|p��͵�LYr��J!������޹���uz��1OzBa�Ec��+�`��&�ۘ�9O�+p�e$���j�I8�1<+)"`P!��zW�>%!��ջ�^{i�
ڽzg��w�Q�6��+�̾�yZ��n��u)�E���S��S�I$Tfq�暿��=���V��Qe1�
�5�x���?h��?�-��]w���8�n2l��M�l�[�=���o[K��Ǥg��A"ܿg�����:5����w�����x�U2��51Z�nDѯ�\EV��e{<�Y���h��x�U߭�-��_���KB
�oݑ�z�)}�a1��WB��πcHM��� �z�c�A,��*����3�j��A]� ��2�2#�����"d���g߸3���0��S	0�e��q]ϴc���h�ve��_=�&�*��
y�cذ��[YYI�A[��aaf��)5z|��"Z�{\� a�/>���T�1�z3��9�>�yT�Vnc��z}y�v��T-��_@l/��s��z��E��݉��f�V�,�0wE��-�r�e�����2�m�Q�<���& ��R`�E���ڿ�b��3_�c����k�� �{�H��e�u]ڟ�m��0 ��+�^�,�YR���i͉[��´"�%鿸AN���;�Z�|8,�U��Z�L�צc��,]�6S��	�G^���ǞJ�^��l���ޏ�-�1@	KI���6�leV�?pk��g(Guuq���=9Sލ(��ɷ
<3�����`����1�Cb�����a�+R2o7�����\U���^��>�uz�zM�s��YZ[ce����˟�)�����@�q��
���j�t������=��b�O��n-ߧ���J�� ;X,l��ʹ��59�}��E������"�^Bj�[qq�|\ӂ�ӂ��B禥�cD�#c��6��F��V���=1h���@�eG�ύEf�����]�۱�"��@�P�aꫪ0��#Xq��ԇ��sr%X���(����+C��E�%�6z]��_C�{�I�|��E��2�Ņ��a��㗾i��^c9�HP�M�ЉIOZ}�����z�g�V)����>��#�`=�V���5�&�������Ȧ�����'����]`Z0�������pѓ��MWE��Q^A)_���$�nT@:���^Td)����YAai�k��]b�X����{�0s�����>w�73�S�Ҫ�y����Z�a��%7�#�"NV��c  �9���;J	�F�	;cp�Ũ�(�\����*��BtW7��Ãy���_>���Nfީ�}&n91�RO�D��X
l��zo���u޿�zH��ó@��|�I��
�M�B�ę�i�A��8/��?j����Hb)�%���bBҼL�﹠ ��=���@7����H�9�=�8�������V�����{�eԝ���D�=*R�`��sqV,��Cy���gU����&JWL����Z<�5�Ȩ�h6���^)))����p���FUn�Y���k]A�޽t{x����j��ШY�Y��}���vh������m��6]���ӺzXR���Iд��Yk���4aXڷBB�&Z�����!;����_����üX�����n��x���'���"���ʝ��@��*u8�i�:���E<�}�&k�T�,�%J�ȫ���Q2�fZ�ߋ��t}<��ochZ/�4�K|��fV���]��_ ����{	K�O��Q"�G7v�&ǡ��N�e��~��kl��:�M������V^^�R�=�G�+���jq�%F�璈���Gv1$(=3"��Y��_�� E�O]L�f�(��Wn�����gj%��~�pf�H�u��!�)�a}��Ƈ�yi*=�J�co������Ѭ^�*_����R o_%�6@pK�Yu$`�	}C�W�8��,�J�W�Z�ז��z���.���2���]lG��7��E�	���/x���wLM��I�jz�p��r���.=�;�\����?����v�݄��{#�.� �D �.ꅌCR�9^�H2�?u�J2��D�_Y��,,�B�*r�"�_K�G��M��$��\B2����?���NP��-����"�gvvv�]��+�$ $����#d��*B�x����5�<�.���#��]����iz���CKVAޕ{]��lw�	�����G�'�C��<�������Y�����-[�C�"�/�?WW�i�����.MƸ�Y��h��sYbl�߫��`�B�j�q�w\���W�@o�]������r��@nalj��Ζ�]#��[�zkǄ������60:( ����
���{�0y
N-�f(A���J� �M?84q�WhH]%�������	)��|�t�!ã��>n>T�#�ت�� �8���k{��<������x�˾���5����7R�n�8z0��
`��X!ϙ&�ht8��ߍ)@m�@^�=E�2�lɣI)+
��^OW [����;�"���Z	������F�0��gm�#s{:TV�[�>�a ���U�0�yc��Ek�g���:���,���<E�<��^#{lfk�Nv���D"W���O9��!�HA%���Iu��	q�6�G�3D.�����|���C��8�~l�d�w�֨������xz���Z{��t �_�`挩-q�B����i%}@������ݨB�V������4K���i�7d�Uf_-Z5�gU�u/H�n��z��8����ItԌ����s���Y�^����6ڿw��n�X����J��f �����߆�gQ�5%jh�X]�_d���O"U���l`���2h1�td��V�Z��\�o�0L��}"���S9���X��!�}m�x����Ui|ä�;*�{�l�����Y����wת��+!�|zz�|��d4�P09yKEs`�_d,�s� �WWl��� �� �{���UUj $�����8�������Qˎg�x`�����ۧZ���-8Q9܃�44��)��������f

������l~�S�`�ANG��-�y��@ �%0J�[�����ٽ��,�m�T��	z����Jj���Y�h�m3�8�����Je>��-�o�|Z�6�����Atξ˯߁/'�����v�ǚ��p�#�=_�ϓh�8�dG! e�{&N48��߻@��{-�v��p��-7�x!��t���lLޙ-\��E��ў���\�Q��&y�'��B����CBd��L?�������2���z~����։��"�����b� ���B�|AAA�FZ��m�@UR�m��N�I"��~N�+n�˙���?J3�;�ŝ��/� �Iޝ�'�jZ�R����Pֺ��$�@Y�kS*U!E;���I�b���0w���%���<�d�>>"ݫ߁�y�����쳘\�(Y�m�27��� ����"�N~쁀.��$���
 �����'k����w�RB˾++���۞o?�A�������}:��u���뻿8�;�F�}C��0BG�� ��.��0F\%�*%|�	�$<�@now��t�c�H96!a�$��T��v&��8 �jeN;2�hc���yt�˽��]��#�������P�n�N_����6��MtΜ��"7������丂b�/�5�w�s�ZS��	HJWW>^�v #�WWW��j����Ғ�},}6�@�)j�f�|j��Vxs���Qt.��O��� k)�>������Vu�͜�0�j���u<{���BL�ɸ-Pܙ�z����yMg�F���_�>���\�2J��m�_�0k?����T���bv4����N��靃F���Z�c듛�4���R�_͛�s�G'c��l�*�N�ep��>w� W=�/�_����"����III�99�Ӈ�0�>h�\�Iin�Rg3m�`���=Vr��]C���3L���}0�d�����6 �~u�������kwX=:D>u���F���N)�L���� f��J��(j�m�WJ��0�����O�Rlű��yB����Ro�b�h���rvy���Bmz��" C�m�mO�H$��S��/���?�+��Q:�l�di�~�� �yR�˥;� ��M�ƙT ����?b��/V�B
d�4O���������h}_/] �))�Y�4M���V����KR���:�	0Ab<�҆s!%h��eb����eD�����zOrd.
�"W\�����x}uQ�ڊ�cаr�Ҍ'{����n��]�-�ȡ�S���ߊ�����̀��I�i�f�pzK����/_Tm_�ݷ����e���=a{7O-�]��y5�6�������c�ޞ�//�B �c/Uh(�ߣ�/����`r�q�)~�U����b��Ʒq�MpN���L'v����*�`�h$�CV�c^�ʗJ�������T���z�b&K6m�f�&K�a��GnO&l�#g�~�P%�<�tM��C,a�}�p�=�)` i>�]=�SxRN|q�'++
T�;@��W\�/�S�6$�
�͙���R��{l'�o����2�l,A>�+޲�҅+S����-��C��e�_�V���A���d�~ٯ��$pd�m@
Z���ҧ��%��5�8�h�j�/���Rn���]8��c$z�QBeQC
|͘iP�է��o�6߄qt�!Y���u�B�>b��"��_ �ɿ�zO#�"�F�9�UF:�5������벷��I	Ɩ���:�-_���y�"��W0�˳�1��f/�r��ܷ5[sd�HOKT-a�;sy�}`���g㬧1dY���G�!�/�<�m��'�"�R_f]C,8�!!����֙��~{G4W��}A� ���������o9͍w�:/&�{��r�ZeI�����g�ia��xn;���x��\�:0!�2~Ϭ���N� �����TڬjwX�O�3�F����j��>?hlh`J����~�qA'y--~G���_�9p��%ܲ�ǟa�]�,
�)�D��𒵤`��RK��8���qF0C��������Am�b���|��L3U�#���N�[�(g�Χ{9t�
h�)-����?�>K�O��>��n��j�\��E�uKWt��2<ti+&eƘ�ރR�+���l���I��~��4[��ݽ#[�&F��.@��ڑ�/m;A��+�#�F���\�[�՘�V�k�~�H�ߥ,��h���h�72��H�TE�NA;��4��/g��-K��x�oF�{ݚ��`�E���n����3��Ds����l�����?������dT�n%{�>���4�j&˧�7�[�=�Sa��m-}}@���&J�������T<N����a����G��[�.f|����^��L�8X�В�Z�c�f��x�j+�^�t1�`�&�0�}�3޶O��Ғ7�5��ֆ���mo6tOO��(j|,C�4��uOk��/�\�K˨���g]���d��B�Z�������n��}9e`+6��z�&����%��R�8�0g��oH���Ѕ�E[�	���#ww����s���'7��9
����!
ڥ��!9X�k��^�>��$1����t�f�J��A6�K�H����-~��2u�rڵ���DqS*��c��r�����R��
x�ĺ��x�)@vp�Pn���P�Nee�-j��t(N#.z��\3W��lDj�it<��BKѵHu�Z�o746����e����FX��]6��:}���o���G��&i|��Nͼ�x���J;s�\��ټ3�Lҗ?��Q��WD_�6n���z��v,$x:c��"M+}�q��O�4�>|Ɇ�c[�^Řh��� ���Ͼ��ʡ�m=�7>�ĮRK_��"j�5����dw9K��������͗C��K��ܸ=�͉\W�}�]E�3��#ˬ�!������7�"�d�%!��!ޣ���E����g�"�0�I��V�5�*/����RA��;�))�?����(w��P[��_?�5��r�K�!�ǃ�z*��ʍ�29+PJ�ez&{�X%�Ú�����2mM�����	��5�Wg@H�H4�0�����_9׏�f߄Oj�9�h����
��I��nND��6����_��?�ʑԇP]$"��"��Y�ْ�� 8�٧1ɸ�hj\��}�:�)� �u�5��y`5&���42�0Č��������g��5�]����%�6V����*qc�O�5l��c�Q���Ֆ<粎4�6������4t��
�XR��_Zj�~��a�վ|���f���y�|�f&ʹ��?����nΉ�P����_�T��|�H�%5+�1y���H��\��#QS�}D\k���Z�2��|��W)6b}��kr������Z�>k0�)��3g�*���|˰��=������𹊑���B�;j���״[;m���s���W�����P9z9��s��XƎ�f�l�c���`.�=j"Md�2��J�C_��ϒ��~�d�G�b�n���쬝8�fC�YMu�6��r�)�J�יF�ffv����`�Y�o>-����vQ�~�E��cmx>`��|�a	�R�p`/�#p�a�E���մ�?����Jx,Co�~�����q�X��@�O��HHُ4~C���y__�@&J:�m�c4F���(0_g%�w1��V?��q���V#8��	4b�i2=?�,��;���ڤ=��<�?,ϻ��=�I��r� *{]��6骽f|�o9���,~lu�7	���zSXK��4��m�渊��DOטḱ_�	�
�q���[?�7���q��P�u/��X��2�Y� #c]���jS�	?���7L�X��J�.$5��[Pi̞�� (�oR����D�1��<G",�p�С<�er�ySY\��[(���^L$@
2���>������ȼ��P��sj\��a�fw�;Q��m�$��v
��%'v�����f���tHR��h3I�އ���5ax��������Z��e�;�e��G�x��ֆF����P2Fi'q�CUG�
#cm*��I1������
����Y�^< ��H��)�f:;1�M>��Y���ۙQ���/�vm�Uҹ&��g�D@\ɯVc�gg|��m6��}֓�rBCn��Ø����g��#,�Y��V��2J8�����֨/�Ն��힧f4�1�̇��g�����_t?2�Qw�Ӑ�>cs%��gmm=��^�{�	�� �T�ܼf��9��Ó��*N.��l� ��4�V���z�;�����v]S煵�Vlh���Yj�{���ljF�M&*[:����+� ��բ���J�I��ѥ��A�~_`2|�����X�b��snm2�2�l�r	Kz63.Fq�c["���4��{q_H@m;BC�� /.-4��\�u���g�֬�+���T{u}��a� :r��	
�/�j�얗�gΛ�_�A	�lN>�`���ٺpڈxɔ�IccZ��K���b�sړc�`
�0�Á%�J���b�ŭR��S�܉a�����MU�H@���rg���Q?�94{Qē�����*z]qt�v��I��B>�wkÓ6�21H����t)[y���K/�SSӬ�ݹ�6�l��v��t	�R<���"ǚ=	Ю�9�E�t�z�� �m�ꏷ��t��[a%�z:�*�$bDA���fٺ������(ZH�y�iru�U�V�cF�1�1�+|R��W��-f�r�rt,����q��o��>��K`9�0�,?�5��K��a�(b"��v�c�W�ߟ[����oW<[x�����,���G2�Y_���?����|K�*a��ʮl�8����<�p��n9��o�zl��!�e?I��)�h����"�
*T���h�_7���e�j���ǂ�xQ]�1��=�-��f��,?��ބo�ױň��&%%�<�/UM���L��@�[pe*��Cph�hyEE#0����O�Ǳ1�*8�T�jkOl�ӿ3:�}�ߚn%��d�^���O3O�v�qE�ë$�����deS�-�[Xy�u�ܦ���cډ#��_.F⦷rT��G.���*ǣ�����h?J���`��^�-+z��Z��|�m�:����q+#���y��4g]^S3��I���
�$� �k߇�gd�)�z.�z2����y^x8A�a���x�w ��[8�%I�m�j�흆Ѓ-S���J��%�?�}=W����MtV;�תB1�g����FbP-}3��nѴ�w-&��5����u���{O�|�#S��~1���*Gu2"�@���TU:D~:6�rf|<p�(��u>y5PN��¥UUj�}[h�
�ͻ�-�n�;�� ����n������PI(���?/Pe	�(�}��Q�_�vE���ϱ<y$[�z2؂[���Z%w��k~�^�����a����W�`3IF�od"�=�WS� �m2N�Q��Qv��$��؂���H<<����0���/�x��^�w;[ {��{o�*����Ɉ��^{v����7@���͢������*�f#�����?��@\g���Lx����wS`�Ķa:dK�G��~W]� :�鉶��߃�����k���qDw���e���YD��a�烬����#ځ�ߦ��6�oF����?�b!�eYb]����ɷ0��>(v8g��B�t�c��5c����-3y|!�ŚV�d��o��avf**+����
++Ui��~c�������Q�EŖ�xސ�����R��D��?���qҪ�Q� u�ew����^�9��d �s6�$�~8��[󙹬"�$���?6���Lr�4�@'���U�۝��~�� �AX�2�>��<����D�9��2���e!^�v89����/4��ae(�T�8999�Ī��l�����de��n9ح�[X��WfOxzT��7�ӧ_�Ѧ�o$�_l~�<���B^ "*���&FmOki>jr���]��@X����Tg5�����Ah�D�������kĜ�?��v�9��JU�Sw����_	�a>�&5 Ky��t�*s���F����Qxxx��af�� ����W����:��"8�Ƭ��ٴ,���e������M�WV����֖Ӄ�3H;[�uKہsUaU���H|W�8�����C�+גu��۞h���@l'�,8�ғ��u�~�Q����:x
�!_���ބ7��WLrL7��e���`g�z�����|P���-!��[�a����J� HɡS6��l����qA��X����^�f4��hb뢪�]��Njų�t͛r��ٹ(i��(z�V��!a�d���er;\H�*~�CR�~
ɤ#|yY��]	�������4)-r'�%.�ֶ9�{8�Y��J`��[>�j
�!��"�����,��vF�����^��bA��x�D���Qx��G�z��a�i.n|�n]o��P���u��bvt�pHy>9�A�����_}_;d��������e�������D^�|�R/5�f���YXE*z�%^$�VK��!���t�L V�h|�<��)x%l���~�[u�3.#�QW"C�H���@22uK�C���-�'1��ݜ�){
��vmoV�ğ���$��h��FCd��q�{(b�]�KGjq:?�w�ݬdg#AC�����P���-�lV��U��G���� ���'���2��C��D5`Վ���W��A5o&"���G�a���sBiI�PD�ۇ�+Y�\e�EJ���mo�7�E�f.��75��S�U��W�mn1z~�ϡ���D�2�Ў+��ڙ*�
��R)�b��b�Y�HdgWڗ��T\ʟ�싕W�ị�J��bs2Ӹ��&]bJ$��X�GU��|�؎����f��wrj-A�qj���-��
�͞�����F����M��KC����>'���ފ���� �y����z�l�����o2��	k�������j�z	Fz�I� ���(�D:c�yp�oz⇹׫�b�(�1���`�N����F�A;_���S����!1e|�-�^�#0���#�޼�Mқ�*�Ma�70Sl���7͔��m�7�vX�ǜ�>͸
���w1��i*�<�:T��@`�1�e�)g25�l!��O�V�7�9l0e��U���ym�d|s��
�EZ���^�3uޓR=Q��X�5n �Oo��up��ƿ�w弆`c.*�o
�I��6��T�B�潋��F������^��6���Z�&<���3��v�mr�`I��r���Z��J��;�gj��-�6)(�}�j)���_o��y �u��%-J���V9>��0lrM�����4F�cj�t4WӕTV$Oߗ � ��m���S��f�oi6�9�<^��T��U��T��8�`_� '����]�����bs�
���u76�/1�o��f��|�q8�����2��sw�۟=Y!�k�Uzs�w�1��9������\���hS�B�uS����=��o�T,͐����F�;xl,�r*C[oa�k���1�d�ū�E��;^����[��ˌ�Պ[�R�#&��}�9;�Ce���P[�W��������������nN�(�7	y^��y���������f���ټ-����e?�Eܺ��L�R�&k���EX�Ұ+�D�aYJ�Lg�B�gC��m Y��9{i.�.�ٙ1-�������ؓ���|i��5}�}���@[�ve�a���ٟ�t�1V���,��t��c��"5��5�n18�z�=��X���k:��/^ v����?~lh�>@u�de��������E��%�Z���f�,VF�fv�WH薲�X��B1��~�{����v��kja�`å���fe8����b�u55�|>B�HǺL��|�s�8�f�أ��9R-�8>��ٲ߼���J�j]��3"5�\70��R����L[.x-,w��zZ�l:/�����v��l�)��^F������dd�p:��F��n�jX� {��1��`}"�E{}j�_v����H`�q�V��\�(���3H��Y�YZ,9�R�պ9=��_��q�*�tW.�c��Z@��!_����ĖOE�.hY��]�>���H�cB��b��z�')��(Y1a\tT�ű;}�ps�����I׭��>�e�����5aүV���v�Ћ�=���]�������Vml�H�*
�T��#s@,un�턉� =D���f��3��H-S��4���~�����4OQ+�힤4Dѳ��c�|��Z�-��7B�=z��*�����mt�t����Y�s��RX�_E/x5H���g	Ҍ��'盌���:�ζP��&h�d/�~�0iրȼy�%��{���(�Q��SP27h�q����~g\|T�W����`��+�(�3��x�q��N��s-?��h�8�8�I�9��lu��xc��j�l���Z���\mb$�)���1^�z�.�G%�D?-!}Ѿ�o*�1�~1P71p�\���f���K�� XD�u�=\�Gu�6]j�v{�r-U�(�����R;z
G6x2�� X�IL_EYذ>�hyl��X��R{���������������͢����-�eGC�@9cwb�3.��<Zѣ�������;��+����Gd�y�ʐ�?��/Ǫ�<[��x+�b������7+�1Я�����3�\0Ȕ���:?��$�0�ArG��&�,~-�0pɳ�&���_RP1�2j↭�6�}�M0���Uj~��a*�������Q8�����jw��b��	�~��Pq��g��6��{���[F��'{���Y��H�r�L�WT C*py�s��B�#�-ϝ�"!�o'�,/��^H�=M�K�q�#�F�$]_]í��&R�o����O�pµj��(G��dA9o3�����B���)W�=:~�d��S]����`�Ҫ��{ӄ��0�c.G�^8�c��~����R���� 2Du*�{�|�&����ߟ��ϛe��"����yu�	C���n Yfk.�]���v5^$&av]7�n�%�(��{�Nj�I�\�Qb8h�v�c���䎊HY��)��uH4<"�=deg```rR�����TEMg9}�_Xiڦ7<�MaQ+�\J� �z�Y\��Խ�BL�&*BBL71_a��>v'�֥ϝ9�,�`��E�e�hk'�H�c��((��m�V!��z��r�,_��Q���G����j�ܸ�I��\��u,?9��z{���(zg�����
�'���|	Sr�@��K��&�ձ
�7�}��I�7� �k:�v3;K�ѕ�.U����b������z��7��Y�⊯<X�l�FWS���ύ��od�Ŀ��;��'��n|�����[7d�<���I��P�ix�h���Oz<"����K����n��4�"�<�,V��*�{�񼾩䰴�Uaͽ����ƴ��0>�cK�!�#'Y�uX���	�l�� ƙ��Xj��
��<kC)��헷"#.T��$��,���H�^G*jf��V���N����@��v�o��l<���w[��s�t���zH����E@"������T�Oևo���qg�N��MQ���~��LNujw�]�J�'�AfH��J�-��\����4�]�Ө�f�Т8ӻ��V>odfT�I��e�x�Ѡ�6��Dx�g�D��nT,'��L���'%�`�4#G��f�>/r����3S�X^��[T^e�c���~�䲷�&���F��Jǧ9�Ь��)^�����Ml)*4�7Y��Ե�BM9]��lv-��[��#�M�;D>��{�uW�{�r�����}����&Ku&r�FJ�">US�W��9q�`g�R�����ey�ynyzKyyWMl��Q�(Q�1��d�ʻ�O����P;���,O�ʵK�{q���3~p����qy$������\��W�~ZJ�`D���68�v�nr�7�R�e��uU�h����~����G�Q@�0��Z�3O��r���tcS�84�xBc.?r�u���
k~��K\�R�J� �V�7g�P�<������`��9å3O��xk����K���prt���(�3x��2�ă�V��C�W���+�\������_17>{ʫҲ��vąr$�BM!M�U2t��cOdIY`iZ���<L�S��
8���d����B��	��ڊ�ֿ��*P$C��	�F@rjN������Ͷ���N��Ӟ���F����ic�?��,�-!n��=�[�ߜ����_[y��k*�EH�(;9+'��8FǦ�j����`FJ	��y���$��R1��J�5�!�Wc/�c]��4����)�Ѷ�=����?���ӆ�~r��+ll�2�̰��E��	�/��^���HE�	r(!�{J�$]���8��Bc((M���v�V�˯u��k��K��|�04+��}����~L*�"��ye���������oK/Տ�%`��W\�n�u����MY)�Hͪ�u�f�����)�1��x���E��UM�!��۬�y�H�fX��x_x٦5�Q�������d������=��t���-5�?�zҩ�t�&�S�\%û����ܾ��&N�#��p�"N���f8��t�O����8۳m�\}@����Ͼ u�6��P;�3cy4oq~=_���N򿞔,Å�{��G��o�Wk��it�
�b6��9fk��Բ�^��-炙o���;���=3?��l>WC݅u���OۧtQ���n��]{�eꈉ���E���sP�������w Gk��D9�RD�Z>B�!�ޗU�K��$_Na@1ap/iP�z9��/b΍
�CCn��L���/�|���b�E#ױ�~"�#����<+�� ��E�D��D�b���c���b�u.�����"��?U�%ϺSc5�$���G����M�v�n\�KT��x�_��j�;:��bP���!�� ���
W�)3տ��Mm�y@����'ծ`��\krw���4⡘���B.�`�G-�N�����&E���z���7�00�7&��_��c�����B�%e��h}�AX��a,Dw�SZ[���:��Y:)�Ԧ���1��]!	�F�#B�4�r�E�05W��������F5�#{�=|i��hp�G���������ϰ��M����� (�x&��)��F�In�|��Ϣ��^�7���-%�X�?���d����p|�*���AB�y�f�	���A���mA�oyZ�r�G�.�;�L�Z=�6��V��A�M�����U#���e��낑#�$�,�����=��! ٺ["��W>u_!���e�^X�lYK��V��3�*�$�=�����p;�/D�v�gzJMJӦJ���J�=�p&M�2���¦7-&gm��8;eVܕ��j�>c���ج!r�/b� ����W�ə�Tp��Eo`��<QL��}K��Ju�*.������9;<���4�α�p�c3F\���X�-]uB_�U�*���5���,�JwǗ[IZ�Қ��`��(�ՉŰ�$o�?B����m�O�F4w<�ow�_����j�5�Y��N��e���u�*�f�Vԉ���|#JT�5.C}�lS-��(j��Y:��";)+{��å&�[3v�L�8��C��̈́��ˎ�ϘdG�kA�W�\�I�r�B�R�M�Y�kp�x�H�vv�D�{3�Îh��1��p���cy��^�1���_����6B���)'n�=먎��:�?5�P�	4��	Q��jqa�b#�����z���U^��U���#v*dR�������#R���k����5�|����r���z/b�[��.���E�[J�;�]�����j�]�o6�7��~��~Vg�.M�L[��e��`����C�˫v�%M�8S0���4^����I��pe�j[�����zp��u]P�u#� Y_(�!?�le��N@��'�MH.�.�=���\ѱ-ά�B��E����Һڥ�m���b縉Ϭ�G!��7�1`�ݛL ��|53!�fU�*��5��.�n1�:�H?y�f����i�/ȠϜ��N�)ȑr�?��b���G�>'�����gṫCS�\�s}?�D��*�$ꄲùK��{5�}Yg�O�D��c�}��?Z_��m7�z��綞����vck�X�<��|R2�h҇J.�{�[^���B���`�#0�����Θ��c��T�|��n�$��eJ{��{=߲����4Q�+������`>��*�����;T�|������al	6D���>b㘘,?�f�����~s�3�x3��yn�(�~���F�y!�a;���"Z�t��=�2B�D�#��g~ʘ��m�F8�R�����Y,�`�!����H���_͡�k�@���=�5{�,	�7��Nam�<5�5ΩSh���D��h�M���t�0���� 'D'P~L���Q�����+B�*���J��K4�C̛��q���Oӎ�_&���
�`,cm�dL1<Yu>��3�����0�����b���)4Z1ݨ��c!����p���؆m�J�z�W�O>��������=�B]��2:I�q�8t�9�x��^�
�W97W 0����bV���&�RZ��@�m�~pm�<7s�G��\�D_�Qp�h�5m_��4��� ���8T��� �ϖ(��q!��'96l�B�a�,u�{i�!�-��|UWy�v�0���n9IF�
�["�^mQ�z�=߹UlAO�C.�,l�)핞`u�^Po��j��J�����?n�k3Lo��UU�k�T�:�s� �S*aR���Я���J��|r�	�l_�	��D	(
����V��"ABa�0�~����-�3���� �n��8��"���W��b��B�E��FZ�gS?�i���pWK�{��k]qi�"��z/�\��/rP~8`��{�դ!+]�Ք$�.�+�O�K��3�$f{�US��`5;��0�g������￰Y��V�Fi�]	&� ����8��J��u�[li7�V�+��>�V
C'\k��+�qZ�s|��|��jժ�u���7%o�q]���fM_��g�[L:�^�^=��]8&�
�p�VUюey<�hc慲7�49�I�X�
�!����y:�D�\��Yz��:sON�&^�2��O��S�	���7�q��B{\��k��
L3;)2��!�k��)���h�8B��ur��;�� �4�4�g�3�d�|�A-آ�ָ�MV�bʱ<�m4�sk��{5�DS��7�bw�b7K�Ϫ�ĸ�՘Ħ;����49%w�	o�>�a�'�]�러Z�R�k<�5)�*�(P�>�uil-/W��c(ʖ]�}���t�q\>���"��2���?�`�Y�k�����$° �4Ֆ�%��P#��y��eqS���Q.`�(�1X�9�k,�k���QO�YC_��I������b��Y�M��yKƣgs6���q����4�Ϩ�w��T�����y%xf�ã�uaL�z����c��!�Q
h�{�,���&ֱB����,z��e/��#@�\����0���	 ֔i%\� ͦ�!9���<�D>��Lc������7�(DJ.2��]a�!kB� ���o�u��+�8#�3�'���e��Vʝ�x�4zI�3M���]���$��<�	Z�{#L�$p-�̜����L��"�u������ �]ܯ?h��G��0�[��>���T���#92�V�3���_T]i#�-�6������eҠ�q�\qq��A���<)���Ա%o>��X�B�������A�u�#O[4LW��ʆ�\��������*�1p�hL`d��'��bMIop �p��ܹ�Cӫ��i��G��G]�ų��[́�2��A����9�y�
��=#\� a#������0���j�M�V���q���W�S��I	�:f����Cx��������7����AȊ����@�/fq������^$�⼨�2�� *e/Jy��o`+t�Z4%���dHZ7ɬp�v�qE���6���;1a%®y�A�u�޽o���V��PK�.~&�ِ�Ϻ�O��ڼߡo� H���t[���%Vނ���|��pŉm�d��{�-�ŜDo���EZʩ�u��i�$jע8c/]�6S�+���7%k
��Hj�~3,ˮmCױ5B���=��Me�!^XKom���Q�0���(SZk�`��_��N������9��SKAb2�+�2�4���P��Pk6S�!>[�4ZK1��0��2Ъ�
���Ŭ�-�A֋7��Ȫ��OYn�!�؄��g���s:Kt�X>	�`x�r�o&�2T�������kZ~Z�Z���zՌZݨ�ĳ#��rf���䵛8�?�D)����aM��f똉�n+T�8��4K1����p�=�i�T�'�a���"�v�M�����a�QɐY��T�Y�'�9��2}Adv�r��e��2}��1�%�#��&%F��8�F������iS1�g;Z'�ʪ�ѵԹA��=+��A���������w�D��î:wT[��,K��}��=1���Y� 9���_�滍JLK+��p�:`~���u[]ï�������g�M�c���*�H	��S-�aG�Jw�ڟlv�)�oޮw�Um�!�~��n�P{���5�>�G��0���V�k��{��7�,D���K��9t�cpT��bN���p�3���`	�0�H���Xh�S��������(�D�~�_�D�wc=B۸9�R�$���s�8�l���ڸ�pӿ������}����i`Ժ�%�_�繉 ,`��;[M��U|d��fgW͐�S�M7�a�Y���U{��i��q����B�)�D|-w�9��+��g��������aN]V�q�~�1��Ⱦ����o�	�B�Ƽ0�o_ȸ�G-��� �ٌ�:�opRB�%H�؅YK��P1�?��(��k{��nA'H�@p�,8wX\�����I��	!��������W5TQ=;ݧ�<�9���S)cWk[�\�؞E(��t��]�N�����T�I�}E�`�����_*6�QK�l���m��>H\��n[�FH��M77��ӫ]��x�S(�؉8��>�=�vu���5�0>7�d�Ϝtȱ�;��W��9�_�	�_l�#�_�믅d����27	��ɩx^�u��Ӂ[*�����2P��(	�t��~�;��%pe��v�y�?�\x�%��O�ԫ4OT�l��r=MB�ή�b�ǎ� �T���۝,n�Z��D���^nzlڸj��
�iN�����ݢ_f՟���_���m	��-l�y;��.[����MH�� ��L�kXG�.eȞ/	�e�qw�0�ǰ�_$5����:�\.��d���}��6�j�+�z�IA�y����Dcf��T��ˮӏ;���& ��q�$=�N�f{��7N���=r���o��q����U�e��TZq�]��?��� c�dZZa���r�U��kD}��}g�"/�ȳy��bsδ�F�ý=�7z/�fYN�����C�����/��Z1�v�#�BT߹2_�"J#��}��Y�e�%`ڠ��Dn�zd������:��@��8ޮ���@1�lҢY��7�F���'�w*`v��@��scO���E&ռ'��[|>�%ϛ^d�(D����})|��٨;�������Z���ķ:����|��s���_ӆ��a���<:�Zt��YRt�iS�Gɫ�����N�f��X�z���\E��,vkJ��rE�(�BL��o�e��y�g�p��5�R����/jc���3�`O_;��J�����x��CYKZ�ք
�~��M�>$��?��#�f9��ζ:�S��?#x�1]��R��t-Wn�n�<�h|�9R�mm�0�Y�Ȗ��K�=��v������l���4�u��,�}�lj׿~l��x����/L��ow7d���t5xj�
m���n-`gmAS6����}0]~�w1Z.հ���AgȢ�,�x�Zl̏��g��9*)�oլU"rg���掭9��H��\Pړ�z���>�h��`r���b�^���!�������_X�@`2;��䐏�B�R@��~�߃ּh�qF��,���r������H��F��a��?*�_���j� X�s�~�&F��,u+7��_�JF�ε�Н*9���@?'.[l�Y�A*#���[Զ#?b��3w}Ѳ�Qܼ�=����	p�>%j��޵ԆZ�Ϯ��O�o���I�.��� jQ����lan��^�V 1ϝ�q�d��^4:�k���-+,z5�����d�b�Y�yn���]0�hk�c^]�ǐ��WȵLԎ�b+[y����Lo�(ʗOojW4������KϞ����P�PI���8�c�O�y,�o�i^�l����
WR�|�i���z���v;��Ղ�⾭ƙ���)������u&�d�5j���Jl�z��F�f%�$׃����y~Tr�����������K"ϰ��xH�����ָ3�/���2�0d���Y���p�(�6/H+V.���M��O.ۥh�Xδ��YU��-�8��N�k�d�5�~�5Q�yv�%��V��_q�}��'m�@�;{q]`&��8K4�˴�1�\'�c�xG�oi�/��b�����?i�8�;�jB�U��_q���Ȝ��P��>\�v�~���1ܨ�E=A��!��w�����$`��[����zD�{s���l��L���#�/tSFT�ǯ�V1m��P�c`����E_�����1������Q����WTbNNz�?��+�����?�>ɟ'�M-�^���HY[1���I�J1���Z�Y� X?��c�p�=y%W���L]N��z*^Ē�m�ZF����j�77��i� 
�*�-+E�y���������~�}#z�KBXֹ-KkByy��4~�����63��=q���0�i�`EZ�ڞ�/<T�T��b5d-~I3�\����1kG����̦jVQB=�y:�n�uOL#7���ʭY<Brj|#�P��^>۞�3��o���Rpd)x�5�96Cs��$i���Kn���ӱ3�!�JAhouR�d�)�"v��X�~/��m�=�zH�����Vm�p���W����ָ������^�֏@0��V��t0�O�1�ԂĻ?ʡ�&�6:�\5�+R��.��ƹ�q��n��8x}ͯL��J)c��<�uV\����Ԥ��w�Q���<Zն�qLO�����+���R����>ğ���/�~ᮌ�!���A�/uL���~�:��1��\V[.}�?{k��RU��0{%���eXl/Ȋ�Т��%|s5M}���u�d���ە������vS+�S�2�?�^�3>"5�U��1=픗hQ%nPi�wU�dW���ӊv�"ū��7���]JdJvkd�,�ˏ���(3�% ����V\���"��*�Z^L����*�r	��C�����rC�V��{� C�����������|�	�����`}�>�i=Y����Ѥ�&e�x���=��X�˄J�4M^�q'��T���T!w��؏j��]z{��W�O��m=J�!x�Q<6UɄ���K�*9S(�=�L���p�ԙW-r�C��-zc�U�r�3B�x�R|!Z�w��3x`��We͇SV�����_�Y�Se��.d��7j��8��΂��w���Y�U��C�?�+��텛%�<奾�<ݙ�&{��?��:��a�8Ԛ����{��7�n�O S�
���՜�4FOTp���v��>rk�(?�'��J�a���:�Z�tB#�Yc�r�o�\F��-�tX4���"��v���e�22�|Q�9�Ѳf��A�o����wٍ��i,U������(w{W�2�\ɚm�vI�)5N|���"��VN#��PU�8>��a�t�ew���h:�!$7�0����~����6.-��P���Z�ah�n����MCĚ@c���%���^����\�g���u���9�Z��.�YS}������=�0z9��,ک$խ|MQ�i���13�������!=`�Ev���r��v����f��ygm�m��5E�����>�B4-9��v-��<��2I1,�J�2��	�u��_��Ki��m����7��O������򷘕W�Np�1����[$�u����Զ��]z�%�>��56s-��o����~�����&^��4n�P���5�P����}V���ܓl�������l�����k�߀�]<�}=��P-:���p���ʄ��VK��E��^H�(��S#E&�v�͠P�9[���H,��7��O���vɖ9�T�v�9� P=Q��������<��᠓?!&�M�?��e��HD�=4��a��z���´j�K��KE9H�~w9��C��f�j3��\���@O�%x���[?���RkILC��P;�)�9�n�*p�#��!{�H��!�?
�߫�����x�r����3�"���*a����������-��?�>������*H�8��t6��L{�7T7�l��q�"���_3>����2�f��:�O�A�1���&�Bx䪊w�-��(L�s��\wT79GZ�.N0���c��7yD�CS�X��K���5�����K��H^��o�������Y�PJpԨ�ԩ�+̲����R5���5�D,�i:��mƳ� S���ŢGo��������F���J<'���a	���;��o�^�4C����].P&������e+�GuӞC��uֿ��s$8�	=��5�w��ԩ��mKV`��)�i���\�2����fd��n�=��,հ�\���8m��?)�"j�9� �o��>�.<&53-#�#� ��y���m�5��T~u|�A�.ҿϏ2v����B����f�����ˀЃ�f�ο=��b)�B`�(���������i��ː���ڡ�:&9�����~�ϣ�M�sǼ�w�l�a|V·F�"����j������?��v�B@��w����;��sIv��T6�%x�����8�Q�mI�1.0L� m[��6�7߰ L����j&��osw�&Ӳ)3g&�p ����V�͈:7_��_�[��cZ�k���� ����2C '+�a$kM����*ьs����F��4��٩��~�RC���?N%�q�W/Yc��UaH他-(��nD�:Ҵ_��YR��h�຿U��r�A;ل�M}e��_�)�4�*gr襹fG���M�/��Ԙ��G�F6S[ �o*G
Ɂ	S����O�뮼�w�[���+�9��F�iC��.�^�bWp��S���ִ:��=�yXp�p�j;�/����p�)	?��N�i�C�\L�"�0C�#CT8���oo����0�cޘ����Vy����*`�J�Ť�ZC�ar��q~���1n��9���:����C��n_A
v�[��w[���G�
�bӼ�?��4c��c`F៿̺����ʏnlf���t���V!���=03���l��ӬW}k�<$ɲ�\�"���t�-s��������h��z��T���ϧuCI�~�����]z:g��|��n9]�`y���ᔻ��OJ�p���g�/�[޷�p:��NSO���-њҌ�`�f-�� �jϔ�q�Q��H���r���|�'a�+0��K1潠�m�'+�����K6ZzQ�@�W6
��6�v��l���§�҇�V�pT�(R�?��}��:Th�8�`��!���5q�IMIB�=��m��#+\}�h�fչ����G�xS�[�Í��V%??*�ݭ�˥��kQ��3llG:i�>iٕ��'S�RN�+��$;=�6��GQ_�N(����YT�H afTB��ǧ��5yiQ]k|��p���I@&���fm�	���� ��w�����ܑ5�;�;iԕ���%�#��d��/_d>��vhs|s%��P�(9�3���:J6�ߋ߭Y���()%�#!�����2G��z��_ȶ�˦^�EwZxK}�e��i�o�PLٙ���������XFO����/E��h��m hy�o)ݰ:�#���w�b��B�c�ՏҦ��
(�I���ؽO��R�׹�~� %<oO� �4A��ң'��%�TW�G�W�N���/�}�l�A��8S�j@O�CTL<�]��\�G�O+���W��v��b��~&�!Vz�s�7�[���/����U�|���	!�
��EC.gɢi�c6gv+�o
��5��	�F�[�)]��h��ty����Ȅ��-?5#�F��ۏ�&�����-�����Y�|������M�w'��X���D����"wd^7A�����U�^`�0y��'G��DL����Td����g�_:�ή
<��,�9�@%e|�5X�f�^�q��:_��:�ҍj�B쩅�o|�gQ(����f����J�]�ß�|�����c�md祸I�� �����-"��d�����J��Lg����m�ꛊ?�CR�p댱���9:FT���E�KFl�BT�i�hIl�P�	�x5!2Ƙ�w�7�Tq���w&(��u��MKFMK��d7U}�y��a�d�u��S�X����ʫ�,C����qȷ�td�5�ݶ��m%��2Fp��ź�#�o1��n�9c���#l�Yd(Eӕ=�%��WRfA����:�{@z�|�þ$%m_p-KT�0`�!|>8a9e$xyY���~��U�RIy�k���X��'�#�I�\y���#>�s\�< bH�H�C�g�^�iI����M5�a�Jr<��p��Og��%�Fp�z����I$���|i�V��v	!�X��ܸ�T�ił��cIA.^^�o##b�����w��Q�q��������GI�����~�|��!sp�
)7��l��0��^��j>a�7���]@��ӯ�թ�`�x��DA�J��<�����r��br�~�Pv,�#��,o;������Hͺ,?��)��	��/�������e5�a�ZQ�S�����9�k�3GY{L}�Ȥ���#�ﾄ�l�j����
KҶ��u��_l���0���_\�<%1.���j���A�a��f��}ݵ�%��>� 	�+p{��B�XY1����E|}��mi�D�H��V�% F����d3 �eK��_���|/��
�G�<�&2��s����*;=��+s��q��d�YXG�5ބ�f�A��%��d�����ji��`ةh�=��е��/�~yF������"���${�����W�I �rX�O|������H�۝�ՈA���@l=�'r����Af\�����������k�̹�̕�e���f��x��Ĉר8.���2_Kl7�`
��Μf��I��aS�48=�ݠ/^ 
�F����L�_�H�������}P^Ղ.���ҫG��
=`��aa��\ ��u,q�N��a�#ƪ��_�I�/#�ÿ�?@�H�Pl�C��-�Z������\��D�d$�����M���J�GF&� � �7T|�
Ӏ<����O�`�����>~��വ��B�>%$������R3k��ɻ�`�D�)��Tx"��O���~�lr�-B���o)9DA�u�5�y�K��y8C̪P!�����������$�p"zډ'�g��n���T�w��/s�J�&aw�R�SCLp�ŋ��yĦ%t��������b::$x(eee��������cj&a(G9��V^�&��AS��ZF�yPՠ~�p��O(�X@N6�t�UQ]�ȃ��~E�����rl_�Cf���!W,~>����N��� ��3 U��T������L��Ԕ��k1GGv���,�6W�K�I�nH�z,:7��)�ݓ;̥l���@ꅦ�s�{-켴ܾ-s%X�ڸ�sͧ.�L*�w>�Y�Ir� 4<<&:���p��>�?�$�[��
��p��&|����ٚ��5|���7��ܒ,�f���Ȇj�?ԣ}��BT,JT�*���w�7c �e�E���G��l�D�դo i��wV0�C=*H�I|�[SQ��o��������}SVWYu��cDL2ql@Re}}��;� _��2Ztz��` �y����I���a��+���z>�����<\�F�7|�í���|CV���g*�y�b�)�騉��շM��E)�mP^Y���� ��9�/���`��yy�\�c;��C+(��%��
�歟LW���@�����c��cS������6-�P|=I)i9@��v������o��ٱ��F�ӻ����:���\�rW�lu����!d���TT>��D���mk�ˌڨm ��@���*�����qQ��mL�o�Kr�E�F��5�_���Sc��H�{���Ar%8M]�;����>	�-;\<$��[W�l_����L ���y��$�8D__4&�����s��&>��T����F*�|�15:*���>F���B	�{ ν84�8��C'!�y
����_�8�,���0����DXT���\�


[�I���C��B��섒-Ҹ��Wl��kkqfgglg�#V�C.��d!\�,��:��eh��'i�;�d+�3�C*n������=ezГ��a(��-KԌ�f��!!�K0%C����[�ߘ��(X���*�۳��cVGI�A�>���� �I�KQʆ��46r�74P��!R�TV��w؄%l8d�ٵW�4�U�ܿF�q�_�&��țM��y���4ꥶ�A��z��=W��w��$L�}����6�Ѽ\��,�𸝨Q��ϡ15�
F��8��r��� aNnV�ޤ�K��Pc�E�־y���������s��[��?z���ۉ"�Ȼ˯3�2�3��y�*rr�β��h�t9����{�W�����W���:~�>���+ap��Z�;`AJ� ��X�n�GWL��C=g���<����$�@�U���wk[���7��S�`�tzsc��UH�nSx���](Y᮴���_�W���� |�Kp����d�j���Y/�������}�W����/���PO�\7~�HJ�AW�v�i0� � �)�f��a�E*+�d��z�j�]
��� Xb��3"�u�ߟ��w��][����E9.����Dp�3�L�(��z�|a��z�(�>FR?ɫRO>�R�l��j����'����2�A9����X��p0Fd�0oh�.�[�jaa��겯l`01�.n����TVb033� ��������<>S3&n���a��� �z�B��M"F~>�^�*�K��'���$|�i2�Vr�g�j��i�q�l+ZH��ݣx���n�M����źEo��#`����1`�w;S^=���B�����z@�=X95TS��4U
Q�����a�1[Y@d�h-*�R�!y��*������oM��p�&���i����F��Q�\{I3���X��ۃ��\a�Y�`u�rI�����>+
�� zm㚗�[��i���Hq���m^�n='amm�WJYQ����&؅��|9 ���	E��>eF?Z]�3)Cuas�M�T�H|����ib��Ylup�ū�����s㷜�Jm��ך�#=�_���M�:�ȵ���b�7�{�;��>\�|�E�j�e��C3[I��=�lA|zů�m����K**~2���a��?�����j9�ui�L㜑�H��)�0}�	�|�K���#T�,D��� K����F��\�d�����K�!�Sq<d;e�.{�^h$�85o+l��w"Eqϝ�c)k�מ^^��k,8�c�ύ�:}x�~"�RHB�}�m�8P'M��΁Q�iϸQ7��i`s6���G��b�g^���po���S��qt�/@�],�/
���P��i�����=9��5���N�Y�q�@�=�^R{�v�7%��I"R�T����'����,vh�G\���, �Ҟ�p\v�a�ݷ���XC�/3�
j��7>@�n��JK�}���繖LBr,]Rk�$1���]��y�A�El@&�j�IbU�UV��b!)�AM�W��|k�u]��@iE�@ܻ��,txqG�3���?�K�m'.&w��SA�M��8�^���Y�4�j�9�CQ�i�_Iİ��CK:oN-Y�l
�� :��H4S�h^�9{�Iد�PVXT�
�"�g�$?�x�R�j�*=��C��U ����}|�ى�'Y���p�tw��a!�`�Uq�D���^ϲw�r�l���W��򂼿�(O㒡2�aA��E����,|���I�����'1>��im�PT���Sm�h|�^DrD�iE�����˗�xJc
���f���G�&xђ��'F:M���Q�<N�Bq))Ľ��j�c���|jl�h,�'s
.��T�*�i��]d�(���s;�:`-8�ei.�&����%$C��f����)�D�Р��]�|��` R����A����fMKW��#e{���yg3�	&��!=��#a����y���Ϫsv��<MZ2
�̭��M�}>���'U�^'�JR�y�j*���'���5�E=�(]ء�T��\c��E]�b��T�&T�?X��r� ���X���A�Ҳ7�}87~�Q��K�/�l=zom�?[�/�ֱ�>`
^�a�Pl7�����qVa�w*�V�H���	����G'��)-v�C{���5�t�U�|dʓ%f��:#��L!��/\S�>d������,��]���V�ʠX�L~-��Y6����$��g����iD>VM�k�2����� �B��Q@,L�uצ[�(�0B��uKO��j׈�ǝ���i%m����b��eE�d�✊@pu5>�5��M�W�����GFݒ>�	U��8y�սϮ�iY��(�4�B�h�T�*F ��E�I`T|ҙ�����M��p�a��Q�
��Yi�J^o��N:x<Pu��7���Mp���S=^��%l|ۏ���H��y}S}}��bBA��ޞ�����Z�2�G 9;⊮��4'��YҀ���'�{	��<-CJb��,��UA������(h��t����"'ۢ��)�^��G�a4�=S��2Ȏ7S�a�p��xY�+��Ȕ�i@:4��C}��u�:��T>;�̥�v�"ie��Çʚ�ϻz��桎�'ihj�r���e�$z��8��E/�����������/�x����7K;2���
!��r�|li�⧝�9��n����s��!��;�ZL��E�;�׎Yd}E&���zfx�<<Z��) T���IA��O�	[�v㶄|Ȳ��6���kc��,,-{B�I�����P^azrn��]�f�r+�躹�@���=+$����঺�9�/0}��g��.�nL���i4�}'�WᠸԄ�{�V��G]ҙ9��7zr�6�����������`s'��.�`�u�z?���mPT��u(�k��?��j1^���~�t�E�?t���V���x��l8��gfg�2�FktGZ<�P:�m��#^��e��7~B֧�uaj�U���LP��D{of�v8�#�}T%,�����`�͟(Q�E:���&
,�{~�V�҂$���Mog;�5�>�-Pd�y��5S_�c¦��\��M�z@�=ဖ�v0]46��bL��`�#��Mhq��@؆�����<�s����I,�q F]�`h,�T�_~꽳�3��^c���6}�H1m�9�#k���侏I�|�UL��?X�h���Ϫ�\���(]�3�����t���j��g"b@܍�J�!,�\��Ւ�|�ۿ~��w봒�D�z'�r�0�ٹ��g����룇�I#W~)1���n4�GX{���E����g�ǹ��C=��@&O2����߯q�׸��"��De���x�).�FQ�
�mD_����|����T�$d���9!�'V���>��h�|s�=����]��6]B?����8��z�M�*�}Z��b��H�>ן��OD:1�-�|I�ap�s͹

�"���mZ�U3�ʘn(�Ǟ:���T�yE�ДN��,=�D���d?$�����1q���Kc jL�����a!���C�|����X�<J�7�;��F�!zJm�M�as+Fӎqԯ�\�I���T��+KمϾQۿ�8��y��d[�d=�c���gK�9�`ũ�L�a;���5\|�̥>����a�w��7amV���^��Rˍ�`�>�#�#�B+�L,�|��"}�/)ߒ0Fخ������g���Z,�N���j��[���~�
W�J'W��0FPs���g�OL�����'��=RS��bCOu�NR�R�V�R���_*�.�&�6B�WK��>��#E���P���	�%�k6>�OUIϐ7n�(>sHHQ ~��]�꿜=���G�9�Zc	��i��0x���x�9���ߍ�.C ���ɶ K|�-N�!��uh�U<����I����%��b A�6|�����c����O���}t-�]{8���M�IK�r���ݼ������ ��:�=����۶��u��1�|��f�O�B�12���v��a��k���!��b�2��ܱ��[���F	)#k�ʭ��~�Y��Ml��� ϵ����P
6�ȝ���ُ#D�*���j*pS�z̀���<����ؚH��F-::z�ّ���&� Aup�>�rZ�X���ǷDz�F4�(�ʮ�	�\Î��?�Z�e�m/����p��~n�U����K~]��.�s|�}�"�Sh=/,pۑ�D�3?V� ɉ�?�0)t�'�ZE�ƱkM��9������<�т��"����S�����M���Q�w3�H�匭Bޙ8���,NϊjHr�������$�Y��{�E��*؍���U����|�%
�󫝪!�6����1WC�1� ����F�E
@��TTC��M���:;� V�sx���FAv�� Dxt�����0D\�'WIIE�>�%!R��������I����\�=?ir�{-_6w�B"#���9)OK�^4����~w��N��| �00���O�C)�i��y��q��/��)0�"��@1p<H���?ގ�m��2�>v�����جI��k�#�T�����Q��|���1נ��[:�Jn���T�g~R�op7�.B�>=+	��Y6�1�òI��j#� uG%�\��������3tz��7�>u�����n�N՟�\;�*�^���"N4|�7o �j�L�6޴�/,��"����{�]�$B������2E�	��iA!�����"�%8pP6� ,���nѮ�W,���<}��_�>�����_;Y�����v�ݧ����tȆd����I��8�m����I�Mf����6�o��Kp��*;-��ةKӺ���?Uj��{�ȡ���m�j��Tf���z���ͳ6dtO������<j�y�5�s_�D:�Hxڵz��>�C��e��LS�����������I濖�\�\�Q �

�C�ǶNs���"o�UPw�L"��N-&]�p�z���V0ͪ�%����-���T;�)넧Æ@�^��Io
�	K��/OS?I��k)7��p�G&��l'1(]Q,)y�Ki೩`���q%��q�Z^v��J�moL���Vt�
~�o	R��`�E#��T�J�N��ޡ}1niɏ�Î�Ϥ5υ�&/�\o�A����X���Ֆ��}>��}�}�'�Kn�(9�Ȳ_ʂ��t*s>�/1�Q{}-�۟0�U�g��}u�j<]���ʿ6���#��j�@  �xr����d�7S��i��'��GPآ�~Ӛ�b_Ն�y�Y;�y�Q.,�A8@�����_��<�*� N�{���ҵ���A�&zZï'%�}m$��o_��>��t�/@�Xa_T�8Wv^ZZ*���U_�6�:��oJ�2���D*��O�@f����[�1���'�\Ͻ��gz���Xu��0f>������pzft���~��^\S�V{|q��;k�#�A=K�HX�K�^YsjND�Pq�.�{�C?�5ؘbT�,��QV�05����히�����9�߳�����1@�&��<��fD���c��F7�071���lg0����������67��J=$xXɡ\΋�����*��B��d��x"��x6X��n�F���\��:�V�%�>��3������q�S���z�״t� �f��F��;�x'}�4� B'���{�F'�K�~=�!!/���󷰰i��۳rٯFe\���c!tq�`��c�-ߋ��$x͛R0'S2eXZ�Y-�,���U��.�,�ɛ�ꌌ�Ԕ�6ĝ��w��L�h����Dht� S����}T�O��>�a5�����@�{E�	h�&��4�	���R����k������&��"7�Y__o��nak�����n���t[�������e�+��r�u����� U,Р#�%���aoxZ�+9D��(�vx�Gq0�܃�R�H^R�z��Y+�L
�]��#���>��3�KЁ��;�Ѳ������lmж�$�r��"��q�t�ܦ�y�����F8�LR� ���d�;\*��[D�-J����')GV�(3l�*�Kd���B�~�B�!���8�%�(��k務%<�&��#����V����W��Oޗ{���K�.bK�6�l|���/�{��^mU20KJ�G�B��2$��ω:��)\_ >/u� 
ll�܁�۔��k�,u�Ѷ���w��Q�Y{�*�����Ş�W�<��!�?���%�Q �i4�ۆ�?�m @K�ME�&˾�l5���$��(�N�A�[Dt�"6��!LU����a]U�Ǟ��QȩO[��d������	��Kxb�l�R��C����� ���<~���6�� ���^j:��[/�V}��3W'5h�@|l���Z񰥞�3+����w��Z��� r8?�b�h#�xݾ
� k�
t�e��x��H�0?I%��
�@)�1�������wI����E6���YCHR��hO���梗`ZjK�u�_����Q�MP��Y�傻q��:Ց���;l��v���$�{_ab�E���NUX~����S���Eh`��K�I�|�D��Gb�G'�B��ow:W�5��HLl���)D�ȣ��+Dۯ�9��Ah")�[
��"���$�B�ե��f߂�-dk�>�0%�2��I�$��<��ב�'�<HM�-��Wl��40������<�&�Kn0m� '���k�����w�[4!���Ee�� ��M��i��*����8��GE����_\��Q��ĶrP�ث�t�n�z���#l����@Lg�}L&d=D�gI�U��%N ��h(���𣭮4��A13�e�������l�n|W*Y��E��Y�
�RPu����N����)I����POnF�zf�GW�������n�
d����/Խ��#�8�mmm����q�3%a��>��ۚ�e�6ކ�q��U:m87��15���u{246�Tԏ�e*[�Q��"N
C;��p��ԗ��C��_9(�*ǙȀű���)n �88	�Aa��8d�� +�3��z�Z�"�A�x�����s#�����|���ݜ���s�wq@t.k'?�� �;y�'�|�Ӆ5�l$f�{Q��gg�jn����3�(X2���ʤB�;���,���h�Z\҉X;Ȏ,6�"��+G#���{����PG�W,Y���\.�I����vW&l�r(�=$���//C��]� F@�����G��*�]c��_��U�Ymf����N�#��j�s=�)��A���#=��yt�3������*�V��SqZ��S�VL-�'�WB��/��|zˬV�k�s\�KK�����b�u���7�!�V���I��kQ#�v��ϻ����	z'��jO����]�� 3������5ow[,���)��
G�#�����ɝ�}{���^'[Gn~��r���<������"PXi��I��v���m�� ��V�O�}�\�5v�F�'�[�k����p~��c�Ŋ�o�(l�t���������:�!o���;�m�	T>/ϑ���E�A��0��GV߳pcy�m*����F�YK{Rq�?���fcB�$Lk�0z���
���}Y�A��������M	D����Xǹ�j��������=���'��&����^8y�Ae	Daa�b�j'�[L�x�_BU�c_���-8�j�U�b�zbU�ry�{=a�i�1c���Z^ֳB�D���|��ª�//i�H�t���d��qK�(1��fY$��S�j��`6�֬j4xEB��.�)PFQF�cFjQNe>��4���OL%�ns3���{�����q矢��G2�F��>���}V�.�=�I�ɤȧN�n��/�S�Ӝ��{%�]�͊�: �
���^�Y���Y���U���"�%���Z�̗VB�+.�I��9to��z��D���<�����j���JB�6��_R��-�:��e�`�q7�t⛿�	O��܋�����q�Ū��us訆�V؈Џ,T�E��H��J�c�4
�m��k�0BO�o�����o�>�v%�<�Z��x���e�����������Unte�M��|�[2ll���"��OW�Cq���i�f+V�x&��V�?r�c�ıC�{;���9�_�i"�9�#���P�_Nj�S�Ǳ��Ce�7[f���6��_�[��]�<��]ߤ�؁���>�y�*ǅ��rTsa�g�<��'!uP���k�����~��N��������A�H��ӝ&9���.�KǛ�]o?����YY���~*���9�����4'>y�r�~���������\���c��7�Q*Ji��&<//9��r7y۞Q�&#�ʹ������.^�C�)d5��%�X�Nf%��q�B�ԝ�є*��٩����n/��a*������P��`���-\���H":��'û���Z�w}����������lkͮ����<�;�{�ʎ�;��[L�c>�%�B �t% O�o����!_���g�G����$W��0������|�!D�&d�� ��(GQy���tݼ��H�M�~j�M���T_�ӆ�MK2�1et�K�&���Lz�����Z�J�����������)��q��-H����&�t�j͙/�������3iT"��>�}�K���d�����.S#�Nx���d$2��	���UՒ��wI��HԼ��1���wS	�ac�܆[�����h��b�2������2��T�e篲V]Oe%G��1��>m��gįo�%�;Fapƛ��ᨯ�F���UE�
���6F[duW��x?�l}��splZG�:r�CwHo�}�zBS�]���l��(�6������]����EZ�o��7��G�������d�������B����>����k'�*�����x��]K�#IT�+���oc,U�����*	��Q��M�k�s��ڎS^;��CP�A��Cr��E���͔`z����d?�gy�^��R��-0��$�\	փIj(qx��6�Qݿvu���44v"�u�u�ǿ#��Jh���.��I�o�ފ�=Y�	���r�dD�|�^-�6{�Fs��"��╖��2�y�?�����o�mB�6�g���_W������c7v�e�B�,�u$*���JCٲƌ5B�m���ٲe�X�f0B5�%�>����y�3��s�9�{��y�$�<�3���(QF�c�흮�@����^	�z�h����AZ-iy�јB�}>8ã��b��k��Z��@�xhs�����9 "����W %?E���(���saqE����\ν�¡�1%z�\ǜ�h<НW��(��r�c�11�g}]�l�K�ro����-�q^[@������V�^3Mr�c-_�~����c9)�O��@Փ��IS�='8뷉������̘���p�oAy|�o���'��:�T�Ey��_�Ηt�fu�������?��`i�T+�6jq��'7/D���T*R.���X+���|_��Mg�ݢ`�(��W��!c
PcR���聠�F�Y[GҏWHXS�I��0�iɊw����{s�
>�����7��z[�F&Rm@Kx��c^U�H$���>3]����l��{N��W &j?�ӑN��ge�M�r%��Q��6/��?�hL�Nc���P.�Ng"�Kı���ݤ��F��L��tPtWAȝޔ��t}f��1t�ř��L���,��O�\!mS]Y�l��Q�U=�� K1V���x�e�Ж��Yh���]��:nD���U��1C�z�;�c�8����Y��_���Y�Ē���f֫��qy�ᣑ
a
2��R���p>{����ZJ�tݒ��taDu	�ֺX$�b���� ƭ����8j�;i'�oE��vri�u��9���%(�!c�|�6�)}�!��u�hQ�l����MDdI�����U����Oe���ǶZ�Y���Ӛtj��V�� %.��%̒�#�Zh�^�I�3ǔh˾st������N��Ȯ����V����K��XЅ^V9�s��1��U���U�M����Q�le9xi��:�D�ب�yWF^�9�1��`���:��A�":=ѓ�g� �~����1��|���_D��@�6��Q	c��Mp���ƠP�� n�x�%.���2{��V�f߳K�q��e˗1�y�a,n|�&�����8E����!�D�&M���h�� ����v"��v����e�&��.ۉ�V>�#�e���!d{����~��]��F���Z�R�H��{Kw����
���r���'S*d5�p���<NL�Fՠ�I=#%���,;�zˊ��re����!-��~ԋ��/��ỨbҺ������|�@4��Yۚ����2��e�c^��	���؝$�wN]F�`����kCm/�G���iS�|x�)�s6�'b���\OIi`1즀����_���+������fق?����x�n'���-4��F��j޺5��Wv^�8�C�ة��e��S�yrWs�VZ��	�����vԙ$��B�1��$*���!�x	���3������-t�1�tN�+1Q@�Y ���s�n���.�O(סo�|��b箋g���8v�MZCn*:}��I�j��N@[i�?<1��UY��p��qay�q��T�ۚ�k��/4�Y���8��6x�4����W���ɐouy�q��vOxL�դ���i�	"������F�����6�./>o���V��1Y��\�3S�_�N�"�==e�h����yZ�L�����Z�bɪl��@\3�d]���?HD�(.��l�+#�P0��Ԡ�ȳ�E�t��m�%q�w��J��L#����8�4b=�"9��S��H���-�F�Nevʺ�<�zr�УHz��Ѐ��2���0VW�3�����6�)_ɿ������b�2���9�;s�W�2��v؋������������jǶ〴�z��_�1?Rd�_-ٽ�f�$__6�oU��/O_��JCBqˀ���	 *�ek۹k�c���)[~!�� b����@;"L���{<T��?~v�f�oO-n���"���i�󏱭eZ�����l� zd@��$�xf�7���ʎod��կ8��������&�4󝰚�3�dPy{	�W��E��+���|�Z��;��p�!�;�[��ﾦ�p�*�|���j󝙺p�9�5ۥ�B�lmY��j7�Ƭ[A��*�Z˜�0��XliP��Sk�k9���H�CEA�v{�j���fs|`M#��8�H��_H9nZ;�J�N�p�Vzu���Mt�;�uϘ�u��o��8Z����V^�����(�5���L@�w��ӟ��}��T����q��qʝN��t�,�Q�<<��z0���!7����,|�9�gVJ;-2@C�P��Wʙ�>�_W��N�o�t!�q�D�0�i�ôg�0>��:�\�k���w�� uw	�h+i��r�Z>l��)KUB��IZ~�9x��A3ơ�n5���[�x�k���Y?:�)��~r��L�a��T@E�b�r�
��񹐤Wx1�,֋��11�r�~Y�)t7!R??��M0�b'������P���d������u�J��_�a�NWBr���m-�v���E�x��M�~Iގ���I}(ET#߳g� �j�۳�V��y�_�	J0v��qPI�Y�`�!Q,ݚ�h�~��5���,��9	�����䍅��y��Ȥ���\$�����f���::���;B�7��A�чF+�Bc�۔�iKm��ˀ�r?1�����DR��ww�w��ܹ��,vwkA��s1S�$�{4��݃���h!��9��KBݞ��y�H߲���n��l�U^�iV�Uy}���w��r��C�3�X�ݫ+־a=�jH�q�q��2
�2�=�4�p�SQZt�B����%��|c��F��o�!��_�V?Կ�9#dgN8�O��Wv�P�o��;M�����C�.:�U�o��4QE��r�����k�Dt�u-s�
(�;�X�������'��ZY�H*�𜨍�tPxXĝ&z���͞
o��[�tؒU��]s��� \q�\�m�7�|��Zed�i���6z�6��x%oS3,	�q%�vt�?�z�?����J�Z�|� ş]�E������ Me��q6�G	���t�y	��ޖ���+*7���q�U�Dl�t��]Z����'F����GI��Z��:�So��^pO����.�_�ߵ-��ՠ�Ի�m��Ф�f'��I���(֘XyOa�/x���eky���LfU���EdF��h4%���w˰r�j�y�]����I5	��u)07��ŭ)j��eB3����~�m�d����G�x�zu�=�� �]k�}	�>�P�fذ]'Ju���*yj�t��� {��P]���:����P8�9u��'a�E ��˅��y����9"#JCn�uZ�"`�)��yz��֥����G� f������0��1�˥�s�W��o������5N`�/A�du�/�;���v?���kv7���g,J�p������G	�x^��m^?:���{�Ч���юߘ�'��:x�� �ҢfZ��'剘S��/;�<+�ԓ�֫�0�!%%��
8�J���齏w��C)����ь�hk��N)d$C�p�$�4��:͎�)�Zpx���*2{S�D�W�ޯd��`�_;�!!%:����fe#�2r��rF�(�����츶�Εk@���{$Np��>�]n��;�xo��(�p^9��aPv����R�"V�� �{��]�J�6����tDx��F���N�8�K�gjJ���H�pC�d�cE@Lŗ]��c$SV�lI\��qd�b������A<�*����x1��>Y�Q�,e̥�پ��ۂ��}4o��ZY�](���(���3�e��\��cK8��gr���?��F����*lp=�)��n�oF�-�D�/��	c��e&�~.td������i#0� �E�"*[�2�'�'w�h��@}W�~
��~`l@������?���$�,V�Ǽl�P���zA
�h���O��x����/��/���/.�7�25*kS�u�<T�+.��ȓ(��g&��
3I��,+[�*�5Ū4_�yyI�y�B ,W�*V����B�zO��Ek�z[�?Y�ؿ�I<��!��#�?��ֺ�2��Ѥt����߁�u=��YDLO�4��P���� �h[Z�ve���޶��dIi	�d^���?�B{`붻�ӓNyYUS4o{'�m_���f~(��Hh����{���F(U6�?'�$`y����).��2 �P��9û��R�Gv@���9vV��\r_�}1�;#+r�X���/v�.�Q���R���\�dc�b?��./������.,�]q��7��t#���fF*�^)z�'�b�H�2��}"����v�?{\�����{���q$149���`5Hԭ���έ�L�UC_���a�P�9�p���ePlov�ÏwX�37�Y��a� M2j���N�A�H=���#��S<�����K?;ɕ���*�J�4A��jZ:����1��uH�5�>ǯ�����j���'�W��^Q�?r�I���j|����q�e-,S���r�s�M��}�+���0?gر!W��-�?��{�q��V��-Ӹ�ί�	�B����>{Y�m{k�'_��ꨔ��;�.P:�/f�/,��ʔpR�uMxRI^��6avu7�E��͊=���r̵��;�����ߘ����)n�z��q���g�Q�~�rV}��!o��493y.��!
����s��Tϔ�w���F����t"�n�MEs��}uEq\� �|�KIO9�	Τ�AzX�R��9����?@�L�g���g��b�g�[s�PK   ���Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   ���X�IM��  � /   images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngt�P�M�ED�~�t>��J��"(�= �	�C("�T���B%� ]�=U:�C�Pn�����Ν;���{��s����Gm͗tԬ�  �N�� �
	 ��s�*��!k��u�Wƞ ������r�}  n�ʋgz~ikxH,;1}�p�'���tn)E�EG;��ſm�3��ͦ�+m���0�΢��d�T�O�B���Țq�8n5���t����!1w��?�#��M��έ=��ݟm����gv�CLŻ�32֋J�։4���VV֋� ! l��!m��)_��.�[��]α�S >]O`�_~(BiJl#r��lI�.� �`֗�0W�a��?ư���+OϽ{Q�����1\��yQ�鉄Lc��l~�}�(	=>\8�(��z画~'w?pt&eHCwQ��xJ���'��XHP�F	sI[�ܛTN��n�e_>̎�8iHLv;��+f3�W���i�tU����\� ��L�o�"pUMI��Ol���@Y���;#o�s��Ōحj8���.aS����G�Yײ���6���)�*f�r��`��������_Z��#�a\x�;���������n<��㛪�k��k@a�����v��@��Dy�]d��PUrֻ�����bJ�/���>����k��c=��BV�V���?�N�=g���#�:�|.ƍR���P�t����B$��9EҾv<�4$�On����â�gP�ֈ��U��o줼�ْ֙���W��� Yr�
��U��2�߂DUͿyv��L "�H��+��P�J��.>Bm&���N���&��ff��c�a\V\}w��<��A�����|}",0��K*2�����k滠4��M��7V�E�A�b���W��CH)amR&R����B	���M���3[<(Y�z1]Ǜ���F�,����\R[���J6���2�&T��,��n�]��%`n�w�4fB\�}4G��7۔�+.g�����k��;�˳��!�W���mQ`5���ϟv�f��kTB!�̄�	��Z�QS�e�~�s��8�����e,�3���"�=�G�;����C���1�\��3���7�i@@M�M�	>w��k�or�X�K�0a��-/iB�Kt�	�%ai�J��W� 俗��W��;kTY�<����H�T�g�[��VS<Zeֈ֓*]|q�F
�����������obE�|W�"�wD�Ԙǒ�+�=5{�n$��Y��{7hl���ͺ�-z�N?��3��?�ܰN+H��`i<y(�y��^�R���"�±_?�w9�M+���g�2���Åg x�����ٙ΋v��������k����l�eD]r0�i����z�2���}�&���]�k��zw8[�~�DRa�K022*���M.��:����S|R|�]%��x��8۔UJ�&���(�W�����]���A������
�	���"ͧ_{���m��{�	b��\��999c�$K���vsf��@śN�nX��c	q����U� <�m��S���������FG��ة��iҌ#օ�q>������q���xT�0��SQ����Sc��YԔ����'��ƭ^�8>N��-�rF�_;�F�)?o@|�ڴ�h{S����w�(�.͠�T��񒕀ُ����_߈_�`��?#�#��z}�V/�/b��Z4�A�%�`��OĉU�Z#A]=���Qe(��A{�� {�nu@<����莮v"��2�Kr�x䱶������Ӝ8yoε��V9(L&W�k�M�r&�D�t�����TW�&�"M{w�\v� ������*��Qm<����2�g�i���wS�G N�[{:Ϻ>�yu%N��k���N��V����F]nI��^Ҹ���3ׯ��~R98�l2)���"�u������_%�����˞8�2@hkԒb%ĳ���_$_�yD�\���/(��K����]N��`��M��o_������X�#���k���G�.E�;�Vʠ 3+G���<;m/H�!{�P��I-+�Wפ%k*e�wih��-���	B��;خc�jD���}����?ybbշ��깠"K�u�J54����-��7hpѫ'�Z�ʘ1�ԑp˦�)�T�&+u�/�F�y��
������7����%H���ތ#sD���rC��\�\u&��'�|�����m�?����[����t��kN�f�9%&&z˝&�V�x4i��bT�^����^����>���:w����?��!/K��j8P���㿹?�&b��=u��	[�<=]��T�᳻(�.��n�YA�x9�{��a���,��Rā��/��|ҏ�˻�+�k;O/��|'U���</��h�J��o��Q�Z���B�f��b΍�A�NfF*�4�f����Ir"ݹF��F�.tX�R�>�1(M�J6�QE?^܏����<b>�]-��)���պ4�%9Y�ʤ��?�߾\�4��a[w%�UD��q�)+S�z�~k_9?�I<��a����G��Jᖻ&��q$���L݂�_ªx_f�BW��"��7���i���*��OX�K�,��M����f�3%�#-�:��3�������B�a��Z0�P%&e��8���Q���h�d(ۗ3��2���#�F��#�[:�El~���e�o���L�G����2���+Cp�zP,�>�^u��e����,�Ӽsݭ�X��.3?���Mx\�~������թy���5��]���F܈��U}-Is9;d���I���q��B n>���7:c)�P=�e��_�
�?v�B��K�<�w�����L�M{EN�� +FF%��=h��Ν�]�tN����<r�y���gha<�We������/�ؙ�^n�~&��t��m|,��pך0�[*�zeZ,Јj����ږ�0������`���G��Wx5x
�9�DO�}/�ǥ�S�2~��Sm�����F^��`dpc6���7�m���F��ݘ�j";�£�#��3�֩�oa{�.�|)fe?�I���7�m,�}��,z1�U�i�ľ�����!Kjo-'�j���)�{0�/W1Ex�ğ��}Z璱�^�F�|�����U�,`0�7:33#���E���f��x�T����nKU��т.��!X2ܻ����%�ť����?-� m<x���k��6dJ��!T(�.������u.##=�cXG��A"(W+�F[[ M�����;�����U��/��P�ØWI@"
��#�ݝ\5]���1���#�^65�XZr?u"�OOO	y�^3�W���yZ֚��6+���T��ZT.�Y��X����Xsã��o0�yD7�Ƶ�,��bXȠ�kx�tT̖�<�Qe����]�5��/�U��ܾIr`6JJV��P��s��Hu����k�$���[�
�s��$n�_��r��!^�$	�F"�#r]�V��Jl;���|�2j��zy���]ש��#1�b�!w�3�B��j����븫.%��d�S[��;�����u_��٩�t�'ߚ�4������;���2��^4߇��=Wk�A�Z��4��K�$�<;�&%W�eR��3���>+�@J���SL8 0�0Q�%������Z��L���V��o�9���>Cw[���OOT}E� �I|��p�u1���Z��}5�\�7��y��_0�3��l���Kf�TK�)�����3�����g��ݱ+�'OV�S�����.��QS4!,\����
\�������,��9gʡ�G�͋�?|~��ZT1?�x��=�`xnLKni�<>dbpz����B����{a�[����d�Cv��(��f�O�'�1�؛Ҿ���-ҿ��F�E�/��/��?hU;���QvBP���'=��|���X;���v��I49��J>��d��c<�ݖ0gRgv Cs9���m�E"�������R��Y��-�[�~�/AԒ;��A���~Z|��� 5�[��<HWT�����Dv!�Q]l�_2�?z�=�W�Mu>���4z2��b��元U����g�T�/�X��_��G�˚L���_�ƪf��=˖d]�o�\��?%\B6ʅ�E�@ �$vp0q�g'���?�N�L  ɸ�-��?,j�����P�o��k��QTj�\���'���\]XX��L5@�+�R���u8��/B긋����$G��͚�a�������ԟM=�:�G��Y6�{��.�~N�nd� h��?���҆3r�Ռ���y�LJ�b&}R'«S,����yH��duõD�ń`�l�����!���A��I��)���ߚ���q��@����	IdR����\�-o������y�]Ҟ�zE��Yb��*l���|G��*!=�A�8G��7}�y")`��<���Ɉ�,$�IB.@�
�z�>�:��u��a������w��ﻲMS`ك�l�\M��Kt>G�hŹӼ�"�x� ��ʵ�qbvd�rJ�����żu�hٺ-2�{����	&c�����_���c�cAT@��Q��|e��?y)���憽+������!������b���U���IaȚڑ�9+��E4-��Z\��z�]�E�(E�-i8�r�7�)�+|f���F��^�
\�Ԕ׏�yJ2{�C[���g��-6 ";���s27�;�Xs7xS��[�[�h��O��j���J>��R�'4���dzs��bAomqV�H���ǆm~�ǌX��ӓ)�ceBT+)uS{��ۤ�{	�}�ʱ[kr��f�i�x�cڂ"C(�`3��Iqx�y�%=
Zrh|�ED�����)��o�)���=}�Qr4�ҚSh�T��5�qu�^kF]�H�������6݃+�w͹&W[ME[-�q��s��`��X���܏3Ԋ �}Rn75�7�W#$�8�	;�z�%U�����JO��v��[A�g��]��	���4��l&|(-yɎΐ���'�ޟ�e��*�K�B}d���K(������������q��z6�X�Xv�!����b������İa@O�_`7,`|WϐT���t։�!
)�4V�d���£�>��ߜ��u؃u�	���
��*��X%_uz����KWT2�.�G���f�"��9��.1�COR��z"n���#�����ɕ&����f �Fۀ폠X~8������K��2Tp�y������c]h���n�ʬK5���5=�7����x����1E3�(
�b��]�3�B����B|�N�e�����VRώ{$��h6��!3�:��f���3d�C3�*V9�)���e�Хp���Q�g�>gux	��e'�Dc�An.�����o��~5���.G�a�����/�:�S3
\��	) 3l��]2j?j�H�ُ��XZ]�2xV}�:�=3�b@���	^!�W4�
�˞5#�5��u�����N�!��%^R�ׇ�¹P;@қ�����ۨ���1ͩ���ƾ���JSZJf*	VLI���a�Ѱ��q�J�)_��������C`�\���otú��ho(��#"��n�Jt��T^&��+7ƾ�n���$t����&ER/�>�HO�\�Eh0��淟UI(�I�=��c^[Ð��Dw�{[T!��bk�d�F'��Y`���_5�ҡ����H�"q&a��4�,[�0�a*0��2�htϓ8 �l��������z)¿���K�#辢6��ݚ���.ݜ�+����ևup?��*!�E�R�ˇ�W]��ee���M��{��5�,���3�s���3�[$��8��%�߱�g�5${\��'<��0'Bhel���1���W����L��Cږ�s�����~t�~"_28="W^�k�j×�o���ع$��s��%}�P��/+,�h4�Y�Y$&���� Fn����I]�n:���,-�x4]R�W�5����_�^R����fי}'o6	@D����R�m���y�<�dI?����Ax^Ĕ���i�D�N���|���Jޝ�~�?�/绉U�Vf3I�ݡ^���N!,�yWVo��͖u�N�/v#EA12O�Py-��Z�<�Wb�?ڷ�T�N~������kgD�a��{w�).�������9��E���f��7H��o�R�ݲzt�U��)�ƽ�J�"�������&h1�����O��l���i��Fo����
�{>���ť����X1Z�O��Y�цE����\yΓ�w̰��&.� ��G&�K��ث�@M���bB)]��E0����3f=좓x�,6!ˮu=_��dZgU�s��}���~D�`/ �O�u7J�&pV̊9
�zS�i1cnkf��WU�Y�wt��f=(!999���X먨(�)����i	�zj5�ͩ2�m�t�F�Q�Q�AS�;�斿�A���~���z/ַ�ʻ�1��)J�=vb������Qtp���gq���߾i]m��|��Le��)�TO��ݽ2V�'��~���퍛`��Ŏ�p
��6��3%�yZm��&��u5a^�3H�pZ�L1;*ڻ�Z�������gt�k����n����y˜3��W=���Q�d�^h�!x�����9XA8�$g��S
�adw��m�p�dw�Cy9t�dȥv�T|(i?�3zf�4��KtAW�_���F��B뽏p�G��X_��Ί�F���]������]-�&����\���ҋ��ME>U��Q�`bx.�#��._�$�Q?�ԨC�H�`��zi���za/�7?�ߨ���<2��)��>󊐡A�{��	./��Գ;"����s?A�܌��͌% �ïfntgʷ q��ϟyZz���N����L=��́A��R�e�!6x��ax	C�H������n���K��j
ds&��'�nb����NSa���[�B��䝶���B,�з߯���h���A�Q���d�Q���Z� �̊o�E�|��?��GD��e��Ų�scY���*e�i��ʑ�5�~=���)������Ň��^d��%L���S�^X�]�"�>������0�i*�R��X�h<mG�+5�����uՊA�B'���+̈��Z��$rt˒9Mf��i�ɕ$����]�i��4�H]&L �]R�c��w���d�&qI���2�@U0^�
�yA5�0aF�,��Cn-�w�#g�l
��Z��L�R8����;��T�>�"3�M޶2�����Y7���wwqI��Af���
���f�Enʹ�3`�J�͵�]G�8�HBs��a:��_��_����I*��uO�<��!a�-َ�A�FB����W�q���3:ۯΐ���v3����
�J<��� ��u4�c��	�Q?�,5d�PEHt<|�����*)��Mq���3��ҵa+%+��w��3�=�r�Q���N&!Y9��o�ƾ����5�e|��.��rf�]Yl̻�	k��o��gV�M�սg�Ş�&�(p�fXI��3��  �6!���[��,A�O���G���	��l-���Q��8�v�*iD��ҷ��]:�~��0h�$f���FqCPЬ���.�E�}��YH=D��7����+����|��'��UN��0��˘>B��g�!jyz�jk�{A���QkqĜ�����
�����T������88��ZpHE����1?�����@zU��-r쟛eu4&�\�jF$8�������b�ī��x�k.�Q�E9�y�-ε��<�	l�ϙ�Q�Y��KCƋ!A��7?��� �j�p��,,"޻Sgt�5u�w�LIT,P�P�u�T(��/��c:
�gqEj��֊�����Rr�9�D��|�r��FF{Fp��!MUE���
&)B���W�YG<��cx���q�wYX��2�;3��m\�QmY���b����+�y4dq��3�"�f�e^.�aAX`>
.���g�L�6p�Dh���m�q������^\o��� �s,�EW�=#��K�`(S�b$��2�Bv��VW��n,�����p��Q~����xg��ƴ�T��+��zۃ?Ͽ��(  j�/�r����h�&xC����\y��%��8X�f��+k�H�͇��-�ܘ8��?�R˝��xD�6Km��te>�|�m�T�Dr��?�|1��w3�4�;c���n،"ո���\���	�U��ĕ�>$r��^�&'�<��"֜2��N�G�|֐T������w3F����w����l2s/͇�M���}�'S�79�)�1oi4�i̔o�ۤ@�[�U6�Q�KI�$ܘC+���� w5!\^R�"m�$K�=��:`YY&�����Q�*[���J�8�͉O��T����>Χ,.�ppY6g�ӛͅ�R���B�	l����Br�8>�wR{���(��6���v<�x���H��"_��l � ���"�����֒�|��'p,b�P��D~b_�5��"�=m)��gh�ܪ�1���\^�(�X|f ��t�ʸu�ΊZ�d��a��=�9 }�M:�8��8,���:��8. A�Sg�u�Vuu�Z)�/��u�g�~BekLW��&$����.����kՙ�Ř�̦�H<@�E�S��9���b��l�����A�'�F$��Q�M@��M!X�rt��!}��x&֦���6����+V?�띣/�j{��Ѩ`SQ�g�B�<8(�n_C�d��oe�����Jy��b��3C���Օ�ޅ����mc���45�(p�S�r���κ��4��z��VB�>�����r�r��H�Ԃ.M��������Z$��p�3�H"���%nD�x}��sa�:T��ۻ,��<!��j���&�%��tvvu�z��Ĥa{/���G�-%hRi4�9�s������1�'	��k+J�,�ܩ���*�I�+�:��+i�� ���Ͽ�j�?���k�#�p��R��&s�>�.�l~�=#E��M�vk	��g�X���WL��|VzLE���`�ׄ�ce���#&����i�19od�dUԆG���Uڔ{�L ,��F����^����-��coY���+1�
|��6��A��'q����~��������Ay�֖�Q����҉7�=d��`���h}�wz����Je��>�M3��X_��!'\�c��x�N���E�Ɔ(����wJ�N��)��8�t��vH�Ը��U�}���[ٗ�T��h���	GM��(�	�1�X*Ze!����[[s�i�
�QV.9���?iʂ�� O*��[:|��=DE1���
�	���!��Ϣ>�ۣՂ�+�º��ӛ������v���B�n�u}�%�?`�Xֻq�����i�P	�c���ս<V�܎��ʠ��$x������Od=�S�K���q�Ay�3)89���u��U��?�yO_u	P���;���q�FxeF�N�Ȼ�lb���h����x��I�ܑӇ�KΝ�OW�cU����u6���T��5B/M�V\���e��}��M���i�	}�G;cL�%$0�1��V]X>\�A����o_KP/"�{�ퟎ�%�t�o�mG�9����(v�v/q=t�j[�ˠ�xJlQ��|��ٮ��k�d�9�~�����@��'�/�=�?'S���|gVfo{q���# �d(�H<=��~�V8��u��h�%���Tk��������'����ϑԫ��ň��v�:W�-�}��=~�A�;�aT�"��_��#P#~rdj
;4����FJ���Փ�t)�m�teZ3akl ���'�/�G��;H��}�Ѐ��H���(UF���K>���ŏ.Ԕsu����]1/ž��$[�����A�F�ݳ�����q6F̤����u<�Đ�3`�2_���P��h�3��
 lsõۢۯ���+�f3[1�����x��ČyL���?`�sx�,���$v�erg�l'�$ˈv����[��+D*�6�\�p�KA�c��򯜁�߶�=�S�1�P��w�( �r�K?1Ì�0�o�ū�D�ӟ��}}W�ژG����y������� u�jŻA8���jߙ�NJ���z]�'}����mj�c���颉����s�D&��͎����X/��.=��A]���׶ݳ��w���d�&�c��#�]ȶ�1��<M����o������1�-h&��ۻ�3$���f������2��7��η���pI�9��Zl�E\�����i��KAxp����%��Qw�qE���|*cfZY�k
n``�
^W���@��3�2����&#k����%�Ϩ(����B��KљK���"��B,.n���\娆����c���޹��m1��9ssJ|ͣGZ�������<��N��a���0�.��avz��^#�����ݘ��gdOt'?c��!�H��p��@!@���G��錄ڵb������ۉ��~�l�����Cc��b��
��ӯ쓛��	�v:BqYo�$_���لM���l��'91��u�=[�+���J����{F�(��愂�)�,�Z���/2�(�4�V�	]SX5�f�e����9��EJd�K�S����.���9�*�!�T�:ι}�DX���k�����=��屚!=F]Ї���v|����zv�K ��2D/��� (ة���-���8��yrM��A�r�J7Xʳ���LL*(���ڿ���v9��- �������;�)S?�����/��?�7���q��������"l�@1�� %]�3鷩Xxٙu;�x���>��)��%��l�[.��IQ�E'��������A\	ԗTR쎤 ���ۗ+����\��{����������YZ��5<Sڊ4s�=����^�'���Џ#98f���.|k"VЀ�ZCs��`7zy�"��d2����*��7���ͪR��C����V�I"\�kQ���˩�5L��"�����v^puw��c����&^7�]����.��"\8��o甪u� �������;[�\�cwoeO�{�?�$75aA���q�n4E8���7��u����^�_���Q�$&v�����^.�4�.w������	��B@���ڴf��+�Ϫ0]�9�@�P�
�l�̉�s�ʟ�����n������]���ȕK(�B����>�!�y�w��6!x�8B�{C�,�Z���j��/�W���W-',����"�:��ȼ]쁂*����G�=�{�*�2�?w��b\�3e��^z�#O�o�y���&q�+�%M����gq��W�"]�WW�2P�HF�)��(���1�f�U$X����6��e�Cc#��x��g�������D��*9�����ۼ��ɼlil(qRTrxi�H����<��_7��!�nV�rrT '�Z|#ь<���_�C���V4]���;��Q5�e?A\	��85+ҵ�l�dۊշVp�W���]���ف9����	aX��S�q�	�r���a@@ �#I�;X��ܗ�=Vͣw���r��*��ߑ� ����ܩ����o�ig�*��[�X�5���1�1�I!�Ͻ�*�nt���T��w�u�Kz��T!���G.dͩ�˛�&,T���E��{r.���5��`����1z�l��"wЧ����7g�Iߘ���GC$��̈́�ֵzK�sSG�s3۴�ӧ߯�M��Wn�� �oR2��N�{���&����i�1��L�o=���^i��=@�Z*⎮&P޴���lsK3w���^5uRW@�i�+�hs��|��$]�m���ɂ�>M�"�9�U�U��ֺF�;�p(�*y�!/"B��f���!^0`�m/|9:�W��8i��5�A/��P��l(�rOku)t?���4!�i�HϱiHC
Zc({�sb������F�+čGA�M��y.������}N"�$+��,����:�t����ְ��n��{p��$e@��0eq;���>�j*�F������P� ��A��
��(E�v�+��G���\�?��=n��2�<<4�B��O�N�o%��t�#O)�ޢ^F(������Dd8�=j��s��3����m�c^�6Ͽ�`3��&5]��㫆O��]lqU���M����g��c1@�_�/°�8�5�*�d����M ��0�O\@z�����O$�2�T�V�SΓYKHc䲬����3����=x��6ZN�9�=�ʘ������(�E�R�'�fOE̵�d����\-6Լ���%����6��휀�6�l�ؓ��α�s�GV��7������J}�㯐����Ϛ�=c���S�{:��$���`�|�Y�>v�=� ���ª���ιo�#��n��斫�SBLa��"u�����?N�<��!&C��O��z��dTI�B+��w��W2�jŁ!g-�^}ԫ�
F؛Q
��=���6�K.�0+�*g�;���'�<�f�>�K �7&��!:i�3�K$8G�����(s�I���+��)9h���򯆦��_ ~��&���p'��r��*�g8vn�KR�y6x�j�;�������U�M����.1�nƇ��y�����V뷮�0{x��9撒��rWc2�?m�1B���ۗ��ub�a,� 8���\X �I{\�k#zKU
`���Q�fX�?���o}�^�B���O�@i�sA���MA<���#�W:��=��f���"�mu|r�T䝄���c�{ބn\�*�zE4?����\n�r�5��^m�z������`7�4Dި{g�"���������4����vKy7�FC�N�>s�<ב�*[�H�ɣ�G޻xhXw8�5�naY��ԾŔl��g�fR��{�B*����p]8��vc0�c�I�s�8��%�fG�[⪤6��fi�TJ(?<o�1۷{S���c;S��Z�o��x��2wQd��t��ӏ̯nG�u���E8R3풤�=��ܸ���١�P�n���ц�`i��ԸyfϢà��CxO����ؕT�*�P�D�
NC	|f6ɷ�QR"�
M�`Wg����<����fv���h'}WmMW�Պ����*+�gɐS��B�F��z�}0���v�t����z�o���l��M9��^�����%���������E?����e�g�����6��Z|}�X����3zNQY��vS�a�S������sMGUģ����-������֭������VS똣Mi��A���z	YY6�oPh���Ij@݋���K�����{���{=� 곆	�������fr��;|>�����sm��Q���V����,.	k�ג�%�̩h@��PS?�R���/䀬p_�ؼ%�[�}CԱ�W�N]�)W�"���©��YB�!{��Z �^,:��*㻮W��G��E���LA��<�B��B�ϠUF�WN�NX�z��BUy��]���ƨ\(bբ��T�[�Н�	[��9���[e�cͳ���9=-�FȖ��,C��Iţ�:���qI�g�< ni�L�~�Y�w�y��ʘ�~}��K�R�柁����|�F�y�OU`�aA�fH�A[���	���b���Ծ=���(����m���K��K�g�q~fM���)\�r$
.a������$��ӹyɲ���+M�m=��P.R_U�[�a���v3�է�Fm���T����"x��7����W��&o*���G�zx�o�S�h뽜^8,Ƃ-b�8Y�0�a��H�\;e��lF対��iV�>&��Ÿ��;1���@�?i�+�9���>��#���7h�%-2�[8����SgSk��W���U�Ee��nd�5=B�X䲂Œ�!t�HR�Vab�EI	={X)�-�#<��V�xFC�ڤ=a�E?�X2H��;u��wY���tv����8��!g�˙��Us!���R�OG2U��m�T����u��j�VLƑNX����)/ܧ"��aI���%���^�_ʜRG�1�ʵ�t����=K�"U��h�B�oZ5�6:d���J &-��KF��H�X��ZLY/I%��稱"WA�Ī �G�FQ�I�@z�|�ƔX�üK����>
H!��#��˒�A5�0w� de�?X�:�2v�úueE5��`�R��O���_jFF�Ǐe8��Ԗ�u�b���A���#��z�4ޡZ7"uq��]�l2��#�G�9�W�6d��E�-=�K�TV>��/Ԋn�ܞ��"�#"S���t�����y1��g�k�f�&:��:�H�����h�B��R��w���cg��f|���7?2YQS�\��no7(6z� ��3..R��u�z9g�o�:��Z�<1�|���̱WaGo4�e�P��KN`ro�wC`ɨ��tW�#�J�
T�jC(��
�lH�:݃�uN���L��5GQ/��v���6��{mN�	��EG���;	�ŕ�P���֬TM��U����2Yp	�phiu���Vݩ�GS��Q	�td0"����_����I�xP?d����[��t'�6+E͔�U -��l��2	�ˡ��[�'�'S��了!�}w�/�w�t�����m_��"_����7� 3Y��� !���ʑ�r#P=�~�B�'p��P��/[�	�l��FNM���|)��Y�Uױ�灐�jtr��<@7t+S�Jl2��T�.�z#^}���wsL��O�Z'�8���s�`���<�x�շ羡�UD��V"_~�ʺ:~ӡ��6�I��.�T�'U���\b��b��X�5E��E��ӓ֖xw�jz۵l�0�Á����������,T��TT� m���+@�����E׌2��d��ISW��1>��KKރ*�^��6����h��+V�R�$�p�Q�1d�9�)��)� A)��냁VS���ဇ}��'}��K��^t�g�"t?�w��
�5���#�;��/����Y�@V����{��L�@�NR���u���������W������\�_����y�^��xt��"v�
 �]���/��}��ywl�>*���us��"��f^hi�2�n��5����~%���m��+����;��'.��2 ��^�b�`U�jC{���<��<�<�-�3�ⶵ;I[��u;���C�����Y��e))A2���Li��-<C��ky��b0�9�/Ä)k��vꞱ���'�C� ��YA	�o=��A+h��lK�@"ָaO�j�r�PBg+V�-���? [�w�N�g�� 2c��z�L"��8ӣz<֙B��P����g����#Z=ߩ�]]]�� ��H���K5�&��S�n�g���g���YQ�9ʣն��F��1��tnʰ���.��R��!�\u{��D�KK��-��IЀ5�B�L�������&ʣ2�T���)L2���x�@G��L�?Ϸ�﹐�qXI'tt*-�t��]����wq��*��n��2��d�+��1�%���� �������Â�󼵷@Z`��B���ު����H8�����7t���/eR����T���|�>*��!�W��$�x�@��M��&�4Ҕ痒�[�������g���A'���Ru���2@f�g����^�#dSðS�%W�am�<�
n������ m��b?��|�]�_���{��=���e�����I�V[;��W�8�D��&�e�[-���T�Css���y��G��>6���G�I�B]�]�������/�n��~��Y�¢�h�E�7y� �'Js>���}{U>xٓ-B[*�>�6Z
���D��L��`9�K8�8��&%�Kv���{H�2�l B=3>@.
�M��?ww���. }�I0Y���Ń������Xv~y��l��Ez�j� �9��1-_��ش���K�_��p洯nd�2�#&ί��k��S����ps/�`P��ϩ�E
�\u��3��4�<W����I��gڌ��JU���*!6U�r�K���;t�[T� �]�A%3d(���:���7�w�6{�	Ts�82ݟ�^��7"?�G������X�]p�U�P�<�
؃������2|䘶���k���A�������#Y���ӓ��'�h��ʶGX�g�hHi���d�T��q�(R�W��@W���w�}��?X@��s����bǎ4����vk�է(4	�3����>��/!��O)C�w?���^)�pv9�QT��X�Vg:����H�agqW�UC���)��$�=������R��IE�L��E'���8B��	�D��LjF����1���?-o��>�a�]���"-c� Q��&a7a�,9�H������E=���I� ���͹G�Qc=?���ߙ��O���E�=�Jb�29����h�-,3��<�6�N@!0�Wa�OJuo�5l�d%]��n4��C������|��w�B�8�@�29�mDN\;�������3'�H�*S	�		���d!�2��rk;'�F���!`�/-����^,ϟE@���
�"��[�7+���[%@:/��)L��0s�O�ݧ�,)�b��z�r� ����vi��A�f��Ɨ��ᶉ�\�p����� +Gӵ���9���J� g����X�i%T/��.ɘ���(�?�����f��n��������ao����OJ��B��.��%;yG%�1ٳ�c�k(%$�:$ی}��6D��}7�R��Xg��o�?���|�����������u���:�\#i*WlW�W�ΐ=�Kp��K��:�A+�k�2O�`��Ce�9�_wl�]L
̥^��on��q�f)��J���ԑ)@Od��c��}z�S�F=͑�X���r��s�@m /Ņ�2����ъa�1�F�(�$�V_*�SH������U�987T��A�7�ʋ �5ٽ��K�(*�3%!.��w�d�������ꆝv�����MO�Q�`��Bb�i�M#M����ktfۏke�b�	􄸷�3����=-���i��^u)������_���ǟ�����_��p�ݲ,1ЀM6B���嶱v���gG���^�,��<����`L�3�Y��%��ÎO^>|�K��'�s(�P�������HA,��qZ�-�|m��"�K�b}�\ �M�����	�V�����Ϗ@�A��~���Fn�y<����t���Dk��&bz�$	���!�X��Yi-FZ��R�a���J�
ms���noyt�At��L������,��V�߃������֖_��zv��-9t�g>�<�cr�x�t?R���J�,Ò7l��a �a�c��
�aN�3�0��
��_�j"�V��s�j���D�av�F�J�#;�����n�Rn��k��{���\�� ]��Tζ��W-�w����.}�(�u���6x�,��`�U���w��_�>�$���ΛtD�S����~�t�Y�G�uKԍC��<�uW��d�,]��\��Ϲl�b�������s^$���@�7+�:uMM��f^ߛi�7��1s�_�_�;�Uu�����gb��� /#qyS#ϴj���:����ZS������0���L��L^����Ҩi�YC�n��l�Z���\�nz��އ������,G�^�n�ؒW�0�lC���Ք�c�^��v0��$Ǖ�{6�^��o��F+���xǵ_���A���� ��_΄ e�=O1]�w[��y�QC�O�l�&�_0,)��`Zm�97cW	���o�4�����c�V��L;��_�7��͸{T���f1��?h��<��S���)�WeI!ۢ3+D�R�61�ѷ+����7�/�,����)���'�;�� ����̕P��z�����_s��mY)ȭj={7��Wߣ�N{�����a��'�4��OU�ú�6�L��QQ��3��`�z���`��"�-r����k:�8
F��c�.L�O^*X��u�f�8O�b�[fǓ�r�^Lb2|�ogLx��VIڀ%;��<�rN3�"P���m��O� �x�ZQ��);<OѦ��H�<���S��]�>W���fQ�r�`^�=��N���|Ԁx�ς%V\���cM����'�K�ݢ��f��,����S��t��B�>p�ǻm���~�S]-;&W���DgeЧd&yt^?��������"�g7	�W1��{���z�F$ai��H3����
c351���\�f�������H��þM������kM]�G��Mj�v�Kb�G��8�Zo̻�a���".�U2���yw�MF�Y��^�o�;3�����偛e���bJQAyY���&/M��?�s�؟-�k�S�j�}�r$M�����r�W�p����Q9��}�HM����=�z� LD��*�-��`o?����2����<-MV�{�������z���A�u���I6=yw�z���)�� F3O�(�&||�/)P&�����j���F���,��+�L��}���}�hP�yO� ���d�d�qDo��  ɾ�m�&7ӑI�%.�S�������8m�vN뗨%�./�VT;!��b:�ӻ-fM;c��ȑʜ�ͼ�Ѡ�]�b���pyA��,�����g������ii��L����Δ�p$�?�t8A!���fyw�Lz�����y��Ȼ��H�P��� ��s�J��¿�)�@��ğQ2�MݘZ¶ފ,s`�=g�5��"�� c�*�:��*I���"\A�--,T	����c�L�f>���*9;������Ҹ�y��,N�̷2�� B����)�,N���~S���4�����ʳc�v޶��,t��� N�������U����mjz����ޮ9��[����$�����c���އ�;�4��9���&b��gHf����o���N/�p�Ҿ��i͹�.n�������ԫ<�v������F����&nT�bl�����'G�kQ�϶XW NT
������ެ�'b���\L
�TƄ��X�~�<X�qr���v�����Q�Ą���F<��& *��/S�AMJ���0&٤�k,�T%����cW	�8�&����QU��m�<�85@!�������.�.���D�&<A���~4��I:��˶z�oA�)��>wo�	�r����({SeI͓�>v|U�*�ýa�O��]37w`;���i�������?o� �+@;�îo\��#���*{�}�����f���L�^Gz���-��I7�Q���=p�
#{r�~U��4Ihr��\���^�~�u��Ʌ��w���u~~_�Q�s(���}��M^R��-6?j�\8��8Kƭ@���>:�UeG{:6譙��(.����2Oo�9Ø� �_�`��s�z+g噑�����e��&yQ�c��M����� ��XO%�z��t�ɭ1�E����}S1U��Akd"�������U~7�?��R� _s���n*z�Dא]����si��Z�eZ�y�@�����������e*�/zȉu@;�<��Jh����>u;�ཷ���Ӕ�A��x��rי O��E8�S�z�5��ϱ�K��[��5����p���X�b�}غ���{��5V0�ݎ��sF����u~_��r�eN�h���F��vW�#�d�Ŏ�_>��B��� -���޳.��k�0.&�(q�5��oQα�/����A1�����.Tğ[O��Ĭj|�F?֝����^�?�_��ۖ�<�-���ƫ�%�;k�P%�0�V��9e��"��T�L�8ƴ�4�S�yz�8���!��9oȷS��Ci$�6��{F{��n?�Dy6�A�I�5���"�3��!9m�s$.g����"���-O�1S_��1  �ɼ�+8��|��ѿ��@5�nX̛�NS���p�A�j�7�n��&U��K[�IN��z����[7S��Ÿ��f
wxj���&�W���ɵ����=���~W��B��L`qW�1�u^��̸g*���;���L���N��e����!�~�������e�\%㎼���nv�|�+�_��܁�2KVje~rܮ�-��k���c�O���i0ip�?-~��i  <��97�S�n�����1�tJMƴ0A����؛��6��%�0H��C}�#��f�0M�r�?�n�ؙ�sě}���J�c�����+��b;1� �{?����� g�VF(�<�Xި�&���%�-?�.J�	3 ĸ��vh���z슌X�W�y[�ϪR���U� g�]|����fA��	�.�z6�e[�l=Sa��<���e���3����W�'��$�ׯľRs�D]j�>k#2Zk�T����}�� ���\��3~w��[F��Go��)V��[d1�oo2d��ĈptXr��I�� �$���.�^��{���`z��ڸ*�ePբ_��l�~�x	r�7���h�������� f@&f��i��(>�ĸ�&`�b��ը��lT�cN���yx3��h�A*ǹ�_����I�ݖ����	1�{��01f����t�V%�p���n���\痋���h��[�F<�ty��M7�x-@J/ܼ�{hbUr���o<,����Z2��H2%t
�CeK�7Qw��]��~��&�q­���>C�L��R�|�Y?��{���b�돋���٘�5��>V^/�͑��i�G��M��]���ظ�:�����WoԺ�m@��	�e\^����Kz�܉oɞ��{{K����c�P�9���\���ȉ5�����lb0��GE:j`��?i5+�^��9��wd0)K
��~�&'q>�o��y��F� �_n~�!���M���ה�f���>p&Q狗��P��Mj|T|�?߯n�'�?I;�n��s�f,�ٕິ�Dj�~;?;7�C��*8u>�E��D�����=�B�:O� ��u	Y��H����OuO<NI����҄c�e@;��Ϭdߢ�D�'vrk|nڬo�v��O��^��$!l06FR5�����"#Mȁ�� c?b���	�;�#E��x�=(aa㑤Pqqi�����ȼ,M[^���$҄zU�Q7�Հو38��1�=�4�x��	q:W��ieD�a���εU�/�{����W��N+ߖj-?�ҁ�ؿ6�"�;V����U?��dWvt�
L�1�I�)B�����8r�_�ȬA����mzg]]]/9��O���_���]��Pa��V�ƨ_v�O��ɗE�2�7m��7R�0#�؊���F3 �?*�g�����Z���-��ˬ��l����9�����!9�ӛ�g.����Ο���;a^���G)�'D�@)L"��?��0�=�.1c��G�vԕʾ�� ��Ƈۖ�b|~��6=R5�}��K�;��43:�M�ۏd�����s7Y. @t�Q�y��u��goe+
;5M�X�$әZ�0���B��V�z��-����;fR�<\��3�Y�`ͭHT�����Sr\5�t��+�<�KԸ4�>��I2-��z�9\l�H�tz����Ѿ#�Z�j��[A���1��j}[Jc�LT���į9��w<�/B"6���[������Q��m�6u���X�d
��������4�ٟ�L	��)�l�6S���y�ޑ����zɑi�NR���罏�+�Z~D�.zE�R7j��n��I�~s��g�EcU��a��K Q\{31*�1��&�Ɂe|�{�	��Z���j���^��@4 ��d���1T��0kwD�1�\G�h�v�*�,����O`�t_��9�T�d�8�X�]w e+Nai��p;���wE6iw��O��h�:F��p*lU���"�}?��X^]�s�~`�M��߆c|����:�UMV�`n�.>�y�~3��dB=�'����<���� g�-Q��'J��u��{�ؐ?�Cg=����v';׍�B�j�H���(�i�E��[#8?E���O�Z��9�Fc�t��y�Pa6�1T�_z�׏�/=:t�8�|?Q�57L��P��y�pR�3LN���T�E��B��ş�]FO-g�6#~Tܨ��tF\�t;GuC��h��"$=�5��6��SSO%�"-��t���N/K��Q*Pk�V,E��=xaÖ9"��t�vΒ]�G�n�c�c��]��X+O���P�i��34r�j�}[�M�Vp��2-Zz
�w�*�h`V<݃6rT>�y%���7鈁i�g��r��lM8��������)�r���8j���-��7��V����j��m�V`�G0���W��@���*��=|��ތ�x���j&a�IM��PnW��wQ�CꖊC-�\~���'���~*��1Z�j���&L��1�vS�� �v�~q��)/����nm� ]ǌ��p��4bW���n�m�#�?��d�'WURkdm���TS�
?E3�h�] �D%h���ܽu������
Ʉ'�OϽ5�$-��ob��~�`���Ǉ�aL�J������=��?ˋs��������uwyr(��J��C�l�)h:�k<�Q���P>FbK�^���ƩI���A���-R�Z�n�x-�s̎
���]�	"j��t�2�� q��N/ �|�����#y��mi~���>�	\��UvG6?�˛����9 ��1��v[������C�,�5�L��W��'A����+���hn��}�G/ʮ~�>��'���q�1_�YR��Fk��   V��mD�1�!Ş)�Ũs+\�z�YY(����Oп�a�{'`�Q ��m�7s�#�����T��:�̣]w�$I��>�کv̈I���p��T||Z��h{S���@���R�$�3W26p<�>��[
�x����q�a�t���.æA�T������^Ml�����|b��&����jTOKe�r1��o�
�^�vŎ_��߆&�,��"�n����)�`�~�y�<��"������ڒ���!���ꬹ�4���#��W����Q=���+Mn��$�O0�o�]}e�]2.'� ?ggg�n}C�8��W���X�Y�!����W5�L",����!�� |�٣�KN�T��ѩ��6����؉��N��+��G ��v**G32��f��׮����8Ώ����i���&~�^��;��vE�7��ZI�t�3a۴��HP�!f�σc�ʐ{�У��F�M���������t�u��[1H9�!�O�& �4�`��}���?����I)��Bp7�Yʢ���#�ת��؉V�t�Y���G��w�e�%׈��u��[���
}��k*~�0jķ���Zw��V �b,;�7s@���磿2�-��)@�����⚪֤ޏy�M��$ªg~b����\|8�K^vC�� 3�w
)I% -SԹ\D�Ŕx�O� ���P��Rn(�������h�sg	w��\�V�F:�QT�HB;��NNHo�}�Z&�M��[ �d�p�����N1����%��o���VBe�g��R�C��<\�y���D�(�Y��}|�+ֆ�Yݷ>_.�m�'k��vՌ*�+�.��t�{�nZ�G���?3x'}�U[���L�E��5H�Drr�2�����@���X�zy��6�<��ל4S94�I��9�=����#`sPض����@��K��)�ئQ'��	�§�N��6>��[���`}ѱ����^�V�����6����Q@���o��7��y�rk�
y�r�9`���,�=� �c�{}�3BJmp��;MPvIy"�I���Z%�7���"�L�[��6�]=<ț��R\s3�@m�����$��Ag�}�]��>��Hd�}�6���� ٟ�<}&����.�xYJ�_{k�!��Ӌ��31�׹k�g	���o����E�D 5��[0G�Θ��l�S�h;�\�VeƈL�K�����N��yP���{�,=0�gK����, QE��(��[=�����]��0���7x%�,FTT\=�@>>��\.H�)�Cp}=%' �����h�ľ����"[]��G���Z�}�,M[!J0�&"�5�4-g
�/���z
�˞B��� �I��ɕ"$NŁ�ʃ����\fnz^�v�嫙�oΫv���}�٩(�s�P2^�ٿ2����{��ջ���o��|8{٩#z�ŋ��������I�^���X�d$�+�h�F^+g/4��^pF���j|�����X!
U�?��-	��LZ<yM(��*��e`������Ķ�)`�:+�'-�V���mMLL��=<<neU�4���]$�d:9}^{Sl�DPZy3� o��/�+�~�	p�:��4�Y�]Su��r�ys���I8Y�i�fQ��\�`)r��C-X�=U��;�7|O���M��$ ���>hfO��2��E� ��U�/-3sT���_����V:fw9���ٝ(���x"�"�1�'��n� R����~��I�[~=(������cff���1P^ڻi�8��7FY�^g�(�m�F��dĈ��D���K�߁�qTd:�s�&x����u"ؼ'�U�����ws�x�t�'����A��0RtG���Ɛ%�������J�6�[t��t��>�
��D�~���H���i�g��gg�u��F�������A.�ZT��ӿ���(��
�e�>)k���V�n4L�W�{�hk]a���NA�겆���uh����%F_�0��:,���4ޛ��o�,�r.6	Lqz�y�ީ� �!Y��sUOe�s25=������P��-M�+�\N�����������n��}��?p����iC�d1�����d�t�	����B@�|��m#uuu���?N�窿ƻ�qƋ@��z����&0|E=� �l�������X����ͷ7X3~�U�M~W�\����yn�4׆��LI�!Z=��e�9
*<��E�P�z{�yF�ز�(���/A� 21�	���&���N�c�0���K��eML(����������y�*�%�����dT����1�B(�� �5}�p�-�e�A�`[�c寅����at��C�kjk=�&���UU��L����b8�g���@r�K�o�{��몯�>D�YH�'<(�q�=����^~M������U��E�/�g�<�h���ݙ�ܴ[
�BS�\V���\��s�IO��}�����^��ع����k<�o&JѴ�����U���U������~�qO5��-�`¡�B�(Y�g"�e���x�X�\�iz��Tp�>+@1�`�3���Y��Ƴ��j�h�Q�s[G �oJB��z���n�����yA>u���?ƌ���t/�l|���9`��z�JPI�w�x�󍪢>�K��)����Ѿs5�/L^:�~g���ݞC,t���5o�(�.�h���$$��� �����Ì�"��yT0�ٽjF)ȰK;��D��T�!* 7�q��R@��KG9/^,KII9Iv�r�6�<c��#�f-y�Y�W]% qб1C�\c�:}zls�����gf�;t|��z���^^^�,�tȌ�����h��@}ȃ��>�wۉq�����7��)����=�Y_��h����F��׶����yz���ـ���ɀ��B�dOUT�[yRH���v�Q�Ea���N{9؟���#6��e����6|�2 �S�z��T3j+t���塟m��Pq6S;:@�ΣU�GS�Ffn�
��-<2�LR��'��T��w��詩��Q�Z۫J�	��(�����������*M$n��cjϽ�G_�gh����Q�5;����bO�C�y�#�t�臡�+���^Jy�(����$��������_\{�v�$�����U/hb7�}�|x���2�������'1?���f����uDJͰϗ���fUˤ7�&峣=+��N�R��!c�{���xē1ğ�5���i��ѧ�nC��z�mgŇy�����5�v��tI����Ww$��_����)���t��?��^�0�T�9��kc�ӄ�l��|���g̦�� l�قA�>�����x�}`�s���������AJj��ȳ�v��n)daxz`��4MwW�r����$�n�[&@r��a��7��
���� ���9��&d��B)�M��ɾ�8�ώ	C�ZS)cc\7ve�ןg��q��7�.vv������򷗖��k��e�!E�Ω߹�s�j����g��kHEhP�aX�k�-��&w��?
>:�	�<�m컷�wJ�Q�ݨ��ny��kך�LM����nn�@&$p5?�͛U��(��@
<B����vy���\�nπh��ji��lE Qi0�0Dy�4��V��D��ρ�ٞO��0� V�pQ�~��h�����X��? �����/eo1�w��!�6^+��k
ս+6��N�d)�aMr��M
�X�޹�h�2=C�i;��Z��p z��vI2H�{��uO�\��!S�|���0�옃߯��w��H���8*�h�|�6~�X\���GE��aT}�Cu-Pͅ��JV�a��f�6���kb|F��Hʬ�>�iG,	ڤX�'=��Y5�&8�Pzm[2l�;ܶ�NF���2�a\s��~z�y�B�|.TV־���P�X���P��XAS7��>�n �vNx~�a��ݠ��y�X'<�02�A���A�p0������ey�)Q�|E�W^���ATޡ���has��n�r�TŐD�X�1Ec���k�j6�Vq����SCL�\=Yt���h�y��y5C'��X��g
���-m?2]�������Ct�6�SGyB�	q����O޷H�a����%� �W�A� �/\(��bA�Vh�eʃ���I�z��ax1i.��k�kۍ�nh��'J9�O�]0�?�q�ٴ�+)sy����*��ƹ��w�j"��ȉ�����1Nx	��/�)�
���jVr;jɋ���%KȂk(cB֠]������G w�q�����$�m�ݜ�����Ъ��Y�S_�!��Ň�G�{��P�NŜffA+��@�L�`��8zr���,�3�����O�����w2	�I[d��3E��)�D� |A��|�٨T�א��kp�>P)�3
U3���dg�m12�d�o�z�dG��k���ő��㟉W�C=>�IX �����M`�ǆE�R�
������,T��f,�ؙ
&׬�cFH���̶&��G5

�j���/� ������z��ޝ�ü�)��vv�P���Ȏn��`�����ߐ��+t黱B���eI�e�D���<��=[5z..9�L�A,��G�[���$x�:;�a���M�`R�:b-[��Lt��W�u4b��L�:�\vz���o�=9A����N���F������="az2hr��k|'��)�?����+�N��*����<r�pM'���;�`�$ҩ̤��a�^T�����bD��|�og���#�����ȡ���N>3|��3Qƽ��'?�l^�*�8�4�� ����9�\�c�8��*ٖ7x���d�����#Jv�M�ȿ�6PD�@%��v�?R~�C���^"d��|����]"���iK�ML<��E����c��A5�����G��vݟ�/2��B���^6��� �,������r��x\1b�M���cVυ�ռ�WM�P<��Q+�m�n=��v�t�� ���~�����|ƍ�����eL���cq7�#UH���~U�m,�㫍��!���M��Y�0	�r�X��7��,�ch��~�;�Hy��A���M��a�B�xWb���ұ�/Q��u^�޳&�I��h��`zG�o�m�7Kx����N3�F�W�����
�$~.)�~�+k�9����c-
��o����ڳ��� �`���2��l��Ğ��=��w]ZYҕ� �$R�{ Tō��;d�����i�]QN���^�L �1���
guqt� ��vm>,}�>�5C���w���9<�]3ܹ��6	��^��z#����kb}4����5\"�\>)���_��04�Y��]ܜZ����
��������-�T�h{���&�c���� 	��)��r.��,Ɍ_`X���p�6}��g1!�p8+�h~q~�Pn��G�e�R$������o�]�؀�U���G�\�z(��� ����L�S��%�s.3����~|�?:Ϭ����/6F�����57�	^q<~���yk�ZM%L��UǉB�v�@y����~c*&��a%�r)l���n�*�UbS&r���;bXc��c''�ba��P�}�W|�߂��a�̀�]���Z�kw�i=�,Pf����?�����=s�\��/���NK�@,yPa��^�I�3��5���r;C�Uכ����bX�Se���R�mv�j�ߛ�[��řSk������Ģ�R{�z��b�dO�]E����5�v>��:M�}.�qP{����0��Ă��Ǥ�% J����� <"
��}U?Y�\�b58��q���Q�C(U��3o�~wW�����慑=���~
��n��_-U�O�H�7sC�E��~șM�qD���	
eF2.��y�p�Jr��/�)���/�+�>�d�A�?QI�
%w��Xy)�:�o$���A��8�s�����6���v�ޞ�u9�:[:�n��̸��c��%
҇��3�M�F�~��8�����	�/R������k��H�bVxr�[[?�@7ϰ�zn,%��{��j�ڈ��j�"/�Tv�o�%����e~BSAu�n<|0V,&�RPd�d�K�=q�����l�l�ئ�|��
�LLh�>~N͞�2��cv�o`̶֙�JCo]��~������Gp����
� �+~�q�Ο�^��V��n�x<~��I��b�<�#;���5�6))�h㞼�aV�C̾X����f����C�ׯ_M!�/�K����y��pԐ�S0�?�Q	���/A@��J�	BN���{:�<5����*����+�K򍿹x�pag����o[5�
r|���rS��>/�q�������@�H���c�q<Z����'���ǯ���yo���R]E��>�<�\�p�6?z[���T��!%Ssk����5m������	�5I�zhn���Urr���9����J)u��a�z���iG��D>i��,����s�ߺI��`�x��/K�))��;��ID����D����m��|�4Y��={?��?r=洸�(�Z�!�V�аp���Z���i���nw�`�p�����O��(d�g�"jd5�;�_�84�08�a{ol�
%e�8��Uw�Ƥ�Y��;���7�6�m���O���͍LG-l%;Kuk}T�+��
��Ɨ:�.��N9����]�ƀJ���������D��-�:S�=��FF��K�w��`(b�^��Z�;��;2��fB�#��:D�i��p��nU]Zz��S 
���bbb�MU� �S�\ۛ��B�J��lXnk��^ y��,9&j���9 ���@U4H���u�|�p�<Wʣ���AW��=h+_-�bov�P���c!���7��������z�ˎ�L�ۘ5�^	j	�/�����k��c�f.��N�O8R��kΥt�I�֨ۑ�g�A��M?Ɲ.i�I�?�ň�A�a�.���t^�����%��t�az���B-h	�C����_U�Tu*)cv�v�Zḋ'�~wNu�ݖ���*�dk�-�7g��Ԡ� ��h�ۀ[⇗�R�r�5�(y�c�lk�������K�]vo$����n(�S�&qRSe꩝��:�ȡm�<G�2Lk�w�_���WUTTƟd�*�FM/���6���'7 ��G�\`7*���Qg��҂b��V�a�4�p� �=۱�J��QW��-�-�s�9����T=�Z�ݵ읝���M��*-��p����A��Uz[���Aנ��4$n���:�,呋Yٍ�Թf�oO��QČN��Ի��(|#8g�ylUVh����ƚV�T�!}t����n��]��Op�����gee��%������!����~��>���n-����%��0�������	�<�X1�z|	9��}���Cq	����lq�k�M��9���#ʮ�įCH"���.�>u�����`��EV���SH���p����m���2���&�ƫ��L�e�c)��]��+Q��2k�}����������.I�L������^�~FXXG7�,����k͈��p��h��i����l;��s���\���B^�&~�?�"����?|�"���+W�"b�¨���s
�j72d� .���g�F�/x�W�+�#d�٣����Q���ю�9���iJ��\8�o��	}�fjH�>��A6���J}p#p�>�y<z�5Z �if����a��DI���x��ʘ\�f�t��3ߥ������B���3�O�3����W|(���^ipG�t�T�|y,eK��=�PE�^h�]/$�&F2��@����s$�Ӄ-�\�/�W�-*�=$g,�f��
-Ɗ��P����D��T�sDZ�ax�C�L'�7����ʞ^y'�}`�돑�.�}�j��i?��
�8'����D��a��'k�|��tGVvy�E ם�ƶY �`L����I(�ь�P���Q �v�_�&�-�j&��רapb[���~��D~���}V��N�@w�0�z�8��Uhm�o@QW�l�Hm��q���?�F��#��'Qp��Z<(�p���z��^	We�w�.B�~��9�V�8�T�w_v�Xﻹ􌈕5�.���6g���~�P
��sK��F�-�>��ρ��~��t��֏/H��� o�Cw䴦�T{f}�@.3�m������h��Ғ^E��DV�o-cbJ�k<ږg@�x���`ƍ�}i���˪խ�6jЁ}�(��\a/,��p��鷛�����z�\g�z�y�o�Ӈ��~ !B��g���r$�qyˠ��M�@���xf I�����39���͍�/����	�R�@�� ������s�Bb%
�T��An�OV��u��J �Mx�|j,����AE�aU�,wuv��M0����5��6��A�]�8�h����Q�W��ey�f`�m1��GA(�o�=���N�(ڪ����i�< ����s�z�ss��1��x	���������5� �_���vc	�'cd"�E䋿�1���>$9k�H��U�����R|�*5hi��Z,���p���ަq"(�f����p)���i�����X3���a}�j�D��R�ӆ�Ө�\��Ɨn2�!6�2Z�/2�rh+����<֍�bs�
��5�}8���ӍB���9�����ڱ&�B;D��}
K~2{����i�y������hZW��1cT:t ���2�*�s]���g������O���'PJ��"*�k�v++������0�P#MMM}2�����x�L$�{�s�����5$J�q�%&LZ�08��yb��8-qw(����16��/�W��(���a_2y�'�RҌ����0���Ws6�r���5���ncz�O#+�KH1g�+z��H(���W"�7{ngJ���?(y�- 6�t0u7@��F^��{���P���o�Alw3Z�T�~��n���C�*	�4��4 ���[��u���j��=E�m�9e�T�aT>k��z��7�}�(9T(���&^v���z	��׭�~oz5!9�����*CG����>rV��1>0/�ի�E���D�P8"g����_��1�:}���ݻYOD9nף�!%В�-|�(h&�ٯ}�E�3퉭����������˷�����չa �{a�B�+L ���V����H<�o1@N�&6;%J��U�̃�����t�?�/���'ZKJ����7��M�8��s)���
3�Eu��f���Ń�2�	����8��@��)I"\����ڝ�s՘+k�ZC��Uƣx-���{7��D�-�H6F� ��]9�n/���ވP��ZbFI�����$�~�I�=Jx%8��S�>-�CLn�D�nd�^���Q;�L�X�v�W�5�3��w�oy���)��H4 �i�~�6�a>�
:Iz�AXv�.�qw`W�G/�)QW-X} Q6���oEC�����n�iff���J�~���|k��\8y���Y��L2�z���wD��V��D��/�> 2���y��tXW�q[g��i��E�bJ������P,��[Rmʴ��A�a#�i�CQQ��rI/x���p����ST��}1 𧨧��Cܗ��.����{���ԏ�}}��>��a�?!P���{;4����p�F]L���w%w-h���{��`?"##p��ǟ�$�6�d�d-�$�ppH�\���yH����X�~-L�|�94��DsOO�:T޲	$@Rԋ��믨K��=�#� �L��S7I�_E�5����#)�������1���%6����
iy�B��Aȹ!)+{i�QSi�{-� �[)g���x~5y����H2�M�=�%F�F�.�ǜH����P3+�_���EH�$�-�鲩�B���f�P��HG�xwk?>74v(�RgA�q��C�@s��\��%_�ӿ��\o8b����������#��HEi�c.��;W��R�;wg�w���<��(���-.a����+Z�X'�ď�w������Q�e`>o��VG���@�d�o�7�2��к�?)ciFQM~J��yQ�� _�=ӌ�H�4�%��N�u����V�J(�3洷yth��p�;�s�-��FY��{��}��)�W�E:���\�]���jx*[�� N�����u��ԟ�@�n&��}ȝ޹������&yH��z�Z�����)�M���e}��|���q�e	1�X�+��Mb��^�<�8_%
��K�����
�uL�7l�p$�� <RrG�䫆�nUS�Mm���6�!c�c�mk�o% ;�y���O��-	�o�:e)�������7�����(�Lh�/����'}�0�h#�̇��*.%�-_b��-1,>���[L|ì��>e����Iס�E�F�[�3z�+㮹څ�v���p5RR7M yN�c+��H逅X\%��c/	��h7�a��wU]�#��F0��^LެA�����t�|�/�տ����ᄌ2�šf��Sм[K�h��r�dA����^1@�J�F �4tˈ8�ძ)�n����v�"��tr�4\�6i����B��K���œj`��g����v�!�ߴu�E��j8���l���C��K�=�PU�����c@	��3���+C^+!�<�}��ٜ�D���%�7�ON�hLكg�T*�;�MOMI�%!+���?.��Q��J ���R�Bw�(Y�Ĺ?�-�r�<��k�#��o��f�ع0cȾ �S�K��³�y����6�̑P��5���z���KX�	�zH����;�+&��,�_\z��.�R~�l���,�_yH�|�����4Ld�	�X�J� �jM�����X2�dx���`7=r�<p{k��;b�&�H�G�G.�/�\���k����ƛ�$IӴ<s��Tyc-=��/\��~��g�ʌl��K�Ӧ����(�5oB�^cL5�r���ǀ����+����Yz&�����#��|��a��@��?fuYE[���J��ؑ�ګ�L�5K[{ob��EK�BlboB"�����|�����"ו����\�q��.�Z-�W���LQ�[�,��>~r^̣����Xw�Dj�g�\�6B�����
9`֚D���K���ۡh?{���gx���r��,͋[��|q�z���"��s�2L�?�}�n],>��)�>�&鱐��7�z�a��r����"�uRꗠ6�����
�4G!p�5{�CD�m���,��ӵ�:��(>�X������GZ?	�iP�C-Q���犆^5�O�i�'�ɽ�PmS`�?�&�h�ٷ�ӱ�cx���F5!9-Ox�[#�ޓ�2�k��i��9 ���\���f�^i�F��0=.�~�l? ab�k$ �'3`��S텼�2����.�c���g��W8�}N�.�"1&I��h0LU%?�VK�^Ɯv�h��<�Y�2��]ﰣ&(��E	6��i�4<�G6���z|���0�b��B�f�6n3��`��|��KU8ը�	c���H�gF�^��1.���5|�%a�����E�N��=K}�a��VD}���Z�)D^ P51X]n�P4i������AȄx@�=�eqi��k4®f�"�P�C)��ΏE��$�%
L�U�}�z�Af����{��:��amQ"�=�VS�Ov��{\ױH2
��R�0�K$hM�	L���.P���{��p���C�ɘ��f%޻�c�{cC����C7�)7���C��<������;_�X���b&Kۏ���MSҠ��F&
�捥B����rk�|mt��^��>��x�?O�0x~�=��!�_j8�*X�f(#mA�����c��=.q��Yv+_f�e�����=��Z˾�u6_�&���3 ��M]'��N@�K��.E�[	�&�$Eu�2�2���R�J-7l�7��a��r̅3��\���N�y��w�y��o5�hn�S\�<�$����Ѽ�s�/�I�]T4�����|HM�ݤ��R._�2\\-�<䛐_�/䗃�{#��v��E}�j��ߐ�|��.�C��f9Jq}&LF��C�; #@���<۟������uO�}Yc�µ��rH��w�����To�o�@�(�`�#�lΕx��a����d{w�M?k�4�>Z벪�����0��rXn�?��Ee<*�k�u&臅䓫�T����7�Z������k���O�����Qɱ�n#*9[)V���3A$�]g�/���Yc�����G�3QA�G�#@F#���=�N8%_��1�k�/٪6���#��IH�y��'B�X&`h��K���m�m6!����5�O��|�w� it$��|��o�����A���:ﳗ��.�s`]��̷���hE�\;b��P=��1(z˞���-FO6�?�"�{c��������D*���.]646fL�-�x�M�ˇ;v��~��uz�ZA���8
��6��cE�kD�p
vV�q��H�$�!�'z�R�?6jRω)�,��1K�z�1�z��}�7��lֆ8�A��N&|*�m(w��X"ͣ�/Tlؕ5)��u����I�ƨ`ǵ!lȤk�Ž`�c�vU���o'�q���j�8V[��4�|�5)�zۣR E�ċe�~]�7�8NcB�iw_^��l��p�֧��Y�żv�pB�vuN('4�����90�H��]8l�;�
A#�o�{��A��4�js~��nq���K�"������Q�J2��}�!.GTF~7 �L�P槻Y��go?",q�`k3L�g7b��� �D�q_�x�V%:�oD�6��:�B3 kI����Q �K��B_Rڦl�;V�O�ةB����=�h_.�3�=$������n���Y/�ދ�,sW��E�3�6(��RP�ʟ��Q;�@��$���K|���X(C�����7v�|����C o�m��S���[�zWl�����CUEn�l�i�F�_�'wk��;�)~jjE���]��}UpU��vN�>�w�����H����(Xn5f^�[ԩC�-�z���h�:ܡnU��8/��{b�vs��T�ҭ�9(HJ����$xGѡ`�@1��<��-�&O�B�F��������q�����y�(+�vK��+D��J��U<Y��DBN?�&v��55���/F���!c���� ��Ec�M�iDS����<Qrh�Z��a������GO]W�~]�S��m|���,�^P�o�U�G�g�Ʌ���<?�������5��n� f)�7Q��1C<Q�f�0��t��-�^�6�ނ'k6GSfk��gz-o�5[D��U̲b|Ф4r)�3���{�R	�/��ܸ��w��r�B`��;=�p(�6�	�ޣcTLY�ku�2Z�_�<��=��h�׵~���ha��de�5d�B\\1��GI`vεeQ�󏩨o��x��!poI��1@��]b��^3��8a��4x��Z�����L-�ue����EU�������6i*rtndq���q�`w{?���̇l#�>��bAQ�7r|�vԟ�����8t�����i *���up�W�^�w/~�hp;�s�����E��D�<�Wl�w�����;\>��i�.qE�Ĝz�K���)����O&�Ӥ�:�|-2���e[�ޠ9�2�1�g�����"a�ޠ�2u%�Ύ�!�r���sj��0��^^��@<�R���|Z�y
��������\��s��R:�|��Ռj�Cd��l��d\,%j�u�x
_�$=�s[�Y�g�2W%���M�"���]zl��Ps35«*s/Y-��j'bTYF;�����:��7����j��@��K�:��A#y�;��B[B�W�;7'�5L>`��Am[�q�7�'�w���f�7��gAF��jw0�0S���E����P���4Za5|�g��2��Xw��o��� V�����-w.M����8?���g�b���}b��O1�Ǐ�N��K���K���}��~�s5ϫ)��UI�Q]���u ��1����n��[�6�.ܚ\~�j�Z�8�*r�<��g� B�>��A�.7�!>KÏN�$
��G������}��H-DV�G�J�4=�S�nY{�>���ﳧ����'M�a􆰷�^C�d_��%�W ��\�b�O���Xl�d�ޘ{���. ���d�c�Q#)^a�ibd�������7ɽi?Ԧ�C�@����9�@�h�x�O�s��J\��K_�ƍa�C���/zi���z����c�ө����WVW+>|���ie����mG����-
)ge�vH��H�2&&d��5�S���*#�ER���1T�e���h���+�Q�� #	甝WE�=���G&<����_u�I�{�t0Oo����!#�6ZcD����վ�����Q�^1��E}�W�1����:U�e
h�c�º�Ӎ��ueu���wZ᭦�S����$���3O��Y-��T9S?�[îak� ێV��Dv��e6Wʭ��;����k�˒B�3��6����$.wݽ#Qu��S4���$75��r�{����U�:_+&E��(����f~̸ۀ�ww���Z�΢�VW�����n��;����yyN�ڷ������`5%Y��W&���%�fj{�eA�O�ʇؚXtZ�-�Y4�d�WkV��8x���Z�Jm�mS����y���@U�٠�Kw�O���/qEJ�a4Z@�hs�l��h �<�yJ����K"��Bw�)��I�֖�f�ۊ��z���Q��$&��-��L�r�S{j���ZR��X9q��n"&�qGKP�������#���r<�H���,�j$��ׅ(j��.�U�8k�E MN$H���߅`n��ma�-ʼ熔F�3k.��wx���\de�)ڝ�ȎXf���/�L��$sz��S�pV�k�¬�qc���N�:b�l�����<���ݘ?�(h�u��s�`��������{FWI� ����+c��zHL���XG��F��<C�R�ȵ3h[Iϋ�_,l<e�4�_�9������-Q:���a||��K$5	��ۂ8u�z�B��xX����鷽�Mt�6���]�=�P�ﳞ��V���`���\��5�}QD��P�����IĞ��f�/���jM���q�i�k�F�����F����G�~�	F`wR�Uy��`�ȔLNZ���'�(�mi���7���y��G�p�����܋Q5¹�!����7�����*�pܿG���8�|8�(#pS*�[�l&��*^"�_� uBh>�R��o�\�w�7�j��+ĝ�Z� �t�g6z&��$�n�q�S�/B�������/�����!=��H��n'+~[g��"LY=���x�D�7��d#܈3l ]j1��R�4jM@0�k��ʍ���d+c(��ﭼ?="����O�:E?T�:���[9�Uv3�;AbE5�����_=R��C��]ЁUש��?K��^T* �WI*�S������__M���5<Yf�N�ŗ	잗4E3՚j���?�{��G�N�q�Τ%��Ɲ��:[	��wo]E�~tQ�������U�/������7�`#1'譜��t����X�՝��8$\d�G[�RK��y��~A��Ҩ�	�M,�4~ �ڰ1��tm,+8d���M�>#.��J��}<���b8���϶��cZ���d�J��jj�c��{�}�1U��A�*�ΝrI������`�n�����i�]Q���p�7���(�Rr���<� O��z<kj���og�?s��`�]_q�V�qqIH̎�5�����J�Nw�h�y�����t
���e�Ct�K���m�����cq)Ѭ��:Y��4���:>��@Vs�#�$�� ��@��obn�ܰ�7<Z�-�b	�au.y��9�`~��NȨ7��I��(��4�k+���r�wP?�����Mz�>����9T�yW����͌��3|�ڨ�b���������C�f�j���s�O�An��(na�P31���6?�M>8�ǵ��������hC��N�`&��t�d�`����|���&A�C*���5�7�k1�<�g<���65�������7�k��[�M����K���ui�ƻ�o��:'xh ҉����H\��絺���2�Q�*�8�U3E��A'�v��ߡ�6��6B�-I���)��9��8�X��q8�������t�;k����l|��7�ohn|y��������R�
�5!OTnm�<E7�c��:�E	�㯜µ��5^�b�U"��7 T�Z(F&�x�Ȋi��ebI>8
�/y���vA��*�	�O��¶�K��0��,�
Ė��M738�6  �`�=�b�[�����9/N� a��Rg^lA?Xt3/sʪ�c��ݿ�e"q5FF?����6:�'3'����:��z-�vf��t�q3��g\ e�w$5�k�8ڮ'��q뱇����Z+��i&l�8���O�$f���|���zl++ѽh~p8��� ���>YΔ����VW���9l�O��4/��
�}NLӤ�Ηn��#s��|d��ƍT��3/�� ���G�X%{�C&��lc�~��y����C]�py|�۴G�6�.ɒ�V+{n���NA�E�
� �`���|�^~8{Z�R��������0��3��R
�A�6���pW-E�'��\�b�~0Ԇ�8�n���Z>Z}4^��p5t����$�q��
�M����U0��J-�aJU�i�9�U��`����p�
�I�������}�v#p[�=z,��iק8����oB�����z߀?�B���ʟ&l���A<.�!�0��w*2t�(=��fj08��y�n4�EAe������$�O��捼�򝨉vb�4���*f�8��!J^��p#��)��'����" x���pe�Ğ��6��O���7�<(��rRTB{��;�a�Ǎw��$�~�X��oa��O냠��O�y���&���ĺ+���ib�E����,y뒧P�����f�e�j;�K5�Z鬴�d���deօg���{�^�Y�T�%�ѻ&����x�*���u�}��n��oSG�
�^'��=&Zs;�Oc8Ӹ�C��F� ��G(�{��f8�7��kxs@h1��wk�i@�5��d{��d�.;���GPص�W��6�� ��4�����R���G�[����ݕk�q�YT-ѥT��F�Y�$���5��ëF��r�i^�s9nsm�T?J�5�1��g�2I3�O�9⪾-A�H\��?��?�	�ؑ&BVO ������L����%�6QSRU����t��zR�:�K}�l�����=0�lnhӠ⋖�:�=/�ȶ�������ˆ[�t��Z/��d��/B?�o�	�̐�@�`�q��*U�BȄ�a���>au�3��d|�-��,�h��(P2�P��(�E��$�KUР��X˪lS��B���װ�H�]['дZ�Y���\0^+�bF��(H�A�7�&Z�Gc�}�t�yɐ�6مi�I�����+�������-?�N�괈�
�Jt�c|-��/p�z��Q.0k�B� ��~i�o8z�6��K�f�#���ۑ�R3-?��5��'/�u��y�V�Ք�<riYu'�ܼ�z%n�o�]�%��Q��%h��~��M��,ۻ�l�v�,z�
�Ū�_x�f�7P*�t��\�#��HA �k�K�����&���		ǳ���f�+I�n�ߟ ��%���dm-���v�����ï*1V�i���`�f��������h��@�޺0 �ٴ�W"�B��,��F���Ij�m���*UH�,6���>n���cAe�魼��B������9_֤T��lI�8� �H����ST�=�n�}��X`*xgQG���̷7i j��O�#]�}-�h�B�HEn��+�?7&����0�3���$�"�;d�O:H�&�|���3J��5K<����qԟ�:� g�/�2Wc�S�sX��NC�=��"�vG!�'��d�"�Gk�}�����XÔN�qe�}NiQ�Q�!+�ѳfH`'_^g$7vh@L0:,cd��^o��_:&���d}�&�S��� =��M�K&�ڠ|�Î��iq�,Ү'G�6�ؼ���7��E�X���H�m��fS���z$}}x�����jZK>z�F\\<Z���:yL������Ja ��i<1<8ɣ��h���-�u5Ё�Dn�	�6�IIr��^!�\!�˟�}���&�5��h��W��\�x��ˤ��A��=i��-��������oed�%�@gZ���*��_���+h����k�+]�y�=��`�ˡ�v�-���P/(֫=�)���o��.�'h��o��<��,a���-�o������#�_��\�ypO�	d
��/N�3P�0Ɣ�]������l>cx�q��2�����r���a��>9�R� �RHh���f�` .<�p����Ǹz��Q(�I�h����QAM��,�\>zN�b�@�v�-wY8 pܒ/XR,;��lx��3,��
~�>���ĥ�f�k��\9\��^���7�n�12ɇܸ����?�vY*��yMy�M=:9�\tc ?�1�d�����>�푝X�fsZiJ�
����ԝ�U���:;�a�嫡�.�09�)�m%�(�tx��?�d���C�CQ�RX\���x[�������\;�f��$��{�Z{�SP�ݸʆ ��|x�\�'�3m7vsT�FTxhJ�-n�%~�a/�\9�_i���if�[�_N��˟�� �W˛���@�}Χ���;����=�pcֆqy�C�1�}�$�aZ��<GC���7Y�ymF:��,x&�$��fj k���%��;�����n�1�b,�`�3*�QE�F^� S��z�H$"�����2>����g���b-����l�"p,z���>֦���:��;:u�Y��r�:��Gvz��#��П�]^Eo��Y��A�O���h��1%�����O�2�)Y�F"���,/@ bm�`����؄�;()�GM<�k۾�Y^6���h�eE6��qV������Ҍ/x��q�@�WGf$���U�h���~�s�4�	`w�����G�`�����p6�&��b�c1`V�h���ϱ[ҙO�^&�9��V�	��ܹ�:p�߬�IÅI��3�hDa�k��BQ"��Z�-o�`W���ԨW���:�?&mTr@Q�okF���w��
l4@fC�g�l�����6��e�i_��0O͸#�d��R�>A12f�q��Ք��R�D�8����䩣�D�J����V���
�CclT@]q!���F{�lđ	��n���֌ri �<�9t�V�B��j_P�nX�� ��ѵY��r��$l\�:�7�=��������+I0��+wl���ۦ��{��j��ҭ�!�0��)r�KvY� _�
�ѽp�ts`� <�]i�v׵������ҫdd�Yn�k��Am��S�2�/���ٯ��߅FysW4��}G�~��3��HŜ�pZ�����vu�/QP�
��@�����:Fi�h>��� ���=�5P�`>u����Y���ft��<zR#�O�2�8tL��y(J��y`����|hO t�6ٜ�V�ٱ�=a��"K@)Q�x���v>S)�^��3Sek"�8��5���R����\�B��{Ò��Pd����7�'���yyۓ�z�[;�Y|~�]�|��8���1��!�
�Ҩ3��MV��lw�^�3��sh[�y����`�'�l�5���؆��#X��-��2;恱��n��RyS�G��ּ�iȸ��u�l��R8���53��v^�Ϟ]y�(��(F����S����]39�Q��t��:Ąmm��� '�<�[�������<���U��v��H�ʼ�����Ν(���|ԭG3��zq55�q$޺Τ�Vg�w���2%�[�@[��Y�h%��uL���^�5k��Z�M��E�懽5K���C����$�b�g��ؾ��M������۱��zM��m���=�/��i|�v��DaJ:%�w�ꨉ�ZM˗�k0���}nޘ�"9���q��h7�1�U;#���|�&.�̘��k��.F�pV/��y�lȽQ���K�Wx�Y��x�櫉o���TY��x�{8M$�ϑ/[%G�u ����n6�d�5�����H�˟�9G�bv)v��]��:֒j��u�2��(�g�{����σ�Y���&�x�1���a��Т4��J�]Mh]>�zgW���hi~�CTh;3L��, '��p�qղ"��*90�SW�jd�Rb��;�#�/322x외]��Q�����Q�ҷq������Խ��ĉ�[<�=��L��U�T�R)�V
L��2~�)���B�و�\�44�(le�@6n��o;�Ub��ew�$��"b�Qjl1�C� �^2CS���L�p��	������X��&� ���r��?Ҽ{�c�`D�]�q�>=�r`����>9�)$������!��*�1BH]1|Ȕi�t��E[�>�.�	"�����-R�9'�	�)���0�]>� uI�9E��՘G;�:��LsFO��2J��Z>\мs� 4��,#""&d�0x������7����@vR!��@�7� g�y��bͩ�Y`�&�yxmNYU\�x.ǩ�U�������~;��Vԭ��T����>;ł�\Cc�8�PF�u�x�M���*AW�9��B|S}���z�+Z���.���r�f�wu��]�~��f�)�b��T�b=��F^d���=�{���U�`ү���	A�1D|@�*p���E��S�{�ָ���o�5������'�^�5Q���n��wXf޹�xa����Ӝ(P㻒+��xp�d@#�V�x��{;�-'oȓ�O~�sY�тء=�s�ۻ����+X:�HqZ��e�:��}_���F��k�dB��8�B�����6�9�#�A���Et�8A��0r��ʨǦ�dOHe��l��� ~j���s��K4j��G=	�\���;����SmkϏ,������n��\v�,b�����I'��J�>;��>�����՝�D¬m��۝��#�ή����qq� ��3Oy�����v;][d͹�ڢ?����wü��r���' h�վ���88�q���H/�f{��z�Q�0��ލ�*g�����/�b	�����r�\���}��^�ԧ�Z�W����ϊ~ҥ?���v��q���誔��G�.KL�@�b��>��n�x����gHct��L��a��1q�kV��J�j��޾~Z���_&fx9� �X;�\7X��z�V{�����tGN�$hY�>Ց^�����(}x��cM��N���rn�ݬ�,��=/zV4 (�<y��?����k�e��b�[�k�3�c�AW){�<�dZ�z=�n^��9�ɺ�%��4oo�l������k����3
4������'��*�C��\�?Ӗ�j��r�_����zw��3;�Al��r�=<$-��Po1�ėӒ5�g�w�� e����:��E)��&���
H����u�D�#�`��W�U�НS9SK�k�����P�C!��"w2�ފK�Zv���R
��z��_fv̾F�o(#i���]�1��xh�m��`����A^18]��W��`ژk�{���7�4��(��t��̴{��璟������%��gUA�_E�����?��8/i�sP����~��!5�"�L>�������REZd"�&����PEin��ߤ|�0Wld �>Fɪ�:��p�U1�kͧ��<�潏P}���&��~�$qе�~�U�� ��/t�_����޳�#n��k�5�N����F�\��\�#l�l�_���F����(/s��$��>|��$n��ݝ6���+.�_[�L��&��`5>shT�
(T�}b�\>����q"[� ��2�_$!&ƈu��WS��H��_NF���/�+QmlC�]3��U��h���7�R��w��ws���
T�SW�tJ��!6���Z�9G����1&��r��ŋ�i$���+��3A���ެ;1���]�Cm�<�3*�(pX���b�yq^D�:/�����-U��l�Z����ej�Kc��n�|��F˧ȇ��ؓ�B_�lNk�3�Dūb��u����C�@�1W���;��o�3�Ѯ�4�V7"_SDY���!�J��Cm�����b������S�V�������q'��g�nU�I�2A�d _�a���뎽�.��M���%Q�g��p����?#&������¿�����]���X�^a����b'I�$'s'�oSP��(���B�"2��*:�|ݶ*Ǟw��ܼ�Y�3���Ԇ?�0ӌu���i�	)k�I�}r���z�h��Z�ZsZ��F�s�r_x���v�%���S����1w| w�޹>�Z�r��}� Co$�j6@��;h)�����r�`�Z��$$h: BسO�.�R��R�!(�=GK��Vq�'����q�\�b�꛼���7�T����_���V44z�Ѩ���V����(�{V�O�mcQ�LѶ����	]����~�'�8���_{>_��J[��6���Mjy���GGs��o�&+��?���-}I����;�
ʟaǰ9�ձ�����KT'�#�=d�ڏ�TD��ƤVx!�?���&��9Tu����;B��ɸA��䢟$^���O����dr���/P�q��UI�2Ϲڛ���h�%F�}4��MU�X"8b`v� >j����d����|�B����xM�2:��n�Ql �>eӎ|P4�����Ǧ�/wY_*g�c�]4)����؛w%Ը4@�߻�iߍ'P"	�o��R�/�2�Dc�r{_q�1^��g�M=�^+���P,{�ra�V���	g��b��`�C�K6NA�0P�nk���J�~�$���u_jL��o�Öp���zk�;N��}��.�e�������ܸ`hd@ؙ�üjs��ro|53����xGHl�0�*���5Q�<���+4���F������ep^��x4�ݽ�MM�Ɍ����+��p)���8��if��*d�[_Y�P\1��d��D=��$W�Z�[G���[�Ř���U
ͫW�j�V.����2���C2v{�z;6��s7�-&P2�贿xS6�TbV<oӲ8}5���&���Χ[&ϛ7K����,�y��J���o�R�z\_OF�����sbw�P)�ٔ��N������+�_��/w���5c����5�)�� ��F鞙�ʝ������2}lD��ÐS����P߷[��Äw�?d(~Ƹ��y~X���ce���PKi�`}��
E�>��"D���Q��.��n�)�2e�;�E���)Lj�����2�� �	)���q|�·�W}>�������y�'g,�[q2���v�@�n�`�!?���+ȎOU�w[�����U�#�vqyLP놓����8f�f+���I�ur��J ��5�`���
0&fb��r�`#wE{2�Cy���cń��?�j]HzN˭����������J�.���@��z�z���a���l �XQS	�y�25]o�l}��î�8�L�@����0�'��mT�g���(gv�o�!I�-7��b��CI|���\�s������h���{GOϑ��ǕIPߊ��4�'���8��d�l���:�X ��i׌ǋn��K��h�!��Ρ�r��'��r8��J)�#ȶ���(�6֤����s��Ub��nQ�������ޚ_Š��NJ���8H���/c�ХP�ye�[�Ӏ��J���}�Шֹ�;��˸ⅉǺZ���rOl��� E8IuY���e�zΏ�B���bi��[���y_��]u���}�{��m�=�d,��;�vz��C��o��;O*a*_����f��7��[vdؽ#k3�{�M�S�\:H�Fw�E2(��j�Q�B>��ɓr�^�?z�ܩ=&�]�Iٔ��~������5�r�Dh�F�zĪ�F2��{�!6��F�����	�^��_*��}k��9��Nu��T\O�prl؋�s��~�0������ُT�%��KorS�֜֠���
��D�ӬvUU챷�kC�I�A7��T����k	�,�$��@�4��Ж1=0�P^��3��@����e����(d����-f�śdd�w�Cb�����ߑ�K��v�O�I�I��c��Å<c�\�=�(0�'o��0�8�m>�)Rcv�����K\�������su
����n�@��!�::�f�IT��c�Q�g)K�z�xO��*"<��p�ݹޛ�����l���\�ZF_8�������T
L�[MR�ZJr��;����H�̦�e��"��a�݊�ؐ�!j�2��a/�_ ���K��N������'$�֚'�ڪ��IՕW���L5���/��v�sƁ��~�{T?��|Ϳ�X�Ʊ��#���s���;BמF�w�9V�D�U��N�̕���=�Ew+���B��˨ڥܤ�.��U�4�(4nkk�b�6�+���N��`V�
�$=Q��j�?�!�q3t��������&U W��y��.�+P)�/�F�ҋ����+>��X1�	/����jT�KF�	���#�{���ħ�z�������Wٓ�]�T�������oI~���ȥ2i\�h=�]���f��[�7Ͻ��{o���@�Z���u�m�[CC�=���f����`h�hϳY�Ց+P�+��?I����Ű2�h1pXT,+��Pl9�v�!�c�'���Pֈ��c��Q��מ�qw�S��aj�/ˡ�w��8Wm��<x$�������ÔI'�^�~�Ξ��יq���χ;�:��&��J�zo���|�(�O�V�~�}m�M�����ʅ+~D��L��;<�!�Gu��l�]f�z���z{�L�6�[��O��R�t!"YYY�K���>����h{D��"�R)�\^s7߹��u�9��m2h��M#Ѕm��;C���^�z�����*u����E��m���4��_l�i�8U�6ӵ�Uˉk������D[#$'��莛&�iL��`(��O�ew�n��W �^y�4�sUd�;�o�|z��ʽ�"J�Ƀ|��X8��W�;�5&iW�jkݭ�9����=�:�Bj�_q�����l��1�F�."�B�IMz�s_T�YЛTU�[oD^1����V��4���X&=�i.ϩp�������3��5���m)��ʮ�?�2xf��'� ��[C�R]����՞��"#Dn�=~M�ٞI2n�({-�ó3k?�,�W��a�AC�R:�\�nٸ�}�[D���2x��oEVښ ՝S���r%�< 6�LǾt �-��rM��-1YB����;E�|��;��&�w4դE�/��5�YD�}g��鵐��z&E�r�}���1����K��д}��#��}y/6�����F"lx��(���yMt��׃�[�9�fƦ6��L�t'�tO���J�6�T�� ���-�Z���pڟ�S�'/9��c���9R���0�:2�����w"����#��-[t%݈7��)dP��#�L�<�"}��W^�K��N����wīX0i~ۼ~� �mt ��jGu���Y7��%���f?Rq[]������i�q�=���=�ĹS��KV54br���,�-�W�?�L�Z�~Gw�\��F�����#�i �׭/#��1`���QK�z���4�^y-Kg��q�����3vz8�
7��D	 �|��/|[���g��L�^�cN�#׫���g^��/��V�%�Ⓝ�ά(݂�"�վ
��p
��L��!	*�ǃy2��	c���߾�x+����E�e��;Ť�sNqDȰ"ߔ���0�G�"u��t��k�ӎ�x�j�e�,��R�L�v�~�/�$w�������| �h����t/Tկ2s�F���5|g����g#@��*��p=N�?Gk~��*�Lo��i�����!:Î�x�tIf
v�W3;���G�҃�uݕp�q߲,;�3�����ޭ����()��5K��e����l0�t寛)%�}
��F�Nc�)-������>�<��u�<>������Zդ{Մ7�g&�;q�?�S|��A�r5�	�'[T�EA�/���<�exN��*3�kF>�SL�M5�٪����kye��ɏ�#9���u���߻U;o����?7�G6�v~:��ݰ�n���?Ќ�Wr7���V�C�Ta^
�A�t��Cp�̚��k������jQ��{�ԧ{ޒ�b��kt���Ov��Y�;�6v'�o��Z7Ґ����2���4�k��>���A��t�>!�li�"���"��y��C�\����~4ݑ[U=w�+k�K�7ՙI{��0�/uN1��ŽV�:��9���=���aj,Ӡ���	 �����؀;��{Ey�%�e�U��;	Ǽ=T{�g��ll�Y�ϐv�t�C.KܹЁٮS�Y��d��<r)𶀝� ��*BI����,l�(s4M��]�J��oLn�lG���� ��w�{�ڴ%��F^�]0��������J�~�C�o�fo���~v~�F�ч�z�f��z@`��:9������r�C�s����������t���.�����؅,�����S���̙�s�ԗv��p���.��M��U��o6J�ì�U˜���J3g��4�]���4�[���!�;���E�� *pq�11v�3�����ҥB�/֛��?sd�l�����e�x����6�L^q�$Ȇ���Q��V�ˢ�*Y�H��d (fH���92*}C�w.��W�*����g�X.6{�R3��Ȣb�=��P8C^����C�v�qL�ªh��R)69��U>B�o�����[j ��х~���@����wY��'������_k<�6,��s��V�=� q�"�8����rx����^��|Z�L�4�V^��g�D5���"�x
�0��gI�ρ�(��.����������v������v�?T��䰝yh;\�o+a��9�&Ө�mQ{�˫�OŖ�w^ϻ����2z��+
�=��=�nt5���|E�D�>_Ӳ�,�?�vz^\Kcu"��B=�ɞ�l�v.6�.;��m�H}ŝ�������k;e-���Hs������ő_/�>�%Q��9����R�L-j��*Yt	F�`0|]v�s����i
�eIy�+�[?��\󒞚V�Q�⻱'�)-�0H݊�8o1rn����P�j�v�x�ko�����U"�f;!?.�7��SO	����$ϙ�Q����`sR~'���x�q�/���#�x����ٲ��w����e��윜k�z�d����� G[�n�{�"�5ۙ��7���e��4kҨS~ݠ}�R���c�΋��*������8���?\2�׸���Ιcj�V듥%8���/A������e�af���:�v����o8���]0���[f��^jE�YTo��9��pc��ʾ���b�W32�*�`�6V��NúE��W�[�5�E��3��VB�Bj���F$�$G
�����Jww��KF�����ހ�P߿o<>���׽�u^���sϹ���{b�l`�@����؋��y����k��^f� n�W��-�=p�S5t� \����E���C1R��+�*x�kט�:�}�O ��|^Pz�ܬM�qu��(��;��.Ŭq9�%a��C�m[�;�[q�;����[������M����[���mY��2�<�4!�I̗�o�Ń��r���F�K��=�Lb`L��+�@����j�j�8�0��<�A:���+ڡJ��p|���9��lV����Q u?,���w�̏Ayzf2�����K�9F&T���M�'�wx��Io���G�6h��.	��X3Mz������?�Hñ�~Xc�$�B�m|W;��w�O��xP[^����zW$�9����$K�dX�{2'�s��8�|��>�84���L���Zr�țH�2:t~�ǻxxl2��+ZK^t��P���j�?j���gt��D>me����,SE6w�ЉA��,���uƕ~���X���}+�ߥ�9��o]��+��2+�l��1򶙀�z�O���age"I�"�f�� ?u��B#�G����XWY|p�����P��vH��_g�OFX2����MHS��3?
fȔja��fJƫ�Vm��8gN�4�~a�>����f�i f����KJl淾����?�0�(5��!5F#���']CޭSY��)���ӈb�f�¦̦1�!AQ6�7\�(�=�T�a@���9+	�u�uF�����܇lN4|ڥ���? l7��4YQ�2&8�x��"cQ�'y%<�}\^[Of�i)n�?[��Z�шC���� �R3�i��ڴ�ʏ������eN"P��_�R��R̞l[e��(�PZ1W'Gh��[+��-���s1K<���d��_���I���m<�H5�5T\1L�"�&)TzJ*]H
U�%:��CzM��P��|����z4FƆͨP�x�'���@Dd��JQ�&.�b�h�<��,=��`������T�vE����R-�V:r��ÊL2�_U)��:3�`��,�ZQ�O�~ՑZ����H���*���Bi'q7;1N:�YM�	-%����J���l7���{��X��֙D��Ż#UlA�Lu�F\^���a�UX��ū��5���-�q�9P�������kk��MBY*�3nh���P�ԃ��z�K�Q�FH��JJ/��h!�vn
����R�ψ?�P�p��Ti�M�G�or�_1��-�Ŷ���7����vz��hM+s�����B)k��J��c�q
l��;�f)��R�<n.�W����E���8�E˶�j�	��Iv��:gyPuZ]gMY�pL����,*F��+�A#����j��>fE+�t+0מPζb�~>"h�.cĩfV���|߼�xew0cx��ƪ��E�ז��;�����G=��`�(��^�y~7�{}}S�l.4×ҕ�]�q�����5�Dv���� Z�b?�mt8�T��b�X�����FXw^�.���T����NM*�f4���o�\e���n��(�(8Z��C�~��Tw�J����,|UJ�J��}��g��2�z	"	U���~�CPJ�=7�Íɖ��sC��=� U���\���"�u�Q��FOl���qy��~��Ƶp��{�HG�p��8b��0��Y�oԁ��_�p�&����X�aQc�Ƃ��ǏΧN��W�Z��ȯ���t���>WV>��X���Y��`Ŭ�*s��~އ|��q�8�3٥eTdӖNm�L)��'����m�NX�hr�]7I�����Y���C�}��H�E_���ވ���1�=E2E��	A�0���J��}�-�ePڑq���'�����CM��O���?��&E�LoiD��6a>9[Jw���q�a'�3��.c�y<�<	�����Θ�wa9�����~��yχ��4�藡��g��p٨Q��,LH���*�2FՑ4��]�����5V�l\5�Ͼ
�
�p���	�h=���[c�.J-�����N�|c���x�!�n,�O"o�Ifl�Tm�-�� ^�&!kD�������x�Ȟ{�m}�<�`�5��#G"����b�|ԏ1gW?�$�(������4������&��YHx�S�<<
���Atÿ�2�}��Ⱦ,�S&A�5U������T��-y��ڊq��*��>�> ���!��RϤ�,ݙ�~���N�u,��sD�gt�[|D�۲{�}9�Iu����jֻ�nwµ�BpF"�F��	!YJz��k_��^~ ��6m��Nhr9R�^y�:Oc��b�<�Ps�Bx-<Ur'T���B))B5�V��q�S2���+5�m��-t��C�����ςxn�ܽ�5�b|��Eځ�;)�OB��'� ֊�S��ܸ��I�U<�F@���g�'[[/7Q�Q�3_��w�v"�q�^QЕ�0�'��{^*�T�����c)fV?��*�U���[K��P��띮����;=���^]�7F��� 7�x86hۇ�ǎ�^"�*J���?�F���?�\�eՙ2<[~��x������Ò����� �a �$��2)�0l��E(�/��P���Yfjţ��i ����̻BU�]{�hQ�K�� ��γu��}Ղ�����uƑ�m>y{��ڂ�=iid�v�+ʿ�k�`��Q�j�̚^AQk�N��2m�횕� 1�tQ'~&�U�
j��� ���u|���%V1�$q>5�Z����<N�q۟xZ@B;I��	�
�$���ٜ^}=��5�*Y��@�=Ƕ^`��d�l���C>�-�m��7y	�nR��t=|=�v���۔�7��Ѷ�mL�ɭ��z;�]��N�½����T/7�((4$=��ۭ����d2(O\Hҿ2Ȳ,���=��M�q$+`�/p'�DWk8�D�Y��q�eyU*a���Sp[[[����N�?;o��i*��w��[v����98���v�i��#ބ��}aߒ�7����'ͷ�׸C�^�R�9r�Ql�'�C�zR}�Γ>z�4wm� )b�#�#���RP� ��CwF<͡�Y�W$r�V}R]�T�D���_�b|PH��)h��_�9@0A���ϼ(y�_�,ភ,Y0���{܎9㗝�J(_/�)������x$�7m�z&8�|�� �|/}�酻K��;ٞ���Ӓx�0��u[�5���%�β"���DOx���b��9�H�\�сî�ae�3��3���l���ʔH\B�����}׃r��NsJ��j���O>'$��7�z�G��p璮���nk��/̗��~J�]*���+6���K�B'A�fR��$���������'�8��
��p�<*��S�S�������w��d @xeQP��/���j�M�s�W"�v.���[k�Fμ�R�4h�[�����%`/�pb��b���$0/����(���3c{H0�G/&Y�c����7k���fl{�)��z�vz�1�8��~��<�-��itFKzaj�M���V��hf�A�s���A��\4>�x�|J:qV�
��S��G�$Q�ް�6������s������}>��1�Z���׹�ş!M�������O�k�n��Q0g�*@N��m��y��-}�-�!�vƆz�w�w��&s��ʘ��=�|�+��i�`-��������My��KE� ���$� d�����C�+�ז�Ӎ-�|�l��(��W��:��d]owI.YC��94�D�+OX^kɞy(�S�!�ͷ��G��������U67���Ư:��kխ/ ����Z�T�uG�ۍ�ӫ� r>|h�����P��V>a��+d�+�ҋ�6�fƨ�������v?d��s\��y{_}�E�](�()��4��)����������4������i�ɞ1��n��~*+
�N#义�@T��D"vΊ��@�Y�.�y$����Y�S�����(�Q���*R@�^%�r��s�H^��wb0�"�'����~f#��;k��c�8�,#�]�>���n��E��$7�N�K{��ΐ��r�����˶e�6P�D�Ojon���~x�����?D#�9��[�H:^�`O���%��^K�	npſl�%�0�Gi����&[��`.7�y8��if̙�������>BS�%.7i�gFW-��G�.����-+3�Q�[����@4t�x����o�����Ic��Y5I&o����"vǆ���糿�ܻ�v�6�m������?����v{|��eW�` ����FȬM��g�2�oc:8|\Vy���X��H�T�_L�5�"11l�"���ة��X��t����Qӟ�@��#�ѪbLi�i�g���&.�y�U$�w�:��eP���L�+dј5m�Q�~N���3����2S�O�͏/�M�B��]$GK�.M,g+���m�f��M*�Sb�7+�-wqi�4�U�o�{�G��n��������P���i��h��I��ǎHIheK�.14Q���}>�;_w�2�[�̟�5;c�;�S����m�w`/�'6�:�9H��5sb"�ؓUO%}My�l���35�X�O���i���豈3z�䀅0ywku,j�U��#����ʎ\��懮���7[�^�����������x�/Ǌ�m�B�u��f�Ƅ;���kƱh|�X��]�Z9��+kZ���6��{P��/r)W_אB�3�M]Z!���G�f��� ڒ��h��I�v���"=��NYx|���\i#b*�h��'��2 �n�O[����?5*��֖��*���Z�*��>�^AAӃx���WT.�C���6��2<��m�,4bZ;b���7șϵ\�m-��4Ɋ�ۋ��(�ppY'Jf�ݮm$ߊ�tT����Ѻ'p�1�4�bPa�4��9gK���M�������Ⳕ{ĕZW�J�W�k�"���w���J+c�W������<�"�a�M7�I6TN��z��)~"�����7��X�(&.w'	����"�~j��a��?F��n0�t�|_m��'�23;ݦ*A�~ـ����U�|��Ҋ���+��~)
e���Ee��M~BM��z���5/w���?ol��e�`C���\��6��N_^]��H�:H�;�U�@F��;��%e�=����+Pj��]�D�0��0<�}����d�j*ǅ�^����N�!�F�1�����1��u��A�Ȳ�:�K U��HX\F���5�6�@e�8��4jw��#|�c��d���N���-Tf�,�*�uBT�f���x�\�;[��!�)M�{*|v��j\�:�Km5�ba�jӟ�=}d���;��?|k�O
��I���eY��2i:ZqI��GFF���J���~�ܑKF���9�=���K9�Ǻ_#�os1?�J�x|&j�*���~|�|;��)�H�����V��-	��쪵ǉ.�/�I_"8Dqܿ�0��&ʦC�|;�M�fK�z/�IH4��o�ۓ�?6r&q�^�=ư�������
ֆ��ğ�����9���=hB�H���,��O�����=Ӿ������R��x�cV�����Z��HR�Hy�/�ޑ��+(ڢ�
:�&n���~�oQ�i~�o��j�@O�������n�h�KOu��㕺{d���#�m}��q�Vo9��^��lY�и��{[բ�����K]�#�������������l�+}�t/O<���( ��K_p�o�[��f��)2L4(%BX������8j��S[�a�|/3�Θ42tugm+�߇� N��� �5�=�8�5S�4>±�^�|."�*��=ŞR�2+�[��3�i���A��7�$sK]����N�?�5�n�xc|u��q�g^闕LM����s[��t���s3�W��*�e�wJ)��ha��ʘ������r��S����H�#������z�#<�koI�\�P���h�e���9��L UmS��Yl-~���&�ilq�Б��~}�a"ՙ���� �Ξmi���WǵO՗��Oc�9�q���E��5��*��[R�� ����?����O�#���(�����Y���r�[�%]��r��'��"m��t�ʖ�|�q7��l��u�%�$D^�㛏RTB���$������f��g����tPW����	��yB&æ# �*�L����?S�?������Rl�R��%J���K�}w:&Vm�����<��N����8ߨ�JW���pg�����4S,U�Wn��:�}�����u,��gXWCH�~m<��'�ʹ�Й���Ɣȶް���6Qv7#��i�ǜ^��j5R��`D�^@�5p����2�3m0̈�Y��%�X%�t?�%f��if���1����l��O�ҝ��M1f��=J�S��{�6�n�2
���>�x���7a��ڃC��'�ؗ	�s4�'����,w��f�%�2|�(sT�#7�=+-��E�/&��/*�\��n0i>�%Y�n4֪��]L}��r�\��s�}O{").$�Oڧ��eU}�mʮ6�O�Nߎ$,>(�Cr�6M����[��7	a�ת���\�����25G�Gz��0�>����۱񢺤bL���ӗ��'��^ZW8���:+ZN����lm����	�5R�cɲ�u:Z�~c�w����gZ䰱��cj���:���pҭ�B�_���밓;���Xs܏F#xj�/%q�UZdBǟ�@�J� ��c�@��sV/��'��"��W�Pd����j�n��He�4U���Sꢜ���w�uv��W:kN��>���R�<a�1�nx���#$$�W����S~�zԫ1E�����	*�E��(��v.�#�;Ub�|f�:CZ�y8��i]L���y\eHv(���=�9�x��u�-�B��*:�j(6Dq���̴ۼd�I���,���9�& �)�E�~�0]djj�;RMx1��D��e�'l�Е��;�xF�w��ޣ��m��ڊN��^.�`�ck���#��̻+�Z5��x�l�o<�o-�]Yc3�l��k�m+�p^F��"�T��ɯ��Q:�D�5�^>�M<��M��xn�f�9c���(꧓D�C�V���A�	�5��g5\�/�tb�Ni$���z5gU�~�ܐ��e�m����t�&��y�w(���}n��[d"��}�FH������(����9�mka�ʏ#=�UsPg#xd�R3�ˊk<(���jp��a�<��Ύ%?o&��~D֒�R�ȇ��^���)���>�Y�o�L-�o�{��$���NTf͛v^�Z%Ia��M�ly0+��Ix2A��J�T����i��q-���Q�Ɓ��[O�Ù�`�Y�X��w�f���%՚F���ᡡ� c�Ӥ�:V�￼��X䔎�h�����N5��,�`9AQ<jH�d�>ƛ���5�{�J�R~��.R���S&E�Z%bV�\3�� kW߻s��D͏/�^�}���;u�yd�x����bo2ݠ���V�W���t�/$������5�/{bڝ�Q	̰�O=�c��Yl7�$aV�`P��h;���7f|)�\�y�ta��"�<��P�!�Ea#X]'l*6�2� 7e��b��4��^���Б��b���T�x��CdC�F���%Rvc7I^��k4�I�Hc��L��r*8�=IaѬJt(�<A��&Gl�!ˀ�#]�ᱪiVKGQ.w��F��j	k��}�|Dݣ�r�ݓ���l��~���L�~Y������2eqG��䱿���[�~z��j��j����X�)?r��5�I��\~��1A%�öQ�x쳨����h~Br�Uf�ؼUz��$�i��i0��Ǌ�D� �;7h��i�{��`j��Ng���V_�I~c�RC��/��s%�Y�Şf.������T��=�n�׷��x%��M	Ij=G��3Hb��Z��?��8��=U�
üx����Ӹ���̿�
}�|8��56AY
��K�<�/��V��]l�c(ސ��x������N�^"���.wo-���K��U'%�3���N5������=2�x�\��v�@�a�wT��t��-��`����+W:|���&=������iydy[M�#N��Z+l���%3kVm��? s�E��5�]�[8��p�a$��l�[�7���w��P���.�:�ĵ�"M�Ү#Br_����w�:|��No�"�� )-���U(�/%ѝ�8>M?�vC�>��@���_�Q�t����[��n�㟓�X�m�r*!�ʶ0B��[��H>�y�uvޭX!��!��� S��6ש����B���
�c^�P�Xp��R�}K��w���JW  U�����Gw�P��qg~�q�H�Ȋ�&=���ڝ����nJ���ė��P�����a�4�準��=QUc��T+:�.�3{���d$`3�RX8ۋ�	=�&l��fH��TȢ��y��O��� ���Q`��N��S�Q����i�^�5�w�/�~/7��N`L`Qk���T�����)�����& �ɤ�8�!��Q$a?��R��.��%�g�k}�������V��C�ɭ� ���]�Gf�tb�$`�]~P����]�b��=D���OIK�:�"lش�'K\8�ھ���LѢ�ݎ�g5��Z���`��g
�<�G�bU>�nL��l�fP�ƹ��R�́� ��/�����e��[kw����<�򍫠%��=7ĝ�l���H�b'��[��uڂ@b���7Z��t`Գ+�<K����n�(��Y��k���Ѻa�S�D�v�^���n����Ƣ�H���[49�U�ϊ��L�b�ê2_� +���
�+:��b���uuhKq���rk#h���M)�2$q[�]b�=���徜���4rh�&|a��{lh�]�6"e��M���+3m䅎O:�v��ߧ,��O�e��ȸw5=-�Z���5�u	�d�,�����bO��>2H:B{�&׽���h�xQg���$�~�:��葮���d�����9u��#��dSzŇ�	�-�8>�fe�Mt;�5jJ:�����#�u���Z�R�㧩� �� �f�^A�G�� )Py����4�����x��GH�U@ͭu��;�D�%T�-'�:
%�W�T�<�_��_�hD��;��,���@����Y]��_XN�"�����cf��^O<���&�D�m����ID�V����S�쬐g�P�Ő;RQ�u��5�'�Vb"�S��U�����b�����(O��C�e��<]�|�����.ɼ�V��ռ�F(>�#��X`*ꮱ�	��0���>Mi�g��2�s�(grN(���1��?�"��[��oށ�e^�g`sI�aV�b[)2�zΎm	π5oE����y�w̪�����OU�u N���S1���%�a�뿾.�dM�{֔pel���j�	'h��pN����ޢ��|oYݗw�&.E�Z8I�)į��������[��5{u��,�FR����<�(��H����8e��OT��������d�x�m�{P-Oǈ7�K^���BC���ł�9���)���:d�R9u�ǔ�C���5xIn� h�mD��;r��l�����=�w�ȷP��X&�/����դMx^���T�\��i�E���p.��Ju۫2v	,�ȉnE�mѴ�j�h�[K�g�������[��k������:����K��U�#�w)�c&z��Ǫ$�I���\�Օ*�o��n�ص�(q�"@bͽ�w����_�	���骤M>���ګ�ԟO����:94���Tz��K�>�c���@�P��XCq��h��}Z�=UK�G��S;�,y�3͍&������6;,���}��"����j*|�/�X��Pb�o���\�5Xx�aDc~���X�X�X/���;Z;��.���B���m�;Q�8�\�Ep�����UT�meo4��˫�Oq���A�"�{�~:����k��C�pW��YXq�[�eo0u��.;8ܯ��ϡ[�n��G8�L�e�)��֚?�naee���zK����ȓ�O'm��<�Jg�I{�Z]���{ځ<�u0�G�"M�/�V�Ty���
�ք���9��Sz�R�e�,�-�y�E��r������We~��\�Z�YG��r�D �!�}R��c�s��C�d�rV���Q��:��'E�x�W��!�Ԙ��k�M�'B1G�&>3k�2�#4F��i��=��¥,�aX��������O88�����H�ɐ:E�������N��S�D|g>���+��rیݙ�b�HL#�����:��E��L�/�&�R��>ʼ��M8��2�j�^[�yqF�$�r����#M*��wcL�M?��</RM�@�/c,6snډ�d���x/X��yd�af����S���+:H�(5������ŞR�1��!�u�(�j/yg�����C� ����p�բ�\�.5������(ђI�[�ފ��r��!Y��1�醗l�ɏl���]j~�A����J,�{�W�J�zh��&am�X��ݙ���o���2s)��+4��97Rݧ��9�.�Η��ܢq�ɵ��<��d������TX�I�D��˷��>�D�R�����b��ˍQH���ƩY	r����,0&v�\�
KNH_T��T�2&g�:rj�;��d�G!*s^�uа=�4�2�%��O�g2߰���T�j��q��Frf�CU���D�G�pzS���׻���""��[��,�J��蟅�Ћ}X�z�H�`�(�j�hy��R�<��KIۓ��&�7���ٕ�3r�]��n=F����H�YW
A&$�B��5C�����b]6�����=#��߼���ﲳ��Fk(���:=�L^��x&u��A)�z�hT�J�#�XE�����`?���z������rr�cz��͘���7Ό��y?��u��P��c�Zſ�%/�zg�D�3��.+��0b:�<�������D&P���tZI6�����]p��$?>^H-c�l�[S�M$�`j2��j���%A�4Ӂ��7�})�۪��ϟ_���[�����<���,,�B*��`w*%J�Dx�6V]�I'�X!}�F��9�`�4�H:W�W�I)�'��f���LA�As��I��溻�/�y�?������Xn�N����3������P��/�-u�(�{t��{Պ�C9{
L�.��-X)j���')�� �x ��C�,G7�5��� X��ؒ����!W"W<��P ��r6M�/�ëټ7��h�Q���}�μ�wFᝬ�vt��0�� i��a}�|BM7��O��O�ioo4d���I����WW�	^+��Dk0%����hWp����g���r��Yw�gKo����G5�/�t�~$s/�����<|3�1���0�D K6�����Z����-�R����x`{�:��	CUC-��',�N;9Q�mEq�]�R��[��m(���2���M�\<�&���q��Y����fj{q_�h��{i8�f� p}��[�n>o��o� h>��&?�������O[�+gq�������)�T�����+h��⡿�ͬ��(�uk9��������,|Y��(�h�	�����9�>
������C-t�MЬm*��]1-�%���f;==��p�%f{c������)j���c)��Ei�w6��滔!�d3%R�l7�Ή�-0��v�_�����;w�z�����8kz�Ii^VY �b��G�Ũq�N�d��#O+}���[��n!btܗI��
�&h���4�\�4�Sn��I�1{�VL}#{<��i���䣶{\���
��Q��n��ߚ�:����"b�;E}�	5!}�K|W�Yg3W�Km�I����͐G/�W�d��WE
�O6��&$���V|- ��X�����O����j����;M~4������qHC�o���7����
K_�~�O�X����#��y����N��ȹ�B���O�8�3r���o}	s��N��%��YҼM�72�Լ�'��w0�U�'&���=����?�9"��Hk[�@f��|�_C�T%�÷ǟ��e�Y���
U~�\0B�]�m�����mNL��������38�~���vr��c1��ƃA�ԝ��/�oI�ѐ7�8<*��\#�{of�L$�=���������:���׆����Ί��*H(�#ض��m�!�\a����9J���5
�����Im�DJ�/lQ ��U�R˜��<������	(; �6�t�q.�9�
CZ?8�=tp��+��_�&)������0/��?�4��x��&g.�FY�׶7>O6�U�߼�I���X�������1��_�]�r\ƾ�^��'�\�q9^W�?���7�QI��u�{O�Kw�di���|�S�s���g�o9 M������=���� )��-Q�v齠|������=#
�op���-��F'Չ4��)�r��w��*HS�L����PK   ���X�1.:�  )  /   images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.png�yeO�-�Bq����.Z(�����-,V(��Rdqw�Xq�w�E�J��H����yor��͝��I�L2�|��d��5U�	100��0%����?t���	��h�#7��'S��s�A_�?��K��K���������ח��孧���-���}�4��-p%}��c�4s�����ݹ��'N�"Ł�`my�׊��Da_����sY��]��`�~!�6F��	q�8�1"&��^��.=U��>������6�^�>1Z���� �Uw���I��1�vd�6ǐm�O�w�#T�7�<Bħ�O�Y�5��/l�8��)��*�ǥ����K���f�G�Dn,*��:��֘�ݜ���oN�`���쪰� �<)UjJ+��-ݞ=�T嬞o����B����0��p�W�	RC��r��",�¦��e��7���P�A�H�1��y�P,�F(�1}O���6ez�>�uby~���I��ڷ3��j��$<�洀H��%��;ϖ�o�V���$�=�+6��� �0����@s�	h'/?4�M�ίC݌ҕSp�u�~���-���x��귾3kF�&�>9�ڭa#|gTLw�ܟl�5�aI_z�߆f�~[%tQ5 ��:5���FjH��������fQU���Sז���_�8�w�:+ ��/ʦ+n�q��n��<�"��Ԑ~|���:�4�1=�ݡ�/'��^�E��8�t�f�x;;|*��ǌL����������4��?Ż)*�9�/��W���/.}�i�d͜���Ss72�6`I��3�������h������پ��I0�R��)#dg2�w �BP�p�N��	�
2�6�R�h���[��[�@�X��(��
O� ��A�޸�������A�m�	�Pn�*E�'��CC*c۱~1Қ"Y���k
�臨�RyL"W�x�E^��x\o�<>�|�z3 Is��$�[�I����*e�m�ȓX �рH)4oD��d
�X��/"d����h��q��}_W. �4H�$�H��E��k!+�k��~��x*{���Ģ��-���( ��h��(�|��7X]D��L��oۜ"I;ZCo
w���;��-kv�5���ID�Z�'䃨#z��[_IY .����S<_����cO[��u��^D����T�yc'�n��N��Y�C�h�ؓ��T��Ҳ���6-~�|j�������\����4�L��%-Q��ٔ�VZz�6��U�N��%Ď"j��\��!����u��I�l_�Q���w|{V��Ⱥ>��Š�����n3|x|��w��r2,p����m�W��s�I)�C��;���T���p��P�g8=�G�렶d��(��|�T����-��iķ�\�d�/w?Q����6��#O�?���ˈZ����c�\֍P�}0��G��۶Yhol���TC��F�%r'��l֮��o�x_���_����GP{0/�Z��Ӭ|F�L@a�.��s���|�3;�٦9���u�%z2=�9���wD�Z~"u�Nk��1y���5wϠE K�<�zzzB*������+��SR~����	G� �yw<QiG莆�������ʭ4�K�{��u���j��Ѩ�ft����q��42>V��CVo�!n�B�����=��!���_ʕ�c��'6��~��f%�k���&@��R��a�5�e��XDo�{n�̀}�wǐ0d����̓ �P�:������jӊͮ�!�Uu�7�Ќ�^o�S����܀��eI�s��|7%r�TK�������K�du1\a;ֳO!�Fz`E�����ބ-�����Uv�����TƳ.��]ܮؖ��.v�bA��.jM�Ǯ���������.��<���2��{r��""��Y���&1Z����׍���u#��G������o��UE�;�~ʰT^���]2*-�J������h8~�����s��:��~�l�h7�Wg�%�`�	_��U��:A��!3:iZ�^T�)��ʴ8Kw4\-�/��~;��e+��1Z�9\�ap�pb��leaE�]7�@s}t����X���� �Cf献/�[��u��kF��[���i�e�`��aS	mH���F�;ўH,�Q}C>�{��gذ|,��Ŗ�`
9�Ӫ
:P6���%� �84�H4G�b�},V���h�Bg�\[��"���0� �o�פ;*��Qv������p��3w�����J�#�G'Xq�i����"����Y��7]���T��'+8�9�$_V�TN��&�|�g���5�a$3����ܷx�fo`��܉?O�j���n����S��+�^rA�n1�b^��U�"(X�$���5��q1SH�J���Ʉ��$K�Qq/���NG�O0�h:�}y�[�.&j� �+�ma��yr���5��З�(����WF�&x&�4��[@9�ɪ�tmF�	����9�E��~�L��$*���\d�o����齬��߶��9�V��@�V�����'yG'X�R��M;�ˆ���%>/�$�� cv���T>��~�I_��~Z�Pv�޳_g�d�
U�/e�p͇����3�s�c�*Mi�!R�ث�8Y�	�N��YSud���d��y[�l����/XJ�v�)��������ٔϾ�fs��a��$�g��5R�����?V��-p�b����3��z'*�~wWe��F���9����W�B�_ZL A�,R�B��,zֲ]y��^ԺR���Y�z���D�J0I�"CA�����0u�]lC��j�� �Kr^!�������Tڸ�8���ϰ $,S����W�k�ì$*�3��,�0檋�K������j��/��s{�É� �	*̓�[|����nM;����3�+��V��G����<�0��4Z0�:G��Ps�Na�:�`U�z��������,đr@(6cV����N�ئP��l��;SE�6}��F���}[UC���v��Y�?6�j��\8�jabU�3�AD�?/��s#���7N���B�Cr�C)=^� 3.�_����1�c�1�t�I�9�t.�`4��
���M&q5�ޞ^J�Z+��1t��8ii(os#�6�(�g�=ϲ^:��Zc�����O��q
S�����!C�*�]]&mQ���%?"_* C�E��#�
��J!�F�]#�L�-s� A��c�t1s�[vn��qۢ6�.�cڶ���7��~jJ��:z�6�A�?B)�լ��c���n�U��ceII-�t���Y#*������Kuv�:�x�<�S�h/\�C@�Ο��˝��9Z_ز"�o�� �Z��].�9�ɵ�/�W����"jQ-�0�+UOQw��8%�ERV�.EbM�J���b��[�AA�&�Xw���5�C����B{�"����R7���$c�R�13���?.�T hS��e٬H�e���̱�*��Ҥ0�D7��(TC_�K��&b�	����zX����>}C��}$c-Ag�H=gwٰz����4V��MRp��ޞ��B�������lyyb6d�`��I��E�d�K�q]p�d��$��U�H�L���D��� �MY���Z�����*��CN���J�[��5KK&�����Q.4���������Kk��U�t,m^}hg�p���^ϻ���Y�6-�ݓ2:N�i��{QK1�@C=�0z�Az�=�PL!´��G.~�:	@��*�{��r�d��%^)�����������/���Ո|�b�_�n�d�'%�%�|��_m��zKW�#�Cͨ��9����I8d�봍��rS9�ʚ<gX��a��z��+�Q��|�l�,+�����U���ƉP�B�Ix����uX��с桨�y�q)>M6[�d� _q02}����IV1��Z�YzVw�|*������\E9L�%|��&���OI^/���P��'�q�M)y���(o�F�����A�3�^(~n��3��¢�Mbt�Q�0��[{�	��@�8���Յ�^�e��5�>j���^�@iI����w�w͜jG�RB���,���qK�qK��_q3�c�	!=uoGi�,���EA4�kk��=ҢB�}R�e�\�ቀ�]��[b�������)�j���#�&�4.�uu-�!�-�T�2��i&ig��p����������	ҙ?VA�Y��^NcU(x��J��ѱ͏p��ص�sf:��3^~#�=2ܲI?���嬸d��xN,��ΤL@���rl��z� *�Pmq#����__7 ��H�B<j'r���I��m�H�3��\�hxi�[�q�ӗ@[,������%����b]�pvR��Q{��̜�޵뤗_2�)y��ѝ,km�R;D����2]�L��R������n�h�9|X�q��a|i�
�W"|6^p�[�Wȳ�븅�`<kN�Ә���?G5�^l��2O�V��]7	��0��m�:���PY���&�%	'j"��,3cj_Ns���+`qA0


M�z�ax�(�)Ƀ<g�5$�0,�t�<�1ֽ���lj(�`/#�g��}���	,�}���8F�&�b
UQ��!;�b�#b'���dV����@f�(���\���S����#h��O�:ݼ��a�XVR}i�һ\`��\`��D�m�K=���}�ITw5!��	���
~�n`()xz=s�3�.B�f�X�i�k�%P=�Ԋ)�jcɶ@��q>t�M}�K�/xW��Iuk�[90��o�A��dy0*�I
0�Ά���}3�?�O�V�m����|4(�e�OӖ.��-Ɨ�����<��ϱ�#E��x���i`C+�D��+൐��T�������1r �^NI�i&c�u	_����xi~��j�o�t�>�d�S��,%��Xd�z�7i���C�_�{���⢫tA@z�.�S�}4%Ь*,�{�4����Dȩ��L�I���%K��g�%q���w�y�_�c�{qʺ�L0n"/�����zt�/0nGt��d��G�=�x�%;9����=�б����&�}�+�m��s_�l�bV��S��;�r�9�.W�i�����F-;6uoN��I�l��i��~C�"�p8�C�� ��؎�הݮ���%���l���ܕ��1k�:�g����=���{������G͈ne���$�(���^�������q���[�N
���D�h*��(�#Oht�aq�|*�t4E9��mK��(T���]a����8���f'��)��z��������\�t)���'�����`05�t>���Mt�=8mx�U��&��@F�<�)�^|�8� ��w5�j'�=�M�w[�� ���&�⸥��n��Ǧn�!��~a����y�
/����'��ڑ�9dW�����2¾5��.�#�쪩͋�@Um���ZlK`v,�]�#�>�7�1�a�d'�#��F\1�c󱢙�5��i]) ^�8PHN�=�"�D1��ǥ����аf��_3I
�G�$"8�0%����������������[�!���8r�kB/��S5c@B�ND��|�X�2��v,����\�)a�]���d:0N�s����o��\��ʈ��Ҥ�!Iu؆Vs��*X�tq�֗}Ȩ\��a��n�ћ>�Vt�ye����w4�F�)����n��oW��y���V��D�e�(/N�#]`z'�`P��ec�����H�Ħt�����O�]��B:�S����I�a@)5�J�z�@�%��9���Y���\�+���)��M���
J
G��y\�Z1'�Xߌ;���T����yS8����:j�!0-a�H<8���f�$��i+ç�t���!>�A-��\���ϵ�� ;��3��4o�u�Iw9f���f�4"�h�m�$H!{�O�g�c��C�C�)��ঢ�S��"5<���3�o�9���fK�!.�������f�^M�Y���T&۴Js����n�"��B�|�o�[�9l`���2ˏ��WC5���-�Z�C���c�zo���=^t$�[&ˑ䨤}�JzgM집D珦=o�M�[N��p��2�u�kx���ڌ�Ȱ��y�+��.�T2-�SJt�-�k��]��.��0zX�h
��ڒs�%�E��>�e��;��ã�/fMۅ�]j$8� LA����F�TM	��{|��EWՅӀ��"�õ���y$6 N��jC�^�&^k�DL�Л鴯SD�i�yr�,?PC�b�^����N�y�P�tm���� w�~�/q㵏���&����Uq�б%@������� �U;��?oT�-�S��4�j����JX�/���yH��v��Iĥڰd}f�kه[�[eo~i6�y+[�2�Pw�2Md��7"a	L�I!$����GNqZ�m�8qI{���;Y��l]�u���������Yʖ+��_��y
�.�h��f7z�\U���}�S"�y,�fP�Q9���5XeYL��?�.�������]���+�Z��9�j���,�S��~���:�=��������t��P����E����@tuX{V8z?Ѕr���k����7����+9�����뢓oC��f,�QM����E�-��M}��r��$����:�v˝�G�4�]Bp)���q��-�o>�����*֏���ץ�R��-�rc\'���F<�"������\t �$m��@p$���]-8�	Ǜ�&����u56CӐ�Q�� o��j�}||}Lk�ů�H˓��W緽 �.z���l�p��drB�1-E�� �G���v#q�߆�[��׿_A����h@f {,��ӤB�0�B�+9@���ȉ����2%]<�Ǜ�9����ɤ�޻��
"+�s5��I���N�t�{+HI�~���Vr��� �D��v<;�n��S<�x�4�at(�B!�n�#��J;�������>�Z˔z���L���:s�	����8���8<4 /���q���>�5���^�P�1�C0˓��2o�y�����o�Q�,VfϞ�իwCR�{�ϐʃo��*�� N�Z�+'M.��mݏr�)����(u`�{�e�M��9|����/GD=/���BJ9��.���{�f���������(��5a�vx�&�V��<䒛4���I��6�K��e�/j�k�Z�s�2+u^�����Xf˻��{k���s��ZY|u�F z}R#��O�:�S_�E�����ho�lW�;�T:��z�K��і.� ����mjr�b��lT:�˒�:T����Q?�y_��_C���]�3�^�I��.�$t��@��K|>��+�%�;&`�1�έ��9�s�@�TN�_&C~ͪp�Z����
HwTS��L�Pq�0;m�i�4�w{,X��+�� ��$�uԡ��ۧ�~{�Y>	#E;�D�YUq�.%�[��E��S�V���R��n
��O��:t�m�D�6TѪh���lF�J�ُڇ��Ev󧟿�
���/�������\N��#�_ J�Za���/�J�κ��Ȕ��w�QI��dˢ������j�%a�dP&���GW��W5v����n$h'Z�r��Q����R�.W?�MW� �Y󜖱���A��S�_��%=x *;��f�eA��y��#&�}�>`�k<+�z&�x���AC2٩���}ŽQ}ָ`��{�T���+�:�Q���}+e��T?P���L�"t��	����-T���hf�[KzGd��Rʦ��7�Ü?��	dX`M�-V]z�#��k�����5�>C-C�PK   ���X�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   ���X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   ���X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ���X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   ���X+L$��� �� /   images/aad47697-5cf4-402f-a095-abba84463b41.png�wT�i�6��;�#��*��2c��T	ő�z/�k:"U 0��@�ޤ
��z���K�S���~�)���Y�k\�<�������~��B���_X~��������TTJ��~?wx�����/���T����[����j:QQq|���{�����,�tV�3sF:�R��h�W�VNƆ��|v���dq*�_�����*&a�ۙ3�%>�Or���������~�����~�����~���������~�ȾP��~�����~�����~�����~�����ʾ�?��?|�p~̘�����\���*�Ηsp��"��'�&�m��׳���C�d��;'�G�=�Z�(���/l���d
ʜ������K�Ͻo<�J0����̚��#�s>q@�}�OJY�n������dR5�/�|�(��'�����ȏ�c�X?֏�c�X?��k�'����?����=��$K���8b�+Y���L�ug��J$L�R�(���2R�]�������²��7�btU�謫4�
.=>��~ӹjWS7�����y��|K�]U����Aw<)�~���w���WK����b��yf_1<��i��\b��}`�/.o�U���(��ͬME�������Ͼ ��+8M���R���XP���m��FC�����Ж�D%�w��2K��e��7qoޫǉe�QfH>_'V�%�oכ�)�p{��ڡ`FS��GՕ�ᾰi�)A��+O�`�+�ع����U�&��:��#�S\-9l60�f}u�����P_I�?A��4�O�����#�W;:Hj����Deg٧���S9�C;�IjE"w��)���0	*0�du�K9>�~�\&�A��L�#��|���+�R},����qM���딴��e=W���a���W]zx��K��G���ޑ��:��=,��j*0���{t<H#f"��rT���
t�՚^'��k<�	7��xn��_����8´vsa�r� �߬:ۛd7Wmv��V�#�u/B橉��x�p��&�r��ix���v��Ǹ�#GY\��US����d�8�Gf�`S�����y×3���O
��:
�F��[��{�̱�Q��.Tb.�d��gh���Q��aQ�]��_��|�Ȕ�[�H{�ȱdo�7cγ�5=g:Ԕ�X�e�+�e��ӗ��ĕ������h
y�E�6�G�g���K.s@�'�K��Wk#�\�ʑ�5~�7�/�ݮ���*��Xֶ�1��\����xޤݮ\}3-���\�����x��~޵$��"y���^���=�}M�4�P���=H>�`o��9�/�k��i���#�B#(���z�~⍄��Edt���'as�
A�X�G��ZM;������{�?]�����	��,�N|9жo�ޑӲ�[��n���x.AO�B:�F��C��7�D���;��2+w�}����g��+��fHVotìkP���Â��%��a2�p��M�[��w����#�������!v���,�$�.��� _�����Y��� 0��uW���R�(RN\�M9� �ò�eūع�����7ޫ|w��v"l���ðw����Z���o�yb֏L��ߍ1Tҽ%�O����Z�:�*��\�)2�w����eb�x%��T�O����&γ���hL�l��Ói?�8�S�S�E�C������{p��s���RS������@3��9�j�㉪��5��5�#Q��gGM�\ݘ�v����;��3k�H�>��ZU*z�[�|��>ʾ�Ԏ�N��e{U��`,d�愈���(���P�lA��K�y�
N�#��x6��+��hQ�J���8׆-/���c�=�?4ݯ�2O�1����lP���[^�K��C�h�Wp,�*A��K�d�mx�N��v/�k�cg*��j�_��t�撃�	P��1��Ć��m�d4u��e�1E���?����~%b��m�����P����,�N�N+$�� N0�1�U�8�lX��vq#����`o���nkJ3k���A��T�L�<ذP��#�[��'�g� ��ڢ��$�ԕ�f�iZ�|?L)w�u����2�*�$t]e������"ߑF�!�g!)	l�kʶ)!C�C�jQgm�g�J�'��&�����q(f
v��d�H�^O���f��yL�����HeQ9� fC�Ͽ�]��n�l��̶l�Z�_�Ex�۽���u�)+�
�7��ǵ&jF���"*İ�Q=��"^����°1����g�8M�j��|����g3��>�J(�՜c�T��kt?O�uU�����Z�C��:\v�S=���	."@r���ӂrT�O���3� 2���!��y����3Uحɀ*]Hyd��/�x�����0kBɽ�9�)�\�5�KFM�1).f�V�y�+�[��WnV�9٥_�V��+ڙ�-�o&�gM��{�����!������z��X�Y��ײg2#�T�e&�:;���f�k���uQ�S�
_�j���パ9F�cL�Q��X| a�ev���_T{�+m=>d�_t�?���b�./$݄���S������8���O�F���t#�F������vQb�򕸓���=[�i4��û&���ڽ��,ӽ�!q�}��(F*ka���?dӯTu�5q`vZ���mp#�N��9��-X�*�����0}�������ai��Lr ���mWg���IYm���Z�=mRyϘ�R�4��A�J@ ��^E�Sl���x97��Vƅ��F�������zեh�I	�vt�P�'�%�lk;�~��ɨ���`WԾs����i�^N�ڍq�S^��x�O�)�%���rH��\���l�۾s���^c��OT��z"���}��+*#�K���-�E�p�5�j���5�+�m G�~q�G������k"��s�뙺��&.��-�ʷ���b4�����Gl`9�x,X�#,%������T��Y���<�e�ۓ�WR��Y��V��G]���eȗ��L��̈:��¹�fqoCMa��p�����-l���W� ��	Ѩx}Kn�JL����,����9�k[��z3U	-�w�l,�$	Ի熸 0�Z�	�06�G�i�s��+�S&���6��n��(��@��j�Ż��w��V����6�>q2���O��+��T&�%�n_ߗG���$�$B$%9��H|ЮEP�>�ZF����k��e��}jx`mU~�j�y��/eAf�)T��ؘ��ƻ�,t�������*aBn6��X��n��;�b���ų��u7�K
��Hv��S����T��	�t����⧖��
��,T�܈�ւ_�b�'��k�|���(�i�iO��a�쫊)v�|���ηzV�
�A��h��K�C�wQ�s)���(�+�s�� �2��1��{�f�-�}�I�"��`��]\N�co�W�������`��4A�z�T<�<5�u+�[�m�Wo��.70)Wǐ9w���5wѡ����\�>�6��L?�:'�|�h�PP��d���m٥.�GY�g	K��_��v]	�C�b��`�V����%/��O�灐0��6��O��9��&@��a��� 5��8�+��\�����;u!�p�P����H�i1���x����FZ��ϣr��H�J!:O�����z���`3ğC;<`��ye+�^b�!e�bq��O�t@�*L?�%E�}����|���ia�P��O{>m$�E�D?��ǚK�ӛ����$��Y,D^�K.A���K�[����:b
�B
pAׁR��� ����i�(@��7��z|���:/WG��s����&��CH�~�'M�;Aƍ8�uo���0����"����Y�H��^G�n�fN����#� �ˑf�>���2�c��$�54�����у��b<[$2�{�A�t��:��4a.�k:��p���b�ݖ{[�ࠚ�p�q$AN�fh�j���F.oA�rF�g������ �9�P��>O"��9^�Ɓ��
�%ȩ�#-�M����W'	i�\A�Y��$���΅*�t�"�E�A7�FRC�Lp�Ǚ9�+1�ϧ�����<�o?�Q5�����e/�pm,�oz+�ٳ7܉ÿ9k�E���s���Uɡ�!o�����]w!�(f�cH�����Â��a�x"�i%���PZ�I~��sj�N��7t��Q�X���������'}��ފ=�+@��=k��M1܌��u���Z� �_�=ߍ�*�{vR�v�rMF�)fҿ�,`�m�,�i �(| ����}|q�s���BML�GR7��:/7�^�d��I�:f���g<�,�-���.yC(��qV~�T�&�΢�7A\��Y�
��uQ��t��L/q�|�ZuR��WZ����Q��L�7����#Ō�e뼕�m*����w�2�)
!PU�/W�p�ȸ�B.*��ʆ�6��k������*3�O��B���tx����!�U��z�eє�L�c��)��<���#O|�h(��n���9hâ�ⱒ2s�����O��6]�A|����c-N\/��h��:M&�d�vg��=�f���}5�W��rf�Hg�IW�]�0Iyu�J�[���*����A2�=��,)�v[:{�i*�K���{X'�����n4�n�v����!YS�`�~,��aS���;�"_�M�o�I���8<~n�G��%K�7H_I���KT�v>iwL����r�@����6��J oĥ�|�Jz.14}�1�&�X_������WΘ�|-� `��az�\vޠ�u#MϏ�7?y��h󛼚oREٓ���W���v�>�boxSq�2�?oN앁��o�۰k��Cɬ�I؎�����^ �5WT�M�|��;��G���?�6"�B���J�wt�������#��r����MO;������v�n[�Ȫ�+*�9|�j�e%)mƶ�/|O�q ��>��W��')�z1�_���f����y��B��ч��4ss�\� �30�y�qW7�_��/���{)�.P1��0{����m���M|���y�uMI���zۚ�H�R��$�4Th���O�i�������/{ގ4�] �xw6�ރHʼe�QF�F/Y�ߟ��Hk�ڱ=�|��==���8�S���W����T��p�#ө~���]��aq�|�{|��W��-����!3�Iv���N���o\YlC�Z򹛗��CB�佅�YXގ�X"��ӥ��C~�9
�ט�L6����{g�����JY~*1zԜu�D�t�'Ɛ3ތmF!��$�莶k��N)~�� jM��J�,�l��h>(И7ׁɯ��+!˷̵�%b*ˉ�Y�A-�\z��@OO�F�Nm-�XH��VЈ��3F�O�*����"L��g��c�c^0�5)�u��_�$emo���,G�1�C�q��1�������ݜ�߈�(��M�� x�qlb�_m�&�w�5z�,��C�&�{�6*r�RU�d�ɗ��A�K�C���>"����_���ʯ��C[EY�1�ַ7�vy����(�;e�C;]�Z'
��{�ϛ�W�-6$C2�3�x����93vF�x�OхS��wk�k@8��l(��ǵ"q�c(;��S?L�6m,���0�N]Q���-={ �?l͠�6/gw�4g�+�F�<��μ�K��%%w���TC�n[�|�������ea?��t}=E�-��_z]���kf�\M~h<B0��L�HL*�o�O��0p��.���f��EY�&��������oQJ���,���3d��'7^IA�XoCO�#_Y.�S�q��{tn��2?���p~�0�����w?gػ����Օ]��`��zKd�d��Y��r��#��D�h$��B���=���Kx	kB�)"1�Vy7=g��z
Q��V�=?=�LHh�_r���"����4�B�z��U��"+B�a��o�Y���>��c������ʅ��=��`�P2s0�q��av�z6��m����N	��R��E��a:#n�|9���\����d�'��Y�\u;C-�A��}��4�X�r^3�S�`ʐ���Z�Q<��5>Sb��X�EH�	���~a�DW/�d��-�ŋ�$�ҧ�i9�k)�=Վj;�>麨�1�Д6W �x#r��s5�3u�B��:��w?}���(Kj:�
���U�;~*Q�t����B�����b� �mx�	t���g�m�r��r~8�`��cJJ)7O������V��͇"�3���^f,�>µ��H���O��H�B�Y�1���x�O�0�)�:����(yM�s�.)$�ZC�Ȭ����!��Yܧ�3v���s�7>IA�p+��nJ�`���p��96N*��Q/0�j
�ǐ�fZ1��&��n���W�{�ǲ3���1Z����"�k�!�>C�<�K�Wz�7Nv���«�tbɤ/�")�aw���D�鍊g�,��*�IR��_���Pl����^�w�o*h�x�����A7N|~G/����o�f+݁>�R�d�d�-��d��R�OI�ba"��]&M�o�����OJ�ӡ��[&ꊈ�Sn�ʦ�d�����qrJ�I��K������w�f6�TE�AG��bPH�<<:V.ܺE�hk��cM9���|���~�XS1�C�R�2��^3�}����f�GU��cц|��Y(��+@ 	��4n���r!>���g7��|%8�ش���1����4��TkIg;�c�Xw�3ۄ!k�-��lo���C��0EE���{�!��Q�������cI���񳧗�tVlI�w`?�ƈh/���H�m-qQa�ѵ��wBt��. �v~����������1F��]_��'���E���ψ?�'9���J��,Z[��Y;+N��S�%�����[tE(:8m������g�"�hE%s���z9AO��۵R�֗�/� vW�O�N��P9ϝ���Ϝ�.�Ij��,oT5����bo\v�`�)vk�|�9��-�||_���8������ڊZzyh�G�̀��=�aŨ' CJ����E�N5ȗ�r5��NN��H�.��5rP�r�Bȱ�
�c�R��O��|g9�����BMTH�P>\��p�ˤ�@S���NTO�$�R\ʑ�.��8麆E�e��1�����d�� VyƓz�i2��Iڐ��a�ZJ)��P� �%g�Zݶ��A�gG�w�h.hc��L�~�˒�_������^y�r����)z��U��=~����V#���Az>%���ҷ�(�&��(�������w�Ps�J�c{�G	�5�F�v,���kP�St*�m��rJ'[��Rm��������h��G?�Ÿ��ny��n�H��fr9xG����
���}I��o�*=�F�[ ��L���|z�"��E��d_S��!�|S����'���ә ����k�����A��-�:�Hs5w�IW6sY��H����堯'T�"�"�6�7<��I�zI[Hs�-n5!��+���Ch{{˨��;y��$�.�5w��M�#/��3g�2�[����'�R�y(mSe1���}��x 3^�X'
T��[|�k�Y��IiI��ꊒWO=������6�{c�xE�p(��Y��J-#r[�ɴ�������)�3�.�sװ����؄�ն�N8O����nο��B�� �d@�+at�qeȩm��B�^$�Ԇ�(��Wi;­":ʯ�	��i�(O6l���L���6�w�P��l��V�w���Pf)���D����QΫ*;��#݋~��.-ʹQtvl�,":����{T�� �0��d�k:���o�`L!0��0���D$����ֺ-4�44�jܫ�M0?�{;�yq���}���{,�ջK�c�[��[���]g���OlSG�Dj��Mh����+�����f��
J�?�'d�<o��w���}��3�*�&��j
��g�bsb
봚�q��kO�O|*У&G�J�+����`Gw�j����Ɔ��>�Ҋn�<�����c�ׅ���;-ꗺ�%�!z��`|.9��Վ�bҸ���̟� �3�t�EڕECA柡�1����9!�r�DOM�.���"(�n�JTey8Z
���˩�c6[�ō+e=����FĦ9�����e뱱���ǯ��Y`�Hx��9~��(K҆��`⪥��0�R�N{k�L��wM5���W�Ym������G�Wd�|�o^���M���RXH�%��՝B�����!���w_�mnV'���f�� w��W�ǵ���7���cY��r-�wJf�h�0�c����I*���΅Z*�m�H����'�ls4�Tv��P0,�'ꉢ���`���w�`�0�;i�+_M5��2�2�{�x?���/��|�L�e[n�@8u�.d��'��4���h;����F{��8�%�Ks+1��Q겨�6���O�[��Qo	�l��� �B�+�W�xK�I�u��a�R��7x7�V4ὣ�����/���Sni�cG:|�\K�����W_WK�?R���([�],l�3rMĊ�ڹ�юV�]~�7�@C����?)�`7��}�T���}�,�#$�$Г����N�߳���e��=7��|hx���w����-�"���T���۽�Ǭ�F�a���8�Kz^f���irճ�(��_f���,U[�R�`C�E@C�qY�����ShƸ!�ɸ����_8m�aF�+��a�]�y;�a���?k�H�nh��aޓ:4�	��oIc������� @6�oT�Ӥ
�;��a��p���9F��cu�y1HQ�٧o%C��@q��Zc���3N���,ݥ�Nq�ec� �ym�Lڥ�j	r�A_9Xr���b㸫�0�Y 3I�������rJ�m^J77��m#p�FRB�������3箿�녲���Į���B[x��~ ��P+���-2v�,��@��]�ud;�ٰ���X�i�����k|%_��|�L0�E�jmNv��)x��G-��m_J��t�*�ɻw@~�q7k�4k�iԕ}�l��43#�����aJ�z�צ��~�;RmI.�<9�9 ���pȉ���8���h;K�t�I�z����fRT���U�c/�sM7)�����?���ƹ��N���L�����+��H!�dm�����`��[2 $��U�M�D*2ŝ3)���n�=��xu��pΏo+����2$���eh�z��`�J�ӚL�>#������;�����J����N�S��|��-��'�F��p%�&K���#�3��)ғա]�)�׸�O�z\��F��D�.ϻ.@�QDqe���؇�������؃&��ͣA��k7W����Zqc�����5|��Z�gQ�C�"���������,=Y(���4'��JD2ڹ�{Gpeʕ���.T�x��e��q9���=Ѹ�� ��`It^j�U|����6 ���8����*�`���}���3�R�I�X��/�'�zH�phC[R���0�KPV&Y7�"���ֱˏ�% ���r�'��\��T�^�r�=Ĭ�3�U�P���f�NT�؂����*��6j2L/�P̡!���)��Q4ԒzAT�T�wa������	����MF�k]�D "?��4�E{�a5�e�Ԡ-�ܩ@�R�u���ĄV���A(�^������&}�@���dN��PkY8fVa9������	���'	%��\YUS�Ͼ�eOW.��2��^��B`Dw��t�wA]�{!\�K�}N���J�tN�ƶ9�4�)B8xB�dfo��C��(3�/�}}����'_ٓ&i���|������^&HzL���pB��Cd�D�Y���3����=q�;o�U�������S_ QP�{��:雏YuF�����5u�������NO|Lg?5֪h�V�67�6�p�7vPt\ך��=3�@�. W�%���؂*m�E��Λ�*���P
ʪP���`�
�
�qN�e�פ�<c�#�y4or���Gib�IZ\��[�X�-�Ĳ��,���������o�h8!��l}��)kzZ-��9��khk���O�	PA�\hC��1���3V�>1�����������w�kN��#�Fi��t�S9������/O(�jm��3o�x����=�v��QT|��϶?!m�2��IO~E�	�5ƛ��`�7�w�Y�g��i%2p8�Z��nsp��_<�fhB�VR�=�e�S�[��?�4����5�B�ݎ�'j�{��Z��x� ��'���2ɯ�N�2�g���]Π��`�q>#�Dg�,w�j�r�Hh�o�FG�ǟА�
��s�^��p`�J�:7��,�MT�r�M�e��Mg�~b�Z��}�Ŋ���4�����*e	����ӳ�5%������I�]g~�O���&�nڦ��c$Ռh���/�MX�}���s����U�=K�ܓ׌灋˂Y���c5�m�&RP3�t>�.�6$��Rh�m�c��w��4�d_#��A�	���[c���'z�ճY�f�pׅ��,�GP���Du�DGO�g���:��2�\���0n��_#ra�J-V����.��{��Ql����LAV牓G	I	>|96L�@V	q�;ܪK�m�42���L(xV(��Yr��m��� lQ&"Gʶ;
��?��@)��5�Y��me��lG��~z�{�G�F2U�n��A����Pd�k xkd��(Б��tx���]��~�>�����q���+.<y��fyl`,/��{�a��f~\�]��+j�����KO��͎3{�if�W_��~��/�3X�[{{b;(���<�G�uj��L|&:<Y9$��Iln^a���@,�ns5�����?�'���LG����^��Z-���\ʖ6Gl���N[���sT>���m�C�f��j�3k����x�+!ʷ��Y ���J:��r�0Fذ2�U%���/2i��::�R�=d��C�.s����hX�.����������oΜbH�]�P"�3�OOS�"�8��o#=.;],r��@�!Ƣ�H�UH�����Z��B�4���^��:���3X!�Yx��`��Hi+k=�r��)�dA%�oL,Y���w��@]�zڼ$�2e�1j0�����x�jG"��ڠ�\j�m�av���D�fGG<��_[���Q���Z̐65��¬Hu���2_�[p�T�S�7�3-��I�w�y5�o��y������@�5���y��*ooJ��U�Ie���"A<E�o�F=@]�'��o) �,�㙜p����Q;��t�X!H��ǉ�����\ȫ8��4��=U��<9ꈫ�+a�C��b�Ni�%��#��Ѱ�2�H�k� '~�k-Vu<*��*5`}M	*�8>~/�R�LG�R)�"���u5�͏���F>�����A����!�ȗ��G�0�H�.xH|��Tg�[�6��b�.Z/�uZ:@z~�S�����tE�/����AM"�au<,�wH�~��
#���CǈybQM��!Es�ᶖ0�3����U4��$U�������{��� ��C����M7 ��X,�K�nS�܄+� a��!���ƚ���,60M���w_���_��Y��cz=��~%)nx�Dա�l��n=Dt#o��q#� i�G��-�y	�T���G;����2�U4A��ШW�'�>yr�k��f�NҨ�O���s[M�������m�g��Dq�҄Տ�q��7�_G�ԃD��5d�A5�t���r��`.S�]Ͽ�S>PR�j�u����\���ۦ����5'����d�[KY&m�]GK#hZ!�[�s�g�jX�.�������������b�.{��=�!�> W��1�8�@��R�j�h%YY��2,f�C��C��՝-� D��m8k����t���>�0�;�TL�b���s��Փ-�7�&����r4+�y!3B{��M��%�駠}�ųGw��".��f[6/q�3!v�DW�+�����m�.�UA�?􎅽�dn����V|��)#�J0`&|���A��]ɚ��ظ�廳X��&E�%:�������	��ꏧniIp�D4���}]/�~}�5�3���,�ƾ�د�V���h5�,�Y�۫�f�^�,g���g�	z4'kT&�/]8~���u��O�k_
,���S1+���O�{����yC��8�xt��T��xV�	��5d�f+� �1�F�W���pD��q�N� ����́)��+�i/`�B����E�:����D���[j5����g��3@r�'��o��I�t57�.�ÎDeFY���uG/�zrC@{�da+x��=Լ��E:��/�X��w�Yɑe~x��K�b�ʥ�����*���ɣ~m���88��7�Y#��P�0��BF��^��8�~������M\lP%��W�@-<G|���̾���jw�E�w���+��Y��_�{�{q���ˎ��l{?��=Vj��2������-���z�]���%��n�����z�JJ���ᜎ�����D���gB�Om�f��s-��]=-����K�Y��h���Or��Ǝ�Z,2fJ�O�]�����Xbи�d�׎6���J�,{���}ח�Ŀ<M�8̘,V\��,�݀�ߞMY�\-�ag�'�{%ӳV��5���rbQU��j���i��MX�o��F�M�!��\m4I%����#c��H���z+����k�C�Pvi��~@�N,[	.9�U�1A��Bw��f���|M4*��3nc3��>��3����Ab���Ӡ�[F�t�������E��B�@tq�Sj��8x��DRDBD9����x�\�!��� �W��m�g�¨�~ٙ��:UH�~�n�|���$�>�U]� 8Ưd�l��)�Oו�JE��⪌��������C� ,�hD18ΐ��j�"����c���`v��J����ma˚�]R�������P>~�q{?/�7���r��vi���-�����&;[ړ�L���{��cu���ǌC�`p'a?�����g�������;�Ͽ��Re髷l�4Nو�X��,-����jl��=��0l����D�(7^��w6�I����{�%z��J�*�V��OɈ�/�wrX�^VƮ=��o�^ך/�L�r�S��B)���)*y��W�q$�l/�}&{�[@����z�%V��U#�6�hm�簅W [u�c�G��\N��_r���kz��2<dw�*�e'�q�%k�/9�b���������`���Ÿj�ib����m�����rS���'Pg �˨���xr9�u�v3_W���� ��bA�K��2>v9�H��5c���?�QG�ԫ����v�#�F)�kV󭔸>���M*��*�z��.���>G�t_�*ky�u���H�T��<�1GB^��H�y���}��Q����[v5׉;�`%x�ؙ<m���v3'�7Y�����_�e�m{��6(]�fJP�捊�iR:*�t��g�s�g{N@����5���&)K|a�'�M��HE���d�}�Ez��\��1����c��j�]S��!������>�1f@�%%����z��;��`zz�z�lQcM̛^�w\��D���~�l�8�o%�@0�n�Y_�6n>��mhD�t�z�.l�$ �`(.{%��)U�t)mF2��o���Ãs_���Y�Ð��Yw��3J䪂���ցd���Wm����׏��\�#Ս�h������s9��ݮ����ݴ�,�4�P_�C����m����!{�	��z@��:�+%�K1�RL�3T<�䷞��y'��u�p�8Ǉ&�^��O�O��xiu�1~h8f[�����3H��c �M�W��K?.���Zj��D���L�z��gd��q���y�h�j�qJÀTe!�|�����i�
Rf�N�t
1nPS���nfꀷ�r�8�G����h'���e�)}6�W$j}	��[ �Ç5wP��8���㜕<�w�詠k��,���7�=��y�����*
����l��c�� /�
�M96U�k.b��`�dQ=���)V�5�gUl<��^�F���=Za)�n�+)͔�h?F��<T�2 �!Fo@rw���4
�3��C�`��ƨ�?ap�zΜ�k�jljѳL�yx���v�Pf�����N�H� ��/֥i�������ԏAId5~�$���2j����C,b���;��>�?�����q2�������<�pqo
�X���Ɋ�#��*P��6�S�, W5u�(Ιl3�=��5�wc
w��L��V'���QQ)��hK>��֮ >�w��Mwn�
�3@�����q��q�*]9������4�k�{�O-�y/�G�+:�Y�ZD(=�a��i�'pmk�P���bB�6k�J\Bt��k�oGx�^=6!�G`dEĜ�E���-������\H��������8�N���h%���N��t��"�>�9�Ɖ9Ip��zp#f������3��n��&¯�P�!��$P�����x?�����ޠ�5���Π����������?�u�לc6f e*����儇_v��ٸP�YK˕���GgRW�w5l�>��·�M|��l��(М��e%yO����]\BY.�]�z���7Sc��ٓ'�f�:}�jw׮_�J���-om#5i�*Ė�N�>L��t��>D�9jY�R���bjzM��㷵'���=����L���g��V��H%����O�:Х��>�F/����Pk�f�
�^=!�)�w���Q/7w]_Ջ��}_�tD~o�6��e�bSb�OSNo��O����zj����Ē�e��M|��j'ܓ��5�E="�T5ʞ������=�Jr�Y�;����[���I��9���C �mi�T>�Si�y}�/�R& g�Z-}%[~F����m~�b��|B˷m+��4�*�\�q��+O2DA���ة&h0u6NR�{��+,��s�=�/J�[�t�F����=�ua�9`�l!Ro��y����݈X��f�5x���{p����&��RlA��F�c�#�\��
�|<Zʥ�}��ҹXn����7���_7Ou�a�6#al�d^��(���8/���ҵ	�5�Έ��8���5�L��;̦�Q����o���V����1JzL�zx�&0�ť�6�aa���C�#��<\��jG���^)h��}>*�����
��m���R����'(��g���2R�Zm��t��[��ֿ��Al����o�m��5�Ey���]��MC���� 5��G��u��N�����-Zݭ�v,�sA@ y��	��0I^O��g�vx�O{��p�s�pjM���A�
��1�G���ذ�_ٴl�C]�{qGF�(ag�
����8yt�|�'��[<$h��>����&}�sF�6��]����F9 ���7"�[j�w���U�E�_<�W��
K62�lɣ�@�w,�z[97 �������?i^�hBHKL��BD��N�s]�]�;�wR{��8+F�@h)M�-�\��4�-��v%�Z�Ҩ'zid�o_�83?D5���&����n����N�%Q�e��۔��@H+�C9ȫ
|���͒�U��Z)�3΃1�'>�f9�Wtf�Tz	$m�q��LZ�C<NF	g���h�&�sR�z<�$�s�4-�)���:Z�u����}�`����曒ݯH�k������Djl/���yos`Llw��#��R�Kѵ�Ո>�'�q��s` &�o����r�i�0@��*���s.
2_�%��n��O֭VVR�F�!Iy@�"�m�kjV,6S�G���P��j'R�� ht��U���ΞϏ��sn�H*%����A?zt��l �ރ�kv$%)���@H���LW.~�YV��iп� �5e	���8�>#�G�6sdX/����\[n�O_iS��#B���0��̀F~+��̭�|�u���A��/5ã��w�A%|�*�9���O���?�(f�Y��X��v�:Y��_�E��WO�]�������*2���z�`������ snN�M#;��(J<K��pDS�s5��ZW��<	WtJfW&sL�p,���sOree�D�h�}�:2����FE�W�ֹ2z���n�^B�3Z喖=�je��#�	�nΘڠ���UFS��J��ѻw��<-��͝�J$ �MzK��P�x@q��j��|�1�ܬ�'Vy)(^��=z������10�M#�c�i9m���J��-T�>��/t��t�=]����gD��,�򧙮����|��c]�u���@��S�瞵5�]�����Hv`5��j��h�N�2�P�����)+(�o�}5�|�!fP�N�<�q�RR<�G+�8�n)��O�TYQv�4���A�$z}|��xlmE�[�Gf��/4;�l�ύ���N���ʻ*����Iz��:�7U�PUZ��s�œWfT����'�kO��X�t 6�̫��
=��ڝqx���� �2�Q��Ҹ���5ۙ�B��!�m<Wj*4��K�D@����}y\��
U�g�$i��G^Mva�1��t /�u�M�zM\ q��	�_��8L��ʏ�8�����<�{��7[���"����#˩$ �l�q
�����'ʋ,����LP�ʳ]k/�:E4�k�u�|���U��2�Uݨ�Lo8��˥��x �0&�<�P�Rt���mfU4�׳�g|LM~�I�*9h�� �fA"%@�����>����,>�ZP}�܍ O�톽���
�ɞ��w*�1.���8��W�׊���-� �����t��C}ׇ_Q!�O��+6ˎ���̀78�}�%�:{d�r��jRb�G 2�,�mR*tlxY��2�Dk�+����潂y3o~4����Ti5PLC��X%��x���HpL���K͖ ֊c�u��U8�[t�"p�z�֒��<�
��[��#%7��͎�����P���}=os<c���p;f�f�wN%~���c;���N9�̬I^�(�X�d�[��Zm����$5a=�����G��偁k��h�F��s���j+R���!���1�ׇ���3�T�ż�F�Y�Z��^�+@_S! p���H\u8��bN�Vb:f�T��jc���#��_�(�3� m<K�|?߸�pf�%��G���ʖm_U	�^=b�̭�]2�R�f^�����nD�]g�{ZTBl�ԏ�=���M�d�`o��(/��v��d����!�-�݂،0�����������2]Bu1.&Ք�ǖj+���=�^�OO�6�}�^�{X3��"3��s1\O@9�H����k�� =��L��d�[V��U-4e��.��{"a�U�!�RJ�PS�iT�G�K}L�$�dn�l��YE�/�A�-�Ԡ�ط�L��\����1�e�}$��'SK���'S�yjc������|�zm���S%w�D
��5k�̀#���ɠ�7�n�O��
UǳL=to9�*v�&��g|:�027��[��g;��/�_S/لz��m��b���4���_�)�@�M�V�����RL���I��!�=��	t�x�/�_��P���nM� q��y<�P�wW(60��mKm�k�0�sã�kFT>���.W��cSY���=EQ� x�I�r����e���R���5?��q`l��ȵ�n����q�JuX��T�S�w<"��τ�Z�~ex琊jO/��,"ȒLg`���6��@c�` �/'���t�ݹڶ?բQ�ë��P�ށT������T�]YY�ܥ�$١��E(���:�cӝQY���C�������{�c��^�����~V������z]
�7��K�k���@��.���H��۴�C��":ǎ����Q!�����jҬw�~��s ��ot�.�:�.��[j��7\��܎�p7L�����:�? 'R�x/R����Rݕ���[�>�1����C�
)�;L�R^���+�����=�I��lzw����s���-��2��K9�8Vվs�hT����z�����>�
�2u02�;��w�|�k/�����2o����#�/c�G�L�6�h�:�D���'1 ����%���)/��<_ � ��0�>._�Ɲz�O�F�\�^�1.(�fV�Ր��V�pؼ��lg7�b�O�'vY���ޫ���}H^_�aMу�K;s_{A~=�}������?�3�wK�(�h\R��	&�1&��=��g�]}P���]PVy�f�����E9���4�S�O%����٩e�_�&��̫ϵ(�0���*��?=�u��e���E>�$~+E��oA���yB �u�?

����go7�v�N���	Q��,�r}1 rt�y������ �;
9�%:��8�15�=�>�$��"��~Wp��}�ܝ���W�	g�	@���x�����S�.�w�z?Z���{�E�5��`���u�d��F�r�I��av|�^�y !� L��cL��]y��RV�b��h�o��Y�=&����2����MB+MC6ǟ�z�MxI:̴߿�v��`��{�<ψ���?���0��
��6[���?���)س#���9ɼ\W���pPoղ���o����&>P���qQ�D���n��z�3��-I��c�2/�ʞ���%���?k�ﵫ�[�W��×��nC�wfe�I����N_��,Q��QbY#6�"����s�Y���t`#���*�N�-�����(�`\":� ���-����g��@�I����Xd��mA>ݛ�C�� &`a�N��"�La0�k�JR�"e@3�z���8��������{ۥ����U����Y$���ֿV�e%y����M��`��s��c��M����bΝ�1c�8OӨ!�o��=�t9�+���o{� �rg���Qw�����c�
<��lvǝ�3��ƀ��_<z����F���9]�B�7��_݌7��Y�lɀ��}#F6uB^�p�ޡ��k,��M���c��CW�v��=���Eʖ���u\���з1���Ą�e�pb�Z�	Xjc�;,
n��Pޥ���VǅәvQ�yݢ0<Z�M�U�@/��v,��7B�a�d�F@r��{��Z�2��f���?H���I-����YxW��5�*r�⸉����Z��Ԥ����=@�����>L���i�U�8�s���j�FW�&}�]����� �I?�
&��'#o0���u��!�K&8����)�y
��~a+D1��c�ɕ&L�o�I�4�Y��?�uI2���pպ�������)���gg �����6�8=`A��%���j���8����Q��r��m*X��WS�6ʊ־��2�E�4��!�{���怟�#s�k�K�JRNJ�>��`o��|�w(�&�+�?ʓ�gTN~r�KP[
-W��6�rfT�g��"q�z�*/�k�'BW� �����5bfT������#�ɪ�Bo<�6Ad��%�fv��vl׮��P�$t�����냤���Ñ�N xs��D��^ό4�=܍$��m���m���mN7"\}9B������6�F���^�2Ň)��=�3�J�qs��L�ՈW�,�I	��rK����k�����Sr�6~��ki�K�aj�)� )�O���\�L��|�ps"�����n�����ZX���f
;��7HW^sx�;zb�i�+&=��3�=4%�����e3ҦO�۷�<w>2a�"z\��{P(��f�S�H��YԄ@�d��Oxt�C��%�I�f�~�JP��VLM���#<���4"/�R�z!}�!'A��)6Q'���s����YJ� ���:�ݫ�A�s��`�-l�#,jc��%��b�G���L�� z|���f-Wb��8�iO0�
S���4�?�R"���/��ʮـi��^-��>��MB�j���gApL$^{��?��ln�;�}���X���4����^��p�h�4f\�L���$Hp�~����騛��(�q�Bmǭ�z��Z���C���P�B�.��{���B����R��%���fO���']n��g�U��4�Z�p�5��N��/w��Up ��z&�U����nCyc(�$��g9W����G�{�������;࢝q6�'�3�n�ìAd�>=H)�:.ۏ}Ks
�N���qK�u�+�-�"��۩�_��'���6���6��Ƶ7��4X I�/_9���+��0+���ejql�hsd����l��ݍUwS*�ސOc�i�_��hg��1�~|�E���H�|,k��Ĺ��VBwK����FB<�f���jd���|!�a��-PZA���sa�D��"�SBHN�ﻙǍ��~��8��OcNri�J�A��)��*T �$46�j��U>cu�P_�l7��YQ#���BN@��en���+.�uE�BS�E�E��D��M��k�����ӯ�U\a u�+n��/,d
+8�i|3����\l�w;�{��*��GV%���+�.g�B���b�I�olnpE{�� eʝ�]���W�w����[����!����!�Ғ�'Ѷa�	�4��<+2di�&�7�X��+��{�տw�J����֭!{���E�R�L�����9������z�о��>D�[Z|�X-K�;r�Rϴ����0g�g����6���i`1h['��,�G-�2�e#^�ְ����[���aL^��[h��Z�?i
}�a��Xv��kz��
ĀV�%��#��G���%����.�g�Ɇ|����P���g���}��݀iL}u��m[�`��H�B�z���n��v���� ;S:���C/D�/JX,���2f��)��9~�k�:���.��0^��~�2⡤�T	yI����?�FE��M�r��D����uc���r1#rN5q�B|�C;���|��C��i7Z����c*6v�T��w��wyG�Z6SY��}�#p��s3��`�5i)���Tx�������%_�e������3���r��������c=��!���x��_��2��m���P6����U�K�H���^�r�hk-�d�}D�����bq��þ$F��Jk��75"<����n�)!2����o_���6W.�z�vyV���%(҅��[����-���:��L�V�b()a�$-���up��oE�F[�n�k\\|�{Z����,hi�vd�d 4�N�tݮ�����u�v�x~� �hI;�~�ԣ/=�m^��1V�&qPc[Ϋp�-{zSj5���K��{�}�)��f��Du�L�,��]���n�,���`��;3�GO����`��;5V�����ln'%V��h�_?��&rh�R��:�]�����'Y��v4oR!�vǨA��sBh*�ƞC���\�ʿL���hp�^����)H����U�� ��=�<&M�v�_����8|o�pX,+���҄����,�r�WP��Ev��R���-��0�5|*�{��:�=���`Ux -s�����P�a4�fxز�G�G��4�Qa����9��'���HP��{G4���}�H���^;4��������h�2�i �|�H^�Y��r'{RZ����ɜ���yx>u�VD�
 *YǳomA>A�	R��g����P��x��W-v�[l͋�͕�q|�:�9�?��?�-X�?U��C*�a��T��N�:9��M��f-�q�@��韈�81�m%��
�K�1�7��z�+w�G<�3"J8C3Y��@�U�؇?��Ѓ۔�P��Y�[�&7���Go�yZT��]%�g�?Xw�w�2234)'�ΝU� ��b����gC��o�ϼ��z�k4j�G���ĥ�:�����i�z~ކǺ=8$�,�@�N�����Fj�w��$~l�VG�Vp���*����ej,��^�e5�k����g��8ۯ�."í�	�k"���_`��W�a�l4����d���~�8��ʣ�&f.��>�����
�ވU'�Ӻ�R�r5n4-vhf��G�,�������ЄC��h/r����ݲx)V�X+ɭO��®�T��x�p�@l�����=F*E_w7CEK$�H;`�5���!)�K�U�}j�Ǻ9[���*[��6#��a۫�AJ��h um
��e���]�'I$��O�P���o��3��q���e �
+Wǘs�Q��߼1�L]ݑ9Ԙ�$���+���WC��2c���ͥ�]�.Jk�{���EBR��Q1vL���T5�ӆ�8����g��?�X�����������X���8�6D$��ɒjQi:+
���Y�KO�];��F�����}N�Զ�p�s��x�9Ah�w���w]NU�l\���)�*��?����Z�=������Ig�﫟	[���@su�CF�. 2�2�c�C�&���@���ծ�Tp]t��al�<�?mҘ0���A��]��<@Õ@�,�M�T�:wh���P���
(37{!��M����l�1����u*���T�o�xF�\��\��b�b78���R�Q���c����;K��Z=ɖ��$��e�Ԫ� 姺쭝y������g������!�jO�Zmb���sd�o��-c�q����K����'^��0�sI���G0xÏ?�2.w^��+���:�\�v�g�W-@�<X���,ÃÈ/ˈ;�Fai8��s��1�m�0�E%D_�b��C(@� 4�HK�+�3&4������B�* %٬�:�lJ�?��Q�����p���Ѫs8�ׯ��{����S)�=�]�̮�'�B�+-��?'-@���s����v]�Y��3B<�_�j6�g6�L=8�
d�t
B�Gޔ�S�-a�J�� ͒&vv����I��0.��Vo��]�D�82������!mg�����+�=��ly��T����B:��eKl�,�-+�K�Gc�^}�t(̈́k���M�q[gש�u([�Kv{����8&���s�y��< �(�1� V
���W�N�����g����H�%3� U�"`�g7,5Z�xlV��Ց��ͪB�
ڢ~ێ.{��50�Z�l�ŕ$>��Z8@5�,���&ٓ���sX���$�D��ō�H�C�nva1q�/z��O��y
�[Nu?�W�Es�ΰT�]V��o�_B?�6_�A�1v���J�h���ƿ��Q9R��:8ד�э�h t;��8�l��\����3��vl�Ƿ�	]����;A��D���q��s����dcݽm%ԐZ�gYN��k����#�=����|�ŵ�
���O_����ڟ�\���JI�����Θo�c��w�˕�*�#�}�����Th���r�O��-�@'%6�
&�K��o�pn_�f��:��?9�oc�����<v+8�E` ��^Zz�ȸRh�~�� Ԉ�������v�<� ,�GyG?K7	)�ѻ�O���uȶ��Ӕ�����U�0b���M��L�+�ƁA���kV;�J�g���ߧv�����E���~�&�	�PT��y�����h�з�fhg�C
	�[嵢�B&�g".j�QHo���A�{�ʹH�����
��ۥ� ��������+�UZ������0��,�&�ρ�aL��<�N��f�~�*����Y�M��W�b݅FE@zN��ތC7iNsK$�-֙�0�����jo'Pm��NBj.>������_SC�vP>��R���ǆN���Vj���7%��H�O:yW?��`�|�.����T{V�1�~�b~
��wa�0����9r���g���D��=�"�l�����\�����o��al��_q��fȯ9�F����I����o�PZ9���?wl�e��e(kw��v}��ؼ:gn%��iɨ���a����il��̧�o}�<�<�t_�(��A@������9�K����*/�����b9�<i;��;��'����i}�(l���̩v�և�J8`�Dfc�h�����ꏓn�UlJ��/'?��	�Q9�QU����~��S랠��z�|�-�p_n3�6&��a9S7���l���~����?�`cZ�`��o����>o����\���ѽ�����yCl�
(��ˢrq��}�������;���Zfɼ�]�:�`����²ژ�_��,�@�4�e�����a�uVH"&âfl���RN�{}��q��6���H��E���3>��C�'ݼ�6��cs�W�i��lZ����t�F����0��:8���;i[�;:�oµ�wٮ��3~|���]�ZW�K���!�r�,�	�Bګ�Ġ�^���Gu���V�E,��s����`c�����"���ؾR����r�r���`{H,{�z�����a��q��AۀN���Y��:��$8�&|�~����Nw�͓�gX�g�׮~ϴ_����|�g��R1�Q�	{���w�����e�@T���<���t�]t�����hu�d�8�A�I>'\ @�4s��W4�>��{�iK�ci�G��\���T�W�U9Fߥv��3_6@��~=h`���h��PuX+�����"�4^O�ߕFK�w�"�*)����Ӹ8�����\v��l��k�&�[B�����۹8:L��o@J0R���aƩ�l����83'��6 � ����	��,{&�Z�W��TY3j�.,<p'e�'� k���|���r��'��/M9��pɛ���,���A�&Q.�2����3�hg��j�m�I�V=���t�\��E:�M�%�n]�S�е�.=h�l�<&����\2���j}�p��?4��>���$��>�DVIs��o;{&��]�,kbZ�Ǹ�V�b�{���i�N�]�=�a?Cc�J�k{������֘̐Wj2]?�m��][��t(ЪĻ��E	�uNq�p���D�CY/@H��c����v`L��z���>��y,���+�^�dP�h����	ԓ׭@`�Rd���$��؈K���`�v1?�*�c�����[�{��� ��P)�zx�=]&�*�Ze�	��v8kJ�H��V���Y!��Clܛ���.g�;¨�eTo����,�=G:���XK�!®����s�U2�r�d�-�
f�a����<�3L�C� �Cc��>�бس,-���V�Z�������3	����{�jl:�D���VΫ�(�_
�85őc��r! :��k�I�5h��+;�H J}c���<�������8UhS�
Ģ*�U@D��y'�8s�c_�}�L~էn����Q���ߨ���z���^",�n>�To�B��ͲvJD��ݫ�% �o/�=T?�Ϡy�*:w'��l|3�_�[�g�:rX���`V"��l*���3�X���ۯ@Vk^ĳ��~b��4ھ@Gn��8�]/�6w}"��ԟ�ʩ���'<]Ӎ�l�8l9=��;Fc=�2w j�~u
��,H�B6�����K_ʩ���Xc'=_�@Dxp"Pi���܉��ˎ{��K��b�.�"���������n,�h��o�Eъ�� ��vMi+�1ʟ	���9��~��ȉ�5�I=;�;L���L&�~'���UcMѓ�H͜{w+��E�$���G�t��l����06�a��:�3`�����Ʈ�40������a4_���Z I�(�A6ZƑ��1�/��0�ИƔ��|��_w�n�d1�0I�E��hcS��ׅ|-�ʟYeE/�P�Y�M9��C��3�=���>������e�����x��-�dc��'T��Z��Րx\=��d9"���z�Y�;�R��Q�,GD��^Q9׀i;D�Qt�0�5�F�#����W��Y���W��R8���){\����S�z��K�z�
i�.F0���V�����n��x�I��As)��߫��7[26�?%�6g!���Y�A�D�OL�Fb�Yuy�2 F�
m-s1�����/�;�w��$sX�VOU�q�8�g���>L����ż4�II:L��c}kܻ��I��+S��藿��S�.D����md�lGf��>]0?�Rsl����L�T`a9!?���AװY��x�%j�A
s��:��g'&�'��2�s<�������讎��<@Xeھj��\:A�P^n\ނ�ݘ����D,Ml���{�������z���n�����B���ZB���9"lsh;#]�~��������^Ċ"/R^m_pQ<�C�wȏ�[c��5�[����������DDJ՟�3y���=r�h'PG^nx_��������/BǥA��M��b�t#�� �%}���6�E�����V��n`�'���:��K<����;�E���d�h��<��eX�*Y3��G/���mB��h��`5�U�h�D(p邕(���O}�C��T�jfɊ��ү+�I}���D�C�ޣ�`�j1l��U�	"�� 
�=O�QH��eѫ�`֥$9s�z5��VuE~��%�-n�խ������wȁ%����c�+_qAt��o� �m����"9�v`�<@
����!�hR4��H��qIz����0�g���6��%��?�wf�߄��Ӻ�=� ��� A��ů�I佚�&���˂,��.n�V��`�j,��h��m�����k+΋��%�.�ZJ�
v�x��q]�E&KBB��]S��4���
7�:n��ߣ����;��VSAY!�B/wTx���$[��:1k��Ł�DU���SX,��o�_|�j�/�T�6վ�p<���B��y��c�Y��~����uL|��;YХYy�Xn�T!2Lf����.���K����f�V|�s�A�[�B��L�x�4��t�dX������Z���4�%W����w� �f���<�O�o9Ԏ̟�5e�x@붼�>���=A�e\�h�pV��)`*�0�o�F��b�B���t��8C}v6n����=�?�{6���^��I`��ͪ��tM���",V��c����wY 0u��|+|��ց,�A�y�u����zkͫ=oU��5]//VWQ8�`)V��a[?���8�k&%F}�����!�l���㥎ڽ��7����I����P���Й�Θ�2=��"'g��Jkw,۫]��&CH)Q[�A���m���{��^�����C^���}ݵ��P`Vl��Wn�y�d,��L����������T�0�����_#��Ǟ�,�%`1�pU�T�YRآjO���� h���?(Y�������yc�\��YX4}����/>�^p��j��r����7^~nw���:��; ���V�,�0�@.#��|�ݐ�013X)]PY-ړ��xs�<���ݸ3z>^,hdz\-�o32��Ǖl�*���!<2�������F7�1m�F���]st���F�^�%-)��$�Lԥ��jQ9�I�ݙ{b���6gD�R��设$wӠ�b��X"��}5�g�W�fk-�V�#3�O1����L�ح�xz$Č\�]��b��BK �K��m�0�w�q� � ��O��*&�4\?Z7���y�����<�\8�g�n�w
U��V����r)�r��P[�=�14����
=�h9����G9�4Ϻ�`���r�Q�BQj�_��L�eٔhV9?��{ �0YU�n*��t:Q=�o��g���lDu��L���k�����<�ߒ�7�/���6p?�U��f4���`Ajʼ�X�]����?`d5��g9<�����7���y5�UI�{-��|R,Ψ�8����GJ]6����9�2�I���``�v�ی^ο�6a1{/���&��oB����LG�\͜�k��m'+Jp���v������Y/��c�k�k�'
[�F$��+:��p:4�@l�ޖ	�Լ�tt1`�ް�p?�q�/����f������,�t����Hv�-y��yJ��e7��թ�� �ɓ^�)����E$���]�����Q.�p�Rڷ�y��r�j����� Q8*'⻲s��7T���ZMM�dms��ԥ���$ș���q7(l��w�.�@���׻�`����D�[4xL�h��]L�У��{�F���u�w���H���u�����u��S�붿r
c"��o���$���a��鬱�u���`�˃1��M��f ���G�ۋ��B�"�C�|�+�qs��+k��ͼ܌x߂�w��
�ˤ�N:�(�zx�������iwW?.Z���]T�r�dx4\�����u���mz�]���ٙ����Q�BC�����?K��~��y^;��Z~:b��s��O.��d�ܾ�x��߯��{N�<m�6@2�AH� �=�y=���Oo���Dk,
N̐�:��}d�y�t�`�v�8��M�<�$�,[>����Ҥͭ�FV���$}�'~\�����ӊ�i������X�F����m�tؼ��IÇ����0�҇s_��9�4���q��]U�}J6qte�;�E�`sa��i7�mYp}S ޠH挺R�����I$��G�?>���1��D&��Ct����{W�^��ZF�Xۏ�hh:I�2��T.���tp �;ʸ$;n7��C�.��fֳJ)lBy�P8�\5s�"*'�Z.��_��A$��]��bm[L"Wv�t;�vu���L�������Qb�Ʌ�{�:���^��21��0� ��y#MD�}�e��ٚ� N����l�к?�����T�E���P�]L/8�:4z����l�l�Ʉ����((���͉��I���:5�>%�X�`3�>�.�%i����_O�K-�11���������{�3��Y#*�Ի��\j9�z�fWg�Q�7���U&�[�Y
*Hy-~��so�s��χ!]�2�z�>����I�s2�,��g�qÂl�o��F�>����8�=�aa���q5!��Q�����8���f�?�VA)X�闓}/{V���&�j��{mj��'a�U.N�����2���i�h��WSm؛A��i���J����7FN�@���
&}��w��w䊔#��:W1���=rNc�5�}`�G�f͞eR3�0_��ED�3_���������@D�T��퇫e�Tq���`�{�����A>�v=��k��ށ��Zf�VH8��B>6���ں���/���Q���ݡVy���=�[yS<�D�ZP� <{�-Y�/����d?j1�X��j�k���TL�s@|�m}qq�� ���j�Xg/��PHr�WƷַ�2;�鹖�=`���%r+�-ez�m"P54x*P� �QÏ������U�g�� ��+H�w�]u�B�:4�ٯ�ǟ6n<���5rRR��R7��J�c�XS�%%�'ٸ9�7���,/�)c�f���$$( �l��n]"�=o:úH��`L[>TY���C|���&���OԘ��RZu����"J�n�F�ÿ7�`��CA�<���]a�]\�9tԄ+>�|�`�pfc��	]��A:zǉ$2v8v/��k/l�p�'�D�?�lR|_8�_������P7�o��| ���	�����z���zdaK�DS ��W�u0�H�=wr28g̡�8Xj��+	�nT-4D���8v���E�,"8*X�	�9��}��t~\4d����2��Phrw�V�}#�g��ſ�.�us��f��o>򀿡���\\�&�R��b�����8��%n��kA�F�ZO_���7�FJ�v�h��[O]X��\��3(��O�o���eP��8J�����'�~�*.�{����� �$Q$��[�\?�e�zS�VK�w
��YV��؎��rYc8����Ԃ���?gʢg�|e��4���ER�m1�Ѭ���W{����8 a�.d1L�1�
��I ��3�MF�I8a��6%!<~ӄ*�&��l���ģ�n��U��M��j>��q��d�!��~���O�6�����1f"�oɁ=��ɴ�`Nda{���V��8ũUE~���s�X6ݹ=�4�m�����I�c��&:�
KwuՒKj�=`����j]��n�N�' 3YubyǼߘUm��$��`
Z��ɏ���K�G��,��U�`$�C�6Rk�eH��Q��<7��E�oz�qN���5l���3�6�����ډ�,-)��A��������'e�D���|M � ��a����VSs�A����>�N֖�/���'R6�FO�~��Ǽgy`��U���>��@�g�oz1� �q��a<9�a�v'|����GOXPܝ�Q����@��1�IΜ��c����
���cNڟ��;+	褄�MJn�3Y�2����r~�������+�R��>��`��{�	!��˸~�Z;ڭ]�	����<RZJ~�� .Y�!�=B-+h��x��֎W�J�b�168������n@�4ܨ�����N�3��7g��Dө���O�&��/X������.�
�E���ї�o���?�ү�0| ��l��ݜg@�{� �4/_���Z�0�J*ϳ�/���>�1��r:��[Pk~E���Nɸ��Ԑ�G4J6MU5��WC�\�ω���U~	��2�֟��J^%����ШT�?ljaѠ�w ��N\�E���6۴��OJvl�Cm���iҢ��W��
ɛZ��IRh۶��֟nTn��5�� �1�	b�|�kq����{��w����L�������|�.���_��4������Q�;�
�k>�[n��k�� d�-��>~�^�z�2��gƇ���UH�RR+_�b�ڇ0j�6@Qv�q�-�c�����#���8��[UĆ�
`귂!s�#S`#���[�Rn��_S��+�H��v�#b!w����o׾#�gt�������]����-7s������@��T}�,��bzI�G����ו[z�� s�U�ˇ��P2�5�Vs�hW����e�>8��c*�bci7�sgG�]m2C.��bi�U����ԔP��ɺ��Ŝ�]��+���K��5����9�����I���.�r�/f�1iǣ�i0O�i�+�ce���.z~�c��U��>��wZ!�ܑL�|�w����x8yb`u�r��a��}`D��p�%L�2Њ�ˋ�sj�����(��iñy�б�9��~�u�/� #��%WE2i��j�w�/}��"�*_�p��J�n��
�1�>k!@�v�(���>�a��&�;�wQa;����O�'u��
D��M�i|L�ꤗk��CL���t�& �;�$��� ㈖6W�i/�i��({G�]Z0�����_��v5v7Se{��bu#���r�[�%o��t�~��M�<��9���w�cb��g�W}�ϤYw\��i3�&���=0:����6���}'���bC���l�g��V�\�?�qC�r����S������ݘ=L�]�y�-y}n���_Y:���RQ���
F2����8�8~:g�i��r��A����ǧ,-'�f�Bh��I��=���k��[`�~�|H6��G7cFj� ����c�%dq��#Xc��.�=������_ ���� �zm<�9�n����,�N6����S�Nu���KKzv�J2���Ĝ�{��Ts4:3�),L������O���/�����aj�o2�9"���^������>����H��#�R+��]�i5a�k�b�����Q�Q�݆@mw-h���w��r��ӟ~���U3�0�e��<~_tO�{ C�~�_)�� 3o �R�G5�јN$�?/p /E�Y3-kC~��8���1d�l�xܠ:��_�}̧s ��c5�hIH���;�P8�j���y��Q������9��J3�����P��b����pS��%��Bv�'yo����  u�G��=uP%X�����#��Ƽ<N3JZ]��V#�@Ka7�����'��z\C���0��� M�޷�m��)$��DaϺ# V�';	  |������DJ�JI@��/&��o�j��j�T,��K���xƄ��?���|h���s��ˮ��K����7�T�Q1��P�VqP��+A	���n������V�@�U������If>��J���a���a��x�u~�w}�@�u���ԣ{xg�����t�_\�U�������%r���sTGc]M�7A6�u���c��.ԞcQ$uu���:Cmc�ʼxh���vM�su���p��`E*}3�Ak[hV�_�d�����&u�V����]�ov�?@�3d��W�n� �
(�5�̖�u�F�L�>�u�)�}���@۾�v?(P{?@Lv�)�i���Nw�0�;���$Z��U�ǜG��cO�`�����YK˨�{`�J��������:d���?���xG;�dP�����]�\�������oz-�h�#�{�)�B:ߥ�V�KO^�@g,�t���?�����/A�A�Vjb�'3�����t	��R�1�����c(�9?�.?���Zކ�'�{U�S������^�
�5��l4��U� T�ĺ5l��Q���[�]���2D�nyW<A3��J^��_17rf�O_���@����,�Ժ���D���XۖŦ8v*�hA��(���S��ʾrrէ���j�Ő�=�wqi��G�5����f(n}��ܕ
�t�[�P<xk�e����TY�b��eT��'�X
?_#�}ua�vWG���;0InYhǡ���Q�O#��{%���� �K-�@3���x%�m+�����Ղ�YbY6c�h���Rlً�JΥ�Q#a-W�1Xb����6�@�S:/7@�z��d��Q.;��I/�<������iW�W���e�! 1�j�H ���ᗡ{�'�nU >�ҐHLf-F��2��C
����]��3�Qs�C�c�n ���s�h�nw��*� i��IIYa9Ǜ�����8�}����Qwմ�Y[����N�T�ǔl��^4�os*8j{I�i6y�f�J�2�>c����%�Y!��������~z� ���5W�Z��{�jg�B�M�c\�N��!��qd�@��*�ul�����% �\��9�d�u;LS���4�J�o��L�6X��I��֒�t	K�ޚ����v��pnlO�:���$�}<��X��ٳ����^��#�Vb��W[�v���`fά��ث�8��4�B	��e-�u_�&�a��Nc�V�"��8��w��0�&�����I�;}I��a�J��1}=����]*��p�n����o��i���7)CŠ�U�bM`�� ����#���������q5ѡ:_F��,��z��O� 8{v�WO�qs���W�̆�����k3�>�GG��_��i���j !X<���9��A������d�δHY:J%,nU��cYk#(8殳kI�v. Ps�G,�N40�� �$���|�,B��������P�<-��lC����������?�J��;����}��u�l��%-������w%3�Y~cӆVXMA��e�Nw�zL�n]���{��O�6[�M:�Id*�v����)��Hvq���cz��e�֏�� D�ų�ߡ�+fS��(�
��%]&@]�����,�m�0�;r����+Y��{��ƃ��ONȿn�jo,�d���?��󂩕Udz�"�"r��9LW�$U�A�+�����ٌ�:���ߡ�8q1��:���%�R���=qӐ�0e�k�a4�l���[��솮�Fk(oU(���~�w��;���x��?�Au�Y����%�ٴ��Xzz���#�a:��û|h�"=���e���d���W�°�Լx�0�}LG�$��P.(Z����D�'T{�o�ܣ���܀g*��RP�5�2֗L���;��)�Y���ӊ�8b�RF�}���J0��	��h��[啨�Ͻ�{��Eq��3����h`wd��_���@꬟a�����d_]�$����n�n��ƙ�?M���=�L��|�H�٠WZ����Le��B\�*�m9>�*]q�J:�nl�D1�%C.ۘO���D@�k��\����jA^(U��� z���h����W�eY͜���/�f&߽��޼.^U&Ņ� OQ���T]���Q��2-Yj�Ļ�RW�WVe�&��������V�)t"�U�V��W�|-�FzZ���lV����}�3P��]���<����ס
���ր���&^/�R؋;J4�q��>���1�-tU9��y-͟f��B�
�Tv��V�z�/�K 0b'�������F�ҟl��6f�SA�F�� ����(7���s9��̀'Y坯BY�;^f�'#j����	۩�������*_cƋ��5�[�9jM����6t���-���F��1��`ʞ]I��/@�ٚ*��xKdSu�2=}��s,���_j��2,�:���Z����L�N�Џ�P�^m�mڍ�x�1�/]�4l��̍�zh�=�,�Ad���&�w�ܒu�������Eh��t]���Ը�__��3)g툷�1bU܋��G���0��<$i�ao�� ;��$�ۧeX�~Śf_����?(n/�(t�1BȲ�fu�6}��Tc�=��- N��?վ簯koi��y��HQ�4��a�j�y�c�t�X~�ϕ3��B��Fc�%��%�R�y`(��s6��g�"�Ƣ��VN�%��!D�GMpgک��uv�UQ���߄4JYՉ�'���Q 1�����F�ۀID��??��y�ެ|'��� 7F���V0�Sl,}G�mrb��$�u��>i˂�^Y��6�{����0�8��O(��Yd(9�����N>S��m��!,)��Y���k]�E!������{iC�l��l�2U��+�,L���vv�����S��%�*}ߍ6�s��PL�w�x��IC@��8�tx����sڹ��<��ޖ�����,Z���Le��ܲ�V��S7
�<./9�_K@MSb;Y3�F�F�[d�@��9�Y�ᗁL��&ƨ��͗7C����S�����7<ng�\p͉����ۢ͒��s�`�\^��%&�=ޗT��&�ip(�ߜ��a��%�kw��cҎ�e\�8��l���s��e�Ia7��tJ^������wIEъ��I��Z��~���6neH�B0��嫹6�tޏrrf�[�A�-_M>�M� $b��O��Mr\{8)��3�@��{��ʐA���Ŋ�?t���xz}��6� �|-����m"��NqT�:w})����\��-�c�7���=^�ZS5K9�]�X{����e����$��g�i�u]�Q󳞁�I�>zҧ��vh������qQ$��𸸀Jr Q�]�$Q�� �"� 9���s�AQPI*9�䌒3��"Ir�4�0�a~U=��|�������Uu�9�[��7� ׼���嘪�Pg%�����\��m����n�-�{���/�������"N����S�����,�ŉ��J�D��Q��`�E��@9�Ԑi��A-�$r�O���te��j��dEհ;�&Eu�5ܕ�ӏ4=�G(��(�+�cx���b
��y޿/�5Y������-�ݻ{Ms͑,X���O�p��?Ű���&����T+����s'	��wq�t�Ě�6C��0��N�2i����)�O��p��1��$��JE7g�mѲ����GqVI���Be=(��������-�k3`ť��Ӌ�7'�����*��J��\�K�9*������W:�R��O#]TvJ9��n�+ˀ�D�B���g��K'�nE�<2&U���h�J����DM}jsŃ��m�R(� R���Toh�����^F�s�;A�b3�n_Z@��
�&R��NͩX�tpM%��S��DP�V�zp�k��B����C@�M]~�X\������p����ƙU��ߚ��\T�g+W�x�����#��Ovg?��_�r���?bǕhjy��SE�?�#Ҿ��ʞ����q�������fU<���y?ٹ��#����YO�럊ˬ��!�wh:cgy�V�;�c��:?�R��n�!�e��l�Ad<�0ǃ�<��Q��*�7�jno��
�T�Avd��������>���X��rr�ZN�0��xF��u2���L��{�3�U�5��kBEsobBf�3gC6�s$@�8��&�Y!/���'G���O��WGG `���[x$^����*�����E���E����)�M��Ծ�ۼ3��@g��l����Q��!�:zb�B! ��%��!���tw'Qe�!]j�Z�"��*|��'��:U91mC�zu�e=h���1�<Ms����˟QF��]oDX�R�Cޥ�e�����$2V~���x5j���<#7s�UÚMT��T+���)6���5X�:(H�ฎ��*7���!ۏTn�*�{��p���������D
!oр^�:s�/��a�P.L�j�uX����ޗ��w���_��C�w_�n^��Y��	����%�r��х��@�6l���(�T�,�R�h�y@�}���g�.B���'�ծF���%k������xo<��O-�ziP��:������z��ӝOa�"�^To�*RNqd}烮��nX<`}�O��3k���QJyp���ȇ�S�&z�X���d(����wǚ^�@CD���6t���$nӛ{89�w��acz�:zN�X��s�|� �v�1�,$9�dY��k���0�O���Q-<9��qw�X�R<E�$�h�W6ܮ��|e��ˑ��ٔ�瀼t��J�2GL�-��T�	���ʭ�$�+e�*u5;��R�7��vܕOfwd�������:$l���Kc%h�+�@G��]���1�����cp� K�	��K>>'3?U��YleS���Q7��a��ٵPk�Y��^4�/�B�{Ng����;�����q�MSٱ6b��1u��f��m��Dt���f��;!�x-i���ܽx�}���g�'�6'z�)�_/�4z�	~��2�i���`wP�r��BY;G�v=���3FO��7�D����&�g�R?��j�|_B��@AN�0��xP��Ձ����β�d�$�5�{#Z�n*Q�cԯO��8i���ʍ@n�p��[\��'>l5�ӥM��,
8��b�Sӛ"@cd�^�8���|�H��#�RLfn����5%�^�v�]ﾏ�2���N��[si��^��J�@|�wծ{5�BƨREm-�^A�R,v��_
�GNS�������8��_�v�&��-OM/z��w������o��A��Jޯ��P���G��/�X.dZ����ֶYD1��τ3;	nP.E�d͵���@������v#�=K��e�(���nފ�A�ɹ�z�y[^�H��gs���|�+���z�[ӣ;��d���7��]�I���a[�S�7�R��a��H��'�)�����N��[��tu���.�vegg"����!���O�Z*I�zގs��`p
ܡUv�J6",��κW=�6�c&��p�����Ҫ,첥���m��9�NVҸJ��� r��.Zx��!�����{8x�Wu��PQ��%/`�VV�%��"T��N�'�7ÌR[n�|������~
�{uS)�vU�y��Kp�8�b	[L�vp��A��X/����	9�m��i�Z����\�L��t�����ˡ�"z{O�ijp����.E���(T �,y'���rv@|���a'/�Gߏ8Qc�	{g��n������̎�*/v���Ce����$l(O�~��<�O����x�Su�
V��)�+���������� �JN�ɖ~�6�B��5�G���8�!yC�f��SQ�h(Z�T����-;�j9��7�l{3����*�Ϯ�>�q�ZB^�AQ��l���	L���ލ�ao��H�!oB�Y�t�JhoV����넕��q��ZbHk`H����09���~hz�d����$�>}��k�"�W2�> ��M�2�6L���qǤe��G�6=�y��}{Z1ٵ1��b����Ĳy>���쐓���wqq����f����c,!C��5�.��e-������<�+Y��dl�^z��892��KiE���6@g���Wfm*/X�H;�����
 �3�'�;�C6�������If����Ip�R����fa�ލ�����s�#�
�I��(�Xi�����_�eQ��"���ٍ�Y4�"�{�$�����3t5e���l�ӄ�dB�r��'|>�2܇��tZO����vUR*��I���͛� ���M�uq[$�yQ����k?x̋���bzGdA|�16Eԉ�M��3iQ����� ��_�硛]L����ʙu��B�ԟ[���]�����_�%ZI�U&|p]�b����<ؿ�3t��!�}��-�&��_�lǻ�:�.���RN�+���H��U��$Nu<���n	]M"xo������F��g-�������.�/l`�k9�ްz
��|3�9@�ft��r,"g�����w-�(�\d��|�hz����o������HU��T����[�u�i0��-;��p)�ߦ,������{K:��)^fh;7�>pTLE�a��>cR����>jԙ+�O��5XK�q`&�����9����?�^Y�8t���e���v��Cр������x�\�Ârl��G�H��C7��{�})A�y�Nթ�`S�ޭc���ǧ�V�;�3Ww��g��IH�P��/U���?��pNNn�m��+`:��芋��(�|�qʄ*�TS&$c��l�-6����2�>��vܪ��E|�`ٜ���i�2t�g��=|_CFT��7����F����l��c�/���|�O�����r*d���@�~��
dԍ�����h���̬���t�����3@�z�g�1�7�d�&�"o	Q�����v�=T����]U&�CMG)n��͆g���,����k@л,���M҇§ʍ ��+��o�L"�3������5 ���mn���!k�Ec�v�fV�4���/3�J7S7�~X�]h���?�Zj���Ju�n�:�R�6)��/'�mʲe��8��R�5�����O��U�%Z����~�RMW[�k�����n
ɝ���P�i��k��'Y��B������h�2���vhZ!�9�`lcq��9v�Z�V���~{����F͛k���8|�0��]��H*f��W���4t�+��	�;7I�{ER��ꛗ�R5���&-�����e�~ys�ڭ��P�U��M�e�I��V���}I�N�ѱ�KT�7j�Tc�%�w&:�ʨ!��8�#%:�����E<���_i�\8|-�@q7/v �$K�sI*3�?��2k�iP�T�m�BXO�njj|�-�?�z��.�7��Wa�i�so�u�n��@���`o��!9� Kl�=��ul/5吾���}��`v�^OK�ow$�ߕ�%�1qϛ���8��/_�7��7�^�L��x��΅{��zɖ�O�7�P\]s��u�V���;O4�z�%��fs��5[U#`��IĹ�Rzn�]R���a:����؝���9,M�j��i�Լ�P���t�e�˕���Eh���_κ_r���iZ?�4W�S���-3=�$dq�<3@���ΎӅ
�d�OG>��Z�&�:�z�+p�o��5�X���/Z%-z=q?��nq����DZ��B7�����G֙�6e+�@���j�z196��"P�B�����wm�a/�g3̮����g9�y��#.?3lrr^>��f���o �fWlDp��+����h�����L�%�n��:��%aNE	������j�(�D#������y$�1`"���7 ���>~�����)6�bnBo��/������bo!~��F�@7��z�wb�]�ٷ�ub����E��m�^lR'�,)�lr�� P�N7*b}�]�������[�	�E8 |�RL�,L���Q�,�bl��d�I����2å9�˲u4��� �-��C薕�p� ���r�1�}ʆ����ɢ���s�B��V�	���A$�$�q1����z1/ďQ��g ��h&H�ϐ�{����
��L�^D3����<��wǘw��e&��@v7aB�x��m��s���D���ٻ�O^�|[d�!�Z2|7BD;����V��|3\��#�F%'�u�8-k`]�e��ߕ�.>8��aN��1���xW�}7����*6�
U�P)�s*�1��58�+����ŨSŖ���QF"G٭<r	V��2#s��)ݰ�����[L��s�3��?����������m��!Q�h�$�r����<�������sT7���5��Ow�I|Ş�s�L%�w⣖���T��cf�x�3��+�<~_UZ)�_�/�zt�b���|�X���tѯ�i�h9���n����0������>��v���,�\�g���h�qT�mwo����=3��^�3��c��/Z�mS�mk��Ź��z����9=\c��+�q��
$4���Z� �ɭ�0�>�4� ,��)�Z-��@yv��|�n荎���4`�"�,�ħ��tɸ���Ġ�����M."��m����m��}��f2��o��>����P�g�鬪�.-z��t��~ΞO�Y�)��sH�x������d��T�<�x@�^Ui|�V��	ź�ȗFQ���3�t�@��ނYk���}[z(���k���M�zw�3�B��r�j�ܧ;�lw���sY�!N}ƭxʮV�R��:����e�Ta̻V��e��.i|�p#����s �f�dd��*&w�!Mg���l����}��T<��:d�%x?d�K�.��8/7��|��g}��g�\�6��Xq]K�5i��7T0�Ҟ+t�`Q�m�9����g3�� Y���n���A���{J>).���i�7ދ���C�;V�>X� v������Z�D[) q���w<�wy��52�]wf~����;��qVg�t��Z_�$����k�V[��1u�@�H�y���c+�����Ob��%B�wg�jΈ|UtY��t��D({=�	V���P�?k������u������1�X�[	���W3��
�O�<����4QRƵ�e�R@}�>�&��c7����X/
�H�*��C)F��Ύ�Lc��l�y>��"�n����t�a%\����x���ݮ�ݻ��5�Q�7�ݽ��<�}apf���>^��>����'/��s�|%��2O�߄[Xrd�a�7���K �I�;�`��y���x	���r�<M�p��2պЄGiP<�PP��T�Xj������Z�9�Vw��=J�y]��y-V�*����ur_�8)2���b7�D����\O��̹�w���PV�3�?#�bq�
X:��-����Q�ﻗŭ�ϚBݤ׃/.w�ݓ���e�1j�)X����vu�I�5%~�l�@���I��?��5t�j|@بa�8�@A�0��Jش�Vl ~�5���.���C�F��>�`-��Y�eߟn�cpf��>X&a��i��Ic�^�Y�]��T@=���	'�<����P;_x�L��lh8͋o����k�����Yj��e.�x���q��բ���& V��9�<hI�����M6�������i0�o���E�[8����=O��cz��C����v��j�"]O�<5
�\��(��B���dOJ�
4�0r�~�0i�����xi�C%^�U9>��/�^�Y��kٺ��H�%�A�)zuw[�C=�7`�=��;�eP=ja/�G�Ul��T"�iR��c
��TV���r�g%��s!��p�%�t0��d$��°�����-�d�*�������=��uu�H�&��P?w�t��6�kT�?@��R�vDH�{������8���9��冷�:m\(�@�?4�--�љ:Gg��ۍY�Q ���|��e�%ȮY�$%7K5�Q��Ke����ʙ���v< ;�ɸ�'�{s�!�P`����Ϋ��C�^�Ul�ԔO����2���*R�:���"����o@J�����Gg�n�U�Z4�%�v�жLͽ�O�SN�~ҡ��b��\r��ʈt��n�����d�UX���&�NX���w��T��b2T�X�Q?R�"�J9{AL^}�@�nfo���'/�σ�MM���/D�]G�qV�{��������\9�3��g ���U��gs(��Q��	X؈�k^tM����K�a:[`}\�c"p�^.�b��(%&ġЪu
��nO�7a��u�Z:�[mR�$�F���軄蝚��f�� ���:g;��	���P�]�J��z��橽-��_nSX��0��%P�,
'��پ�K��#�ًE��Bx"�"`X�(���?
����wy͞��%�[��fQ��I����n�nX�G�#�&/�?�n�=����#t[˔���U�M�AY�c@�+��U(B��P�d�t�g7��LC�����TvY�!��B�SҘ�F@��}���5�o��\�͘y�P�D�� Ƿ�`��+�[7|~$�NXظ;�߲� �*�G�>z ����("��.�k؉p��-����*���t����ށC�v<ē6TC��s'�IND xѠ����h�q �WI9�y�ݦ�E_P��l�U�i�Z���&;�(�"X@F3F�I�s�2����ݕC}{�.yu��"�ɍz}}�<q���s�֫L7��n�P�����s�W�5�R������^�ON6���B��1'�U2ӻ���-,�����^�7d�$�R9�w��{|�9!Sro��/z�H�Vi��E�*�ȣTf�d�<���� <@`�I��?ΰs�>�f'�
������v"E��D,�)|mU�����T��S��]rG,����7�e�N�d�,���EK�;�����-ܑ)��q�/�_ƛ�a(fŷ���4��g��҇?&-�b��$!}�Y�����!�	E�@j! ��٣LۊB���FJ��$�:(5D��lm�ƍ�X���bĘ�N���b@8��>�d{��!�^-W��!9��i1���ы�C�)�^B��}�:}P�
��X�+�J��.ƹ_d�D�/��{`����֙����	�.ŴIh�ZD>j*�����7-��$:đ_l6،X� �S�R�N)��	��{m���}�Hbaьߣ�-��ߪYF/��Lah�(�>iH�R椂��x�����5I"��.;P����r�e~�%`�i�~��4	����R�k*+�&��~g�_w�@��%���p��c ���lZ��K���{�Dgl��q႕C� �T`��^�����@E��,7�\��o]g>�K�?fF�8��2g�]h�`��{,��P��:8h��ijzZ�	���=.�v�5�	�E(T�C���j�MqZ��j��̞7�4�X��P����ooX٬�;�IA���M7��g���O��'��4(]�14�h� 9,�ssT��;I6j͢M���IN��kL!��2HTJ�1g�l��ʋ��kb2�K��ސ�[w�])R�d-�J���-��uޮ�"w�;�c�:��[��:��%��ݭ���D������I�<�F�)NՆ��EJ���(�����X���|�]J����i��Dr	։;��ðc�YS�P%|��әX�Oi��������������F�1U�|fծA�H&}{�eF��9��� �i��(��s���4�ޯH����[_��/B��9S�Oʲ[��8�E+�$�IH�N�u��lnW����*#���pΖ��6�K�����#�ࣦĀ��v*ƽJ�e�<Hz�����"qmw^�� .9���ΦU�m ���a�n?�| ���o4ܾ߲��d2�Ñ��qc�eb�~ā�I���XQFl�qB� 
5������8�^n�~�Z��"�*2�%��a�*��ׯ�����zG9��rj�dA�I����j�ì���ү��?㴺�H�d��rl��!�@^�}�ZL��a9�B�n�������, Q[�S?�>�P�Pc �f�>���N#z�$݄H��L�|�	��?���,m�[;.u�b[���ٸTߠ��I�,(��]3AҾq��NW-PTh��e��ϱ&��ND͔Џo��ޖ"�B�b�WF\�1X����u>���/ƹ�k��R��M�,�c���[�p܌e�]���¬���y�U����sX����|��T���G��*U)&N�*���,fFG����X�|_h��� O���l���qGD�x�U��X�
�6�u���t-O.�c<L��)�@k�������S�k�j�Lv�CC��j�uN�BU<�$�/�����`]��DܷVLC��9[0�h�;2���g��l��5�@�NO/.^N�D=~��t6�dO��0Cߗ��R0�����/��! w��i@��d�
z��b�j�z.?�A;��%�l���ޯ��aV�}Чښ }�Grُߍ}}�,8�=m��=��K����no]�\[�>"�lw?]d�о�ߨ�:E�\8�$s�p����<ii:K��^ �������3'����o�p���D�}�)?�|9��'^�d�1X�[x��Oo��R{��@#����7)��8�D�t����i�d�	����2v[�ݩ��=����R7��Q޿�Wxn����򽟢�QӍ�P���V�S2�P��H�G��J=	]��i5{��!l
�x�$pu�7�䊘iE��n��M_-!3xGL�{��6{x�~�����s����MmeP�ɤ�n�6����k!�X��JfEd&����k�2� ��
����٥��C).۔�����?��خ�#T����I�E�&w7�H�
�i��:�����o,X��`�\H�9�'S��$��
p-04���j$
��ݚ�f{P�E���W�{:�w���F ��#Ce�M��0�^�8�~�p�F��)_E�S�H��t���ws���R쎭�������X:���vPyoM~���XR�Mҡ�޺���uFF�V��D�ѯk��Ѳy�~J����.]��.�S�s8�hɃ��ǲu]g�"*kw&�s���!�E��| Lt�Z��<� ��Ώ�FEm����c���_�M���|������z�#(Æ��'��jݐ޲�]K�e��i��<�C��h�h���X �+D�V`i?���:~ �O��*���7��V�v8-�煮2$���ݟ��L�� h�x�$J,.��4�"7�mȻ��D�?5�Q���HSr��T B�ݣ6�X��	:΂�5}���`!s��v gʤm�m�����L!�\������7J��o�X\�b��2�L�bi�%R�Z��f�^�/�D��jTL��>��S5d;���|��G��ES޸�D���J�۷�)�P���%�bI�p>�`մک�
#��I�8	�	�ЄQ��OJ�Y�,�/�4�
��f%�k��y�Z/��A�O�'~}��8��ڸ��
B�G��}T���~Ҹ(��FJ���5xx;g,@� ?����T�=�q��n�1z&"�#Ч1P��W>M�/�P�Ӱ�)�3-H�G�uf��)<�c{
Ghf:��ȿi��ٶ���K�:O��Y��'�)Dq�0N�=�E�?	�%��D�؟�����h5�xBj��	�*[T������XS���{�(���j ���}���sp�WM��� ��<�����t+��)`�I����1��|̧##�ܬ�����|�$2oI�L���L=Bg*@̮�q�O�Ty��*_(9=g/d_?�E;�/��LZ�����z��LH�]p�^v#>�2o�`�x�Fo��hD�ڴ�?F�m�v�%���"���7�s�
DJ��W�f��~�FR���$o�J$�7B�D�Q����*@�%�g	f8��w�`�1h���TNf�.��[� ~��ӡ�� �J��<��0R0�bS�z
7���n��e&$t�T�Oӄ��P���3-*pb��En�ju�t$$0f�M�I�mS��3�3���-D����2�t�p ��t���9�v�@U��9̯ˮ�%Bd� �M�!a�4��P'�ר���s���9> }	*���E3"LO��(g8]܅���������2l����!�5^�Ϝ��R{y��s����Nɖ^�M�t@q���Ĺ�d#�T��ƻ�c���0�obBჯ�~{�����.;Ӡ�;2O,l�ʐ����������"�xc]')�U�cu�,��bت�v���gia��>&ٳ@�����a�AB��}.�'��p}.fg>�3L���O�u���/ �&��;ޞ��V���q��U�f��-my���$t���b�3��t7�j��#����M����&!����1Н�TV��1����K�`7�=��T>L���9t��'e
���B��A���2���Pv>����I�,`�� #2�D����#�z���&�^�-]��|����O����gu��ch%�.��1�\]�$�\�e�ZN���υ�q���ۻ�d�*�n<m�1Q"Q�#��u5_K����:3!��Uy}eO	�ӯ5 xՁ�M����=]1�9j�@n%$�M]��ɽG����7�&1a�Qg&�x�%�.F�NRu4�yqI�\3�c�-� ��t��6�`ǫ�
0�ÿ���n6a�b�@}$W�W�f�AY�$��N 	��CJ"��/5���
���!MSѻ�W!�� @�F��:��|�[���|2զ�6f���]r���i�D�'w��fe�K�����^��-�!�βȁ B�\��*r�ut�fZ� �b���ں4*���(j<��N��P�&g r�JT[���g�����B>����tk�L����>Zo����0Cݓ�. ��-��`a(4�����T�C�Sg#_�6�e2i%��t�Q
��haS�Z�G1�5_Gr9�k��+==�O��]'l6�@�o�ıN��i�ݍ��1�m���8b�P ǩ�����
ÿ�O���`�����`H�Q��&���~�*�;���O�8H:ȁ�7_�~�+���8̆:�!'���Y�q��t�dT^���+<yk��Q`���=�v~��Ab�U��}���A�6���RlbH�{��=���ٱB�J&����ן'�v�9A÷��,�� ��~�z'p7gw���h��\)�7k��+��'���%��J�	�|�L���6�9�� O���~ޝ(JG�El	Xr���QYP�a�R.��#ϸq��D�h�mk���7��R�]�Ӓ[*�7ϑD��R[@���1�F`����9Ӎb1q�"�F$8<��
]
���EU!o����8�w���UN��i���8����Ɩ駞�M����+����:yP�4�����UX��1gŋ��_ix\haU���X9� ��z@3�޼H?���c �M��GAz,FM�KDBP�9T�w��8!J�jf(e��
:��u�XRrS�I'@��۔�6$鐇5�a�k`7����o�tmJ*Qd�u�b�EdKB`K=���` ��wY�����Tp[��;(b*����{'k��	��L�B����"|^G��.��
�C���Z����&��;PVVI�%��?ݶ���yaf�"DU�Q/�84aX�Ab��E�����yE�@��Fd��A�	����"�bl;K���b|�'�6�	h\��E�@��Xd~�\b�Yk�����z�,6��~Ŏ�柃 ��m"
�
�;���y���`� ��ʆi����K�D�"f�k��}��Od���a�9Q9��P�X������{$�O.�,����k�j
M#���(@�_�R���>����a܃V�������O2��	�͡����] �� ��Z�rXʿm�.a��DiN�e�v��anԑ��M\&��|`Q{_�*p�`���'Y�+��-�H�f�Ɠ�uC�II�� (G=�<�0%�/�j��f��e�������P^cc��_�V�{�.:�G�n~��Zq�8��?����re��%`�5D��`A�s�f��O�cAfE� e���f�9P�᣽3�5߀Vq�ƾ��4�EϺ��������D�]��;M`F�n@>0ǂf�4|�o]��*�2�L$��ɽ�rr4�>&{Q��_�qp6�y�`��D�F�~�NGJ:�E%$m�.��F���2_>�+	͟L�o��qU�J���D�h�2;z"��� �7�L��z|�G+�6�������x��D)%��b�I���Y
��o�'�������ƒ{��或/3� r	1U�h 2���=�7��=�Gu"��(so��J&���\|8a��������=�J�
2�w�)�j�`��\�Q[R@�`S|B4�����
�k��]��%��2��K4E� ��}�6K�F�J:M����>���k�6b<H�̩d��3Rg�����I���$]4�?'m���Ue	�Z}-����Q2?��cD��R������a����:I�-�֕����^��P�~`�V6"-N��ȸ�e�&�T6�t�
��%��vւ�i�`���xݾK��/K/���X���1������w"
���G��0�|�p��p��7g)�T{�\i�G�Ư�bc����8��Ѷ>bS�qc��!����_�=���s.٣©�*:�zK�"�ܽ�׋�o��elOq�������ҡ�򪝎\F�X"[�Tg�?B���pa6�2�b���Ŭrmn�O�
��Z��qHオ���',`�{?�0��]H[�:}dҿ�[��������9wu����wJy�8��=H�5�z��-h���=�3h�A���;ҽ�]DN��?	P���6l�[��a�;�xKɒGG�
��>9>th�yot!�T�`P`^��#{2����.P��n}8G���̌+�����MzW��9�4?�;K{�-�g$��+�y[!�Has���E||�_D�B�<o�I��C3.{���4b'��,�8��8Y]�|ʑ���~~���j��Ü�x�����0��Wh�xө��`IdXslL��v��t��Xn�j���Aȷ��=Db	o�ֽy�G��՘+��	a��DD^��1��W����~�3E��4���--[��X��bQ��u�����&��U�H{a23�
�P9��4S��i^�v�R�/dO�|#\�$�V{U����i�i4H��Q��hGS��@���<T}7%2=�eq� F�N�W�6�p�0u���+���og���pu�B,g���O������ XK��L�d�]�i�8�b�F��+Mu�W�6`��h�֯�Y�!_��\>�͝���I��o��Al�_PI��xK���3퇂;
�� ���z�Ņ����G:2�H��d.z�D�4 ��W�
2�̭�S���z�e��Ce�����1h��q��ۍ��u9�N����N�������+��o��`#�m��3P֍eNI�`*��䊾09C�U��ŷ ��u�2[�f�l�3���[x�ԃp=���{�.�e׵-�|���Y�!��e����]�'���=:�`:���5����k��V:�5{���*F���t-`��eaY�*n"��"jkw*�Cֿ��^�d�<A�Hw�&)*}�_.^�j��PD���c� �hj��?�F�܄ݱ��S4wʤ�k�m���<��r,���>J�ƀ�����:5��؂��:��}%��Q��r�ޱ-�cNB����6��_����b�O����&,%�fl?�v|e=c'(j�^k5%���DϬ�ܣC�r�M���!#L���z�3��a��a��!`�m�L�R��v�l[hZ�ÌB	y���vwC��(�����=�.i{���v\!W����u9��jPX�cw�OY�w'��}��V���#� ��;۵3��J���ɤ�T�M6�mA�F�ֵߗ�v@�I-�f��b�2����z���M!Z������y��Z�1X�`K(�Z�0�@�w��-V��d)�<H�ӧ�(ں�v����'{Oמ�Z�n��1��V�a3�#�l�;{��kO>oѳ-���;}enh`���Ə�1��k���K�t@Q ��sx�~���C(�`k��
ZS�k� �$d8��S\4�J
{���=q���Au�L�X�]�$��þ_���44Jy�a^��b�IQ�-\��&����RnP�eNh0�~��RH6I�x+U��b�\*�@��K�9��!I5�o����R(v�J:)��\�v_g��Kh,$��R��+O"[����#�`j[E,
}3;IE� 7�*�6S�i��]���
��W;�N��R[U�lQU�_���8T��pngq�:]KD���"�?z�6.kW��T��&q�אۻ��.=�4n�C~�)
��DB?VU�n�m$G"��u�2=�LQV�gh�N �g�B<�����ˇ��9�z̭;!*���SvIp�V��Is}��g�.�nJ����U�F�`�<㞢sU�����)�S�(u'�c�H��A�K�h�B8*	j�z�	z�
'���u��
�ỵ�V�:�DI������p�'���s8�b@��	v�u�ťKҚ����V������=C�-e��N�-���}<F���-�>4tp��-`�[n8�c��_M�	v2;y�D�,-b���)2Uz�rn_K@8
t_R\�_��8���+�`��`&1]����g,D���o�<��%Q�9�%7�%Go��$3zk�c��奊Y�R�� ���I]N�H�M@��זn�_K��{Ҭ�/����[0��;�G�-m�~%�P���J;Sݟo�wP)u8ϥ�z��l��0ɜT�`}?�FUG�8�=�\Г��C�~3���>纁�a#�Dyu�e7���d���j��\=Tf�&��K�SZ�Ɏ`���a�"��P��'45A%Yۘp��Bo��N�f
��ն�^%[����wk@���Y����q��ѥ'e;��^��6]jq�g{ 8���‐S�&��%�5	��fʌ�X�d�������UK��CI4�îvẀ�	%lKݯP��D-P��Wf����GZ�˖%�=g��%�-��Xr{�^hK�VI͇����G-I+�_��8�Pj�0t�~ �m^�D䱯.�?�XN�U	��'��i4g��Q���c��j���ޔH=��]��^5D\�A�K@s
��-�n@^��
�2�[�:9snu!8�T���(�����H?H�v37P�a�{�3���z�*StT� "훽8'H���:�mqE�^j*{l��&�'���a4�A���7^^I�����`멜S>����f{��{�٘v�ZZ�Ǎq��L^ۮ��g?��I9�i9 ������o�om��`G��\�������b3�)q��u«NBP�:�d�6 Zo�*%���wڤ�&��&���ý�8�j�+wl����N$<�%����-/J��"��}��'�g��Y��~����!�$3�k����u�5&�t`�&��V �z���\����~
X�B��Pv@p���N��lS����.�k�\X2��U̫h��5�~�|?��o��7�b�^)c?oX�W��}�G<�U, ��l� �;�����$���Í�0��*7���;�L�9��N���t8��w��^M�����Y���]�f���z�AS��֑���W�b}��� (��@�:��La<c ���vo�a���i��L|�Ui�1c�`r9�1�5el[�I�s�a�U"���#w
�qP��
��6�2��du?h�S�A�
w���� ,����MtH`�; t�K���D<���3���׊��N0�-O��$��\fwH��P�B�'�Ã�f
���P+Y����s������-Q�K���@y���(�!H��L��uA�|�NuŦ���p_�rX	��U��n	�� ��WP&����m�@�a�������@�;W_,�zt�7��7������a���O����;�% r�O���Ђ��\���,�G��4^c/
�R�-S�� \J��vY�i�$P�Z�w�N��S|�BTD>mP���pT���\</���M
��qD%ᮬg�C�s�Ⲫ5=�n��u��E��M�M��g�M���v��b��x�2s�M�}�
��vGi�KRa}����;���M�G�Ѿ�<��Wjȸu�� t?h$�;πK��)�g�_!���=^Y���ֳ;B.�Ly����7�����f� ⍭)�����D�w݁���k�� �ۺ/Ht|^oC�t���򕌻{��{�VZ�~�e�)06w��z������fD�)�ϑ&�B*���x�#����������uW�4�mP����h�ڈʔՍ�������O��1?�@��m�����Oqۣg7:T)��������K
��ʮp�ܚ1O���M,���˹��Dn.���!]W�Ө�G%���:,��Jl]d"��Q����<���j��B�<��`x�PZV��f�� �IW�����ӂƵ������zt뿤�%}�uS{���Z?�݈NRQ�H�����b��&�W��Tb���|�dܭ�;�;�qU,�VPK�^������S'@�֎J�%�l����/�m bbQw�넧�ϭ�~ᇽ�-���X�_T�Ӵ�i$��RǛXLд����,Qx2z��-^��?����_���Uۍ�h$��.�I:js-?:>Ls�J�y�h��+x��6q��b�?�K��$�
ťTk��\R��:P��č�pX~��V����f�D��F=<H2�ۅH�L5=���n9f�eS��B76s��i�-��X��[B�����bs���u�x�c��nm�,����V�]����영Nb��1�ZŃ}9��ڟG 󵚥���0ԩぴy&����?k&1��?U�}����Z_��v�������L��'�嬔dHf3>nv�^%�Md�2�2}��4��p9�x/��q�eg1Ym�YX�=2����qb܏%��*�KCCu�&�9쏉�� �ۤrG�H�+���-�(}w㒪��Ĳ���Q	v`ij[^�g]�� d�y�o&�����ub�W)�%J���2s����)z��s�*�S0��W�<3�����\`Kw��q�J\F����]�o�ג���Yų��뻇��w]l�~7ch���$\cB��W@A	��K��f�3��r���yKMR��=�Zu�E��v�C��{��幞���>;�X-*��Hz*��r'�o���287��g顿�����p[��IM�+�!�;#i�%��,E��I�����j���s�6�w�;�{,��}�������?�e-�y�n�dp���#�Թ��jb�OW����w`-Q�j[	�S�e)��Ph��s�A�s�W���z������u����\a�ҙ��K+�J$y��M�~E���'�`����3��Y5�լ+�w��;1�� $�ق�p�]���ݽ��fC\#���Ϲ
(���+Tևڥ�w���'/a���iR����]���V<P���{?�7+��aVs�׼�$}����Yw�m=a<�L|���>���*(�g��<d���^k܄��{-llE�U>�GLR�� z%9;P'z�G�YF�S�n[#�d����]��׍V��`Q&�[}[����s����9i�Ѷ=f핽����4�q��������33�xC��Ps���o�ՎZi�حng�q�d+�&ƀ����LU��]����d�T��!�)��fef~R3X���-TGo��8�=ʇT�G��tn��O-x�B�r|�m'���DHٔifpG�rf�Í�π5�qv{I�!J�9T��KE�\��+�k+Ʃ��O%+b�
���q[�r�xB�\z�_π��1�T>+U�D�� ���J���i���Nm�jo��m?Iqg�, O\���ki��!�~j#�>0A}��u.�|��ĝsS��T���	�;Ol���I�/0燛��E������x��7�so��[��VTJJ��P2��m�PIȘB�1dO?E7�.�2V�̉�1���J(2�$�1�޵�^�{?���������g}���}�����*_�� 3���v'�˘�Ï@��}}1�����[o	w�ybG>
�+��z���2FTCދ0c�����6>{� s;|�{d���*+]�ٝH�]��<i0E���~��F��Č����fOl;�����%�ڿ13,�㬿�(.MƖ ���>KH���0ad�J%����B�녧�~ �o}k�7�_;-r��O�nJ��b�v��`����|�P`:a,� �x��Ir4��,Y����%Z�N}}��B��r�O7 X�Z����IL,#X4���6|��U��f��	�7��iH2$�lqX��K�"��%�STJ���T�+�뛋ϸ���V;b-���%�j�~t(,�B�������v	Pw)�BUװ��i�S�!�Yl�;����e���R4�G�s����R&���A��)�"S\�	�;��T����mT@Hqi�y�ga��:��&��,�z�
�zJ^���{tF�
<�?��"��/gO����w��xU�Y��#�bi����^�84�+����~Ք}(�O���@���ҹ�͏bJ�re�UJ/�q��8��w�H5 c%�8��	�u44��Xu��!#\QRH�8٣�̕Zc��S%��|�ٗg	��p�p=��1��롊J2�}�Gkp�N���O3�l�T�ʴ<'<Ɩ��6$��'x�pUZ�<���Aȹ�|�f�����E��s2k�H�R#@R��A��S���ւ��[��\��Kq$���)�����xH�uvV֠U)b����k�7r��[ ��S�>1렔}�ίn�8���= ��U0$�w����"���*7� t��v���O* .��7��N�8g,��7R��̯?�A���c	t �"u^\U�ʲ׽��w&�rIي��^O�[��m��.�j0�V�m���圣���,�7�4~8��~RS��'A�tv)�J�; �Ȉ}�>Tx���{�z���p�n�b2������V)��V)8L�m[eoo�G��KJD�?�v��5?��˫�I?��R|�#�����Τ�?i����+#�{)�t��/L%<8C��Ɲ�/��6k#5�4v�2q
=���l�uo�/L9�b[e�����̯z�ƀG��Є����d�NԸ[��6�Wӧ���{[�L���5�n�1�U6 V�|p�X�⾆���Θ�#������D�#�p�O<����5�E|1~��ͱ+�7�^?�EX/��ǿ�U�-�4-��0�aS3�@��ӧ�+�$�
e�I����U'�U!jqj]2nݭ�m#+�����c�4�Fs���ރ���e�$��^�x9��*UF�韍����Mw35�,U��r$����)-�Y�p#���{�u�K�,t5>�M[����^ԑ�{��a�z��N5���s���x5�q�><��68/��E��F?�oߦ�	�Ur]�}�\�UO_E5X�-Y�f����}Ʌ~���J bo��(��DD�7�뢈m
#3'y�B�J�I�9C��Dr�l�s^�0棹�{U��0�wDzM��� �< ������u����v;旳oߴ��vϖGj��=v_�����NKň���$oϗÐ �ג.���!R7D� C��ex�ǿa�p��z��yfr�*���`k�}V��N������Gtoh���-`���%�N/���4��_��K��/�^.s�耕���%��hu�I�X��nL�u���g�6�R,�>�{԰�.�1�;�4�d�Q�]:�0?��� #u�_�v��m�I/~��DaER]%�A.��υj�O�ֲK�>s�ݛUU������77�Ϥ�uț�?'��<
�j� ���%�G��]���t.��ːܮ�^�fߛu����ԩ]�!��~QI/Ĵ"�ވ;Ʒ�rD��\|G�V����?_V~�w5(���k	���_����c�����������~�ߏ���?�����~�z���F��ܲ��}5����{�	x�?��d<F���"Աd������QgϜ�����=Q7r_'����^k��b@��]Zk3$�m���`PǨ��$��B�4_Y;$��,MS��rjω+{&�"�M$��c/i�y��D�vy���oX��b)>�48b��k꽋Pӂϻz'+8��/���z̎��>\���Q���?�Y,H��@VBM�A�⧭wE��L���O��61�;��sF*<2�\���.��,��#�5N9S{F0#L��O�ч����|�9!���_[(C�;f~o���X��͏.���`���7�@�{~#��M��kpKt�u����Tǵ��Ϩ�*�^��DiE�%y��fGJ�-�6~�&r����=ﱥț��r�����,�y���;�	2��������71	�\hLa�/��&.�>Pݑh_*r��m�M)��k^���"rY�J������-bm\�������hB����\TQ.fJ���ٴ�/]�2�/�_�W��v�\���C{|+��R�H��ZΔ�������zXLaޱj�?<�s���/)��X�}ؓ����	^̮rQf��k	�����}�/<�4�i����_���B7�j�0)�Oo���/A�af4^|����욯ƕ��W�8���Q��U�r�]�{�U���Tj�8W�>�^�]�Z��p�3��?�͸�9vL��#h�-u2�W�
m��l��G�fv�;�\lx�O�o�L�������W��G����n$�F5��qa���W6�J�:��m�ae��t���u�r�� 0�8�t��s�^L��@l��u�u�:��.�&7�z��A��a��/�z����h��܌n�>�!���eei"5��C��[3dQ�`��o/���2�X���g�]�2\���N�;`�5��Sȓ+PL�cT�G{G���2+i��d�`�������?.�W}�f��(�b��r���Ć����.�	�����5r�~�ƭ��T��]#��:u1��Z������+wjB�L��].v)%=�&�C;8�U�e>tG/|e�Qs�rًS�T=\>��Z<�"����/�4j�"���Z��t���S<�%#�D��q�j��>]���Z�A��'�C��%�h���(�����$kQ��� �D���&�~�`��&-]#��\HG���l�[��4��Ы7a�o��m+!�x�Ջ��N�&����4h��Q�"��j�W9_�ӶR;a.�Y��ġnZok��W]nl 
#_��%�fT@SUw{���e���*x�gZ(�f����
f�e��5-��?�I��L䉔5z�����fx�R�KZ����x�)l��5���� 
�WjS{a�_�O���ܛ�;���S{�#�qD͞į�I5oe��r3�֪���8�l�]�cba+���B?XM�'f�vLˉD�0̅[�9�]58/K�ay�E���,�j�U���f@��Q�-?Ř+ze�6��q[�?|��/R5���EC�/��-��� �2� C|JBw=����vls6��$��԰<x�.E`��I	�}`4ou9#�ί��o\�K̼��D��'�m�X���&#��8��C^N~f{�\��Q�,	m�}-ݮ��=��z�T޲��$["�=�r���Z+���y��%��Cͽ�-Z�J��Iz��ݦ�H��%�ư��.�8����e�l9��"sS nQ�i�Bw�h�ё����㱘�_?���P���q�� �o��iZU��rގ��n±`� �o��Py_R�9�'|<��@D�	����O�����r�'�6Pِ��ˌ��n6�ij*7�7lpBȾC�ø?L�:O~�8�r&	Rzb�q};hԝ��bq6E��K����7�f���n���E�4Ʃ�FQVsaL�t�v|�j8=� t�q-3����m�h���N�\�z�\���t���7Y�����6�Ӵ
��@1�NO^�|ޝX����a�Y	�/���] �M���	��w���7��5��6�¿�9��o��7���ݒ�1��uMQ7^��^������/�in�>��>�Z�?�^���0�}P�n������/�����)R����m��k�6����H��<\�� ���x}{E�iL �XP�9ܥ�S�:��w�V>c��BU��7-_��Y�ϧ�ǅ���? y����~�� E�;�6@/Tyf=�?:Tje\��������謊�$��<�Ǭ��������G�Sc??Q�6���?B`�C�D��pg���q2l��.�~��2���%��{h�(4JB��(�{YF����J/S����r��w�@]��z��1]]�\��1g��h�e��Bb��փ�!��?/�v^�6��i�A�[�V����/5�0+o���v������gJ��W�B���N�8+���(S"�s|_0��+W��g����n�z9g⫓�Q�~ʄs��d{MB�-\��B��K�MW<�U�b�Ɓ/a��{�D�h�iQr����b��\�B�\�B$���D1��Q�� N��et_.1���_Hjۮ�3�zq:�]��l�v���xܷ͋(B�r�����,d|�A�T����emw�B#��8��!SGm�U%��R�#�8��)����q[�S�n�-�.��\��[s��ͭb�& �ҍa�5쩢B��1�}�\dzx����������&�·���ޑ���Z���1|͋1��2U�!f��)�����G{"�����DP��;��!�~V�eum|'��4�3�%\���co?;�Z���Y!�;�t p;p������O�!�

3}�P�n����/WU�E�i.(��n� �J�c$��Z��Z,�mw?�A�j�<���r�\�ǂ�NݵP���bx�j��v2�N�*�����0��:����d���@���j��.������󮓍7���Є�>�I{�r�g��q�&��K�}�m㋑0��6�Y]�^^sã�% ���<ئf����!�#P̓]!�%5�d	��B0�bDA�g�E5�=[�۶m����G0A��HO�P��'�O���e@��<��&j\/��#L6Z�h�vt:�#+�o*Y��ǣ�>��ͷ�5]�A����]�75�r5]�#<7>Xδ���	���mkZz�o��&��w�XZV��K�D������8���P��D��ti��RU�d�gM������z��W�d&�)]�N�_�O�"�ޞn�T�*������A���8���]Z3SF+�~�-�p��6S��S��^@�1�w�?�]Z�YPu��3?oR{���'�i�ԏ��m-�:�:���Q�����,����e�J'R]�^���s�"���PI�x`�o�S��	�\�I��eX��)�(y�}��#�Ȧ�Ar���.��$O4�w��"b7\#�����u��G�bXWi3���IQo:�r�c�b��1�84=�H�r�[�#p��e�� ��3�{ŃF�1�]f��� ��KD����Q^+;��9�~��&�U.�W�b�\��0�M�%�z��X�;u���p�惤��MZn�Q�2�ۤ�t���4��!>�pi���vm�MѰ��@�m�okT������y�>&��%�1A[ZA����v��qW�����6ǽ�d�H8s�NT���J6W�+w��1�R�d{:�$9���x�K��/8��ZV��{��Ymz&]'�sk�Lȁ��������t�t`Ya9��1c�<�a�*� ��M�-���sig��Ʒ�Ąw9;��H7�]�=YI���t�E?���J+��׼�r�ϟ,�t1�J�	ty�_ENI��z�x0�Ct>մE�,�P��i�["��xX?I���d�`��6_�������K�������?��1�b;Y_��6�okoh����oQ^�V`����1��e���Ԫ[��]%vXhCy��z�{@�l�ʹNUb���K�p�����oZ�E�Z�f�V�n���+�J)������
6�sl�8�㻣�l&�쉣�!gC���q:��W?��0V5�W������E"7+����
�Cb� ���,�9mR�[���ݲ{�o�7e�^�ͤ�(��d��!_/N�&׬c�&٦��3�*�M&Q�'l������C�w�n�TG��1q��5���DM�y��5f0i�� ׳��1�,���Q�
�_��4�F���~c����\����6>;m�i���6Fo�SC��	I������yե0�`���;��4=���HЀ��9�#1���/!�w=��`{.��n &*�/��U2���Ӱ3ig7b��گXb�bc�����V���%{�cD,8#>	|�(Ӏ��՘r��aʟk���4�n��s���C�Z��1�ˣt��S:zl|t�m���ʵ>�@ڐЦ���M�P�7������{�m�ct���>B�%�ٴ�.g��h� ޔ�ؼl[}����2�0e�O��fw�ϥ����9� cV�E&�>�x�-nߍׅ�h%�
 ��a�ܬ�E/���Maʒcv`yG�-'�`�Lq�̮1yU�<$���&o�(�΅�� ���-��$�%�N%G9'C�`-������Y��.��ECp������8����U�?��nw��d��
�����Jx�C�{B��e6>xTM�/��߾�0�M��p�K�Ʀ���n� o>�ax�~��ݔb����=����<�� ؼQO��=+qs�Yk%hg�R�����l,S�b��o�U�<\����o��S��ȟ��M�-hq�l��ܴLL�R��X�][A���B+<�����Vc��5�,��h۝`#i_T���AGK��Vt��}��{�rtDBR�$;%��衏��� �a�5ϛӼ��j�;��;�abp�A�V���~�������-��	L��Z]%^/Z�\�*��Z�x�~M���y�@��1np���$���0%�5�������]���?'���f�%�7��z�ѳX�o�q�F���I�o@f϶�;�q VU�@��]��nPu_�@\�'WE/&���}�5ƃ�+pL��'�B��2�����r������;���N�a�&6Uq�{�m?�o{uDɳ�|���tzL��苨82+o�v�Baoz�`�@�� u�0���b��W�z��D���U���'"9�w�[ԫ�.Nq���di������d�2[�Nnƽ#,�̲*C1ꃄ�o��;�����0�'�݄��ԝ\`Ru�E7�m�"e#].�{[$�O�eMg�MQ?�Sv;\�j�dP������2�*y]�	Rɍ�Ó�	I�X��"�s?�7����o��F�v]�����y��}���fc?5�<K`�{�
�d�HӁ��e]�&A 1��#=�o	��(���`�3����Y��1�Y
4ܰw�T9_�H��ݍ10\����%vPo.an���D�NƃӍ���I�E��5Ly�!a�
rVL�^�Hvx��J%S�����)RHy�܌�����)q�}�"*�M������j*Y�?^�%�]�v~^� �~��i�P�V9�\�ĜxM�{;[�2Q2�Q�\ @R�^�e�g�U��jƱf�&�M���6nH�-��\�7㹊�$����ʲ��ɦ�b�=.��E�<1j��u}Co�E�X�����@��Et�7
C�4$�����u_�Z�&Z���	ZS�M�^��tQ;�Ά^ÿ��v�X���ޞ񂖋�$�Z3�ܰvv8r����'Ԏ���poJ��H��'.̺Be�����W�~5���>�H��\�d<H������� 8v#�AkH,o���D���#^����o`�O��Z�d�as��ôF5�ީ��.U� �vk`eBF]e�/?���7L9ɯEOQ2��]w�l�zE�%�MQW v�3��4�i�R���d
�e����[�p�|P��0���G��7�}���F;p�ob�ڍ�>%�V���ז��i;�ڇ�ə�%#ҬvH�����(>�v�l�O�f�{Q3��S�X++�� ���([2�����ؔ�Y��)���Z	U��٦�o���\^�p��p`��&���֍�2��:3%�V����Ԥ����!!���ۈ7C�e���F�����X��e8��f1d~핥s�J�i Jd6���(��L�C~�
�N�ץE�4���H���ca�$��8~�qri?�����<̚��1��K9ylh�)�&���h����O�*d�4��Yax�MC�
�mf �q��ݩ�;r��1�Hu���#�"��Q����KY�\�}%�}��.!xt+t�~6���!��-����J���.�Ƴ3�NTA\#�f�7:�����u�J6���8��纜��!����s�&��x?afDd�TFCN�#\ْ|�{���H���|����'jMO�5�Z+1�ؿe�j�Y}e�0nW�U��Ƌ�,�$�|�>�%�>�i#�>y)jn	�&��niN��iDhRX���� G.�����@tġ�G=./EqF��g,��*��ɍ@F/1�?W)/E4y��_C�0��w[��8���9��6�|-~��Z�EOh�*䔏�.�$:3$����C�$l�0[I�E�0�iI��n��Ʈxd'	�"3�k�h��ů�v����CMV���q-3g���	wbz�A|�8aj��KbX��2�=M\!�F�.p��pjA2b�(��FH�� M�~��k��^����%JJ� eС��[�)��5(S�mS�WZJJ�8���(���N4#ޜܾ���K�<��%`����Z+��#������`��3�af�zF�N��֋��q�,�[��H�Į�����bI7䮟FH�	C;���B%�4g����61D�Ǫ�w���clG$1ʼ}����&��\��d<r�A���!,�$$�F��ɷ7�v8X��:�E��ߚ1��U�*�!����]׀&�)�y<ćP2-�i�x('�GQu�F��w&&�0ٲ �t�e�����X,mKI��M�:��������'a���J]��(�8�O�-�+�o�����Z�R�/�`>d^#6;��+�]�|O|n�`��-��Er$��J��.:+������|b񚘿J��H�f�\H���b�r�J��]g���s�7+\ΦJZ�2e�oVR����7����`���c����c��ذP���Bt�n������~��n�C��G�v�N̦2mBp-} �����Ǳ/j � ��nݍ>�J�Ϙ��Q�j�!u_v}������ ���'�סX�)ȵ�M��O�N(>��j��e&�� ��e#+�ݴa�z���g�ŗ�Ѱ7Zg��2]@Ӥ��~���vπ!Dh$�'��3#�J]g���KV�H��ã��;�V^@MW`��3�5��~�	���x+����Ճ���X���(,��!�_����b�r}��Y�mr����d��-�F:�mA�Z�p���$yo���-QӢ~�`a�+?xǟ0 ���9�5P��j���y�a?�H=n x?|3_���rb%���e���`��\�#������G�f�24�$�a�ċᾀ,��pl�Q�j���"�v3�X�	����347��W�}�ي��s[��Ԛ��;�Q�XP�T�����cs{̴y	��:jqѳ5=^�rǁ��u��/w���p�����Ȍ� Pn!Z�7���W�يE�C�bEE�Ǽ�L#G�x��.=5�0�������%�~6먇����F�a9+ݼ>\ݓ���a��@eS�����<�2�Z�����¦cĳ �����q:'0h`���$�^�/ʼ���)��P��+��\��f>��-�*����̜s�H<�����'��`��"��^�S�1N�,"W7�E���`�	��X�2�*L�a�}���F�{�}��ZVe�_u=�
�g,���0�&��=e;��◗�P�H��3|�w��\�%
�bv�`J��^���`�2�A��֚�|�P�Ա:�a�8,
�]R:���&bUab�`]�ƶO�j-�=K1F���GB�qU#<�++E�*`pV��Q�5x�#dĵkq��p[	+�/ʮC%[T�˽QB���R���@�J	�ׇA��;�E	&��j�����6��H*8��Uݳ��<S��e��7��VĶJ-Ω��Aj�@�����5Q�tB�$c^t�@�hA��n�6���+���M��fk��(�H^�5��}C�l��7�� #�8���0rd.'ZF�K"��c$�����Lb��eՄ�E�� [a�k�}�}���z�x�|¤����1{�~���g?`�8���;�u"�> �q�N�0��t^��K���	B(��V�M�pR���I;:�j$9DO� ������xT�%Io��_䰼Z�xz��������)�E� ����\B�|	��" �@ ����7o�(I��g'y��6��m�1�vPe�\)�V��M�*H�Ы��z��^{oY 4�k���>��3��eYab�c9�����N拘���b��q��J:p	���wk�ܨ1D5�kw@��(��91%�z-/��F�Xo��1�>��5���F9�Zk`o�S��+<R�"ho�	?�
7,��Y�ȁ~'u��*r��
h�T����A��������h�+�^|S�D�e�W(�t�Q�0#�`q2�c��dNx�ؾ�x:�U�H��!Xh[ޛ��)r��~�I�`��2ў��
�jE7;�~��2��$o�ްP���f�|�S��w��
� �S���*̓>~���K,��2�&F�k@L�"������6Xc����ɲ`jڙ�G�'��D����ب41"X�6=��G%	ψ��`&��̤���/�"��&��v9�`����}B/� ��yQf"��6�7�����k�yyNs�]��G�n �\Zz�xO�'�yjl���
�'jί��Ѝ�cqF�Bl�;W:�ܛ@����b���F'��A�N�CkBq��8�Qö��0�ʒ�ѭ`ʅv���5|�>=�S$g8�a�&��=��>��S��퇸�1]|��M�X���ؠI��!XV7}���;D-i.qQF����wE��k�M1�oBya��}�
�c�BN�����̏�7��S��ߏ�W���}��V�|�W� CRl�j�V��'7�x�`uI�z��4*�Q����M�Y3�*,��B��Q��`��Լ��4Zz�ۤ�ˉOD��~Gt��eK��4�t�B(����]�o�rl�D�ƫ\M d��4��hg���!�_�@� ��i����G�e�ns��Ԉ�!�r��M*��t%1����;��J�O��J�:����M�w�/u̡�
f�Řo��_Ҟ4a��ꨍ���-��g��%h敿�̬�=��E&9 �� �JX����L��m�s�Kx��=�(��F� ��B2&���9W�ί�Κ�#ƃ7�m�>'3m6P�U�15?��`$_�mP����
��g�-[�"Ttb�t���+�����"C�k�1"��Y~_�'q�丶�7����F�<uv"5F�{HMx\�/u?_�l{�8��dXUk$��KG4w�q���j_@�/n������G���炣��w>�7�1����ݐ��V�jK�ܒ��Dy��sa��^em=eI��R����!�=+����+XV��췚[��q��l[h�4�䫊,�M*�o�[e�����{�ݟ'��Ow�GPuE�-%�)�,̝��EN�̰A;?���xJ�F�\qt����ϚL �J����o��a�NG�-a��c;�6�ǻ1������-�,�뺁1�F��g����^sK,}��t����n�H)��K�����e�a-?��0P�|�d�N{ؗ��"fv�X;x'���Ό�9α_��Zv#[8�{�K��l��}�Q5�(����t*�N�#�a>3e��e�ߙ�64;6��K��Ʊﮊy�D?�Y1=��3�4�V df6�0}f�7g�Ydۛ7=<���h���a���w�:�S�B�@��p�l��q���&����*����h�����q����)��������6��(%²V2(r�8.SxЂ��4z?o�Y��p}�`E�Κ�����S����h�^��ͳ��3f:�\��BG{:�U*��{����_9ƍ�b�f�P��
ռ�`�D��ݿC��U����B���K�b�Z~Rq25��7���zF�C/d�sU|y�Iք+PHD@���f&��ۯ_�ꚒEǰ��4�?X�{z&L���1�ì0/�y��T+��;����j�KD@�څ����X
�fz��J�n)�~���=�YhG6!�(�d��]z8kz�x��.s�����.-� y�X��t�L���,���D*ϴ}�x)#4,u��(�TyQ���x��q���7����ǕE���uVNuN�X������Co��- #��#���#? �A��q�eH���Z����Z�P8aέ����2�NAs�_�j�_g;xK_���{��/����/c�ª�ݠ/5;�2X�����tߡ;�|)�N���w�S
oJwD4:�rTfN|�E��5B�WT�<ؙ������X'���ΓE��n�
i��k��#��Æ"zsw]����/�<�s� ����([����f�p�ه&g/�ȇ�A[E1�>w�[8p�}�l���3N-"y�t'߅��_��x�ܨ���M�e�i�����8�E����j��%u<�ͻ_��?���L�k�С���;�J�6/���0^����7�'~s�a��v�~x�O֤�[�GV�e�7g�^�ΛG����MᎰ��Ǆ߬�����U�%����W��o7���Pp��'w'�d�j����o%3���dl��+�3����vr�D'��Q�{��)׎q&��H|�t�7�I�.�dw���RvQmyd�p~���s_Ů���w�s�t�����]s����v�
�=�B�!St��Š��?뙴���z����i�u��d�lNM �-���T:�x��-�yBc󏞚�ޯeT=�VWUUj��?ک�5��3'f����9o�@�!�_v<4���n뜥I��g�5��B<��^l�J���j�gP*�J��^�5�!N	"���u�Ӝ����������z�w�1��e��n�E1|)�U})o�s���qZ�l4شR���d��~�/�0X��,�D�i�u��F�]�Q��F�#�YĜ�%�&�����P��O홟�����t�wt޻�f
�Ea�ofEv������T��%�c���:{���Έ8ģ[����ךª��J��rL�+�N���Z
\ԉ@�F��}��)k;b�t����wz�.�4$?)��<��ɻ����w
o>�jѹ)=&m�1�S4m��~�%@:AD,˫dc�����Zz��-��^f
�I�d�����FX�YS/!H���;eg��Ɨ���Kۃ�~B�P|݌o�2�_�lKCy���s����]��X�Z�W�����C:�t���҃�d0�
�b�.N�=�I��fzk���5��\�B4��r�8s�e,�$^����l;wYTHPtX8�CE���e����,�6n*8}뉟G�tJS�0��]�[1|T��YOu��f`�˗e
="w�e]�w_�B��5�|�v�Ts!����F����">x7��dP���PG��4�6��4+�69�'{M�s9g����݂�a���ԂN����t9-�|S��L&����ҁ��j����3�O��q�����r�)kl������-�]��J,����ٱO�I���{��p�	�$u7X�:���
�W>��m����m�"��Q���ck�a9�V��Y 6Yl�s��=~�b�a�oS}�yƪ�ƌw�Y����NU�0��5�
Pex�S�C�i��G$�����;eş2ݓW�c&���.�6k��I����s�%��z���zs��X�"�Dq�:\��(���a���3�\��0�,�:V��p7�XK�_�<��U���F"��mb�T�tT���>1>�^%*����Z0R-��a�$ �'Zn��ʏ�0c��~����uq����tܤӄ$�n�Ġ#4�oYN��H��.Ȋm!|8`��l����փB���s��'�k�5p�D1=�f����cNn����|^��G�/W�̌��r��Bu�����]'_��DjE�wH��?bg�J�%GǬ-����D#/�]�oq�hֆ��,Hƚ���՞.i���4r *R;�����.�0\�������C��˨ҋ�8�Ӱ���ؓ��3&(�ƣH*q?٦��;K�	-+v���0�~��Ȅ2���=�M�2RlB�k_���cU�mv ���h��x8��w?��"O_��6��!�[�J��Ϻ�*���O%.R}{xZO ��P�Ns�؎6�֦j��+�(����bM`Oy���>ۈ��p�����:}��|{��o�{��s�a՗�e��@���Q8֕�؝-p��%�-��46��yd�� *%��ĝF �r���=�Φp�$� �.���nХTuw$Q�uAa)ɬ�"9B���v#>�a6�ch/�)�б�#4k�nˆ�g;7 gx0��L�P�V �Ca-��G]e���>�Vy�:�p���@kP���~�,9|d8k�v�q��9����]�n���g3xdi{B�k�v�q�<�N��/D�G��߾�ΣP��Z���d�Q��$�s�b��w����@�ԇ�M����IdD�����tjR�aS�߸��>��$Z��e܃�f���e&V�#��$6\3XB����$�|����SWD!?5&f�Tġ�����	~?r�`Z:$��`k��9���h�N�,m�������L[�����1�sJ����xG���+l*�$Ԙ8L4�D4�9�"B�jj�-ְe���H�Ь���h�uL���K���Q���׎&~Ca"-%BWδ����}�շi;V������?�h����5擓G�y2�Ө��zDO�Df���k�o>l�����fs��_��a�v������� ��vRf�u:�oº��������nEJn����;�0��&c}i�{��놞�\�}�'1��������F���DFᱥ��}�"r"!L�N�o�S8����b�Vj,�z��A�+*�
�/�ɳ9��.:��$��Ȣz���G**  ����K;���Byr�ۋ�� �Z�ϕ]c�6�y������N��� $t�wV�=f�Iė�h}[*���\t�2�禙+7�A]Y�5l��M�onZE�#� �G�9'cC�
�j�3��!%`<��`C�dJ�4x�gv��/C���u��)"��/A#%wOZwy٧(�i4�bY��-?!�٪���ic/(���$�vP�N��h���If��i75%@���	0%ċ�z���1,@]�t���E:pk��%:��^w�z|�d\s�X����]8�7���z:� ��2&e�V7q���q��o�;㚱�1�<�@�b�TTۏd��&<���G��4�
����(%�`[�6c]s�}H��ج�̮ϕ9�d_�s _/�)��Z`�ۇg���(�����$/	 �w�5R��4E���J�D����{����3�<�����(��(�/.�2�cU��,U+Ԉ��p�l�%�"̍*�H<�;��o��mhFKF/qƵ[��4;�0���˨��ɞ�Uz��`>ߴ#h �����'݂����0���ml?V�"cd&��d���w9ixeD@ w*sAn���6�Hr��Kf�kJ%ώcHHHp~�8��/"qԗ��I4�To*���=�y�X#�����O���)���ď&���S�f�Pg��LV�3�(��?h%Rm̍��>��f>j���t��:�w������S͂@��:����'���0�e��PM�B�b�D�݈�2�i�����t��M�NW|�l�c)kQ|hBΰj=�s�`��<w�X�C|}�h��̂4�5J߇7J+:,�q�vPp\�o3h��ό���D�rN�jUp��3HT���"X�S�j�����:�;N]��V2D�b��@��>�)�8Zo����D�M�8θ�҉r��2rz��<�ޤQo�⒕�]����kc2��&e�F�0�،g3�A�5nޣC�$8;���ѻ��-u �c��hE7HعW��������n�c��h�����dϣ�̍����nc!�8��S1�O�.���P��ZP�� �X �$1���8�a���Uq;lO]׺�r�[#����DS�Rt��,�7�Q&p���mbU�8{>���İ�r�L�%�A8�S�����{��@�5�e�x z9���B�j��>{s\y� ���
ehYӨ��O+�̳UM�����m@�Ҋғ�ŕx�j�}<j��myHz�o6}�_�YI����O�F���W���'{� ө�M�o:�8��J�LY�[�B�y/8�XU�����%��g!�q�o��3��U��?5��z	܏��R+&���_����~�ű.��o'A����%�����PD۽A�(��`�|��Q"*���+��;�&cq/;�4��P��I�A
�bm3�T"(�'��s���'^X�~�M5n������x��8s��]4_$0���0��r6��?F���D2f��LyXG���凌��	�0��$&8L�2�VM�UF� ȉ��Q�)�.����Wdզ��҅T����"���R��l�Ȩ���b�pw��נ�6��I-��94̴j:��x��'��`�Q��PQM��xCɆ�
��d��-��+��J��4P�>����=s:J���o��ݦ�$K���c�2w~� K�=8`�~޳;6vW��))��U�<�vxdmd!��ϟ��z!�BA�H��&� %�y�� �%�
O]i�'2���>aq��@�h@~[�7��=P���h��83��֏��KF��՗	�a�`�S�xqi�F׹���V5D��)���NI/���vQj��/2X��7��Qz����y��#���X�p��T%���>�
P�i׺m��C�ޖ�t~��m Td�ƴyP����X���,l�����)�T�+m',k#A���::VR|m1ʁ/�77ȶBW^�Ԫ'iO&d�G�H�aA�}�S&�}p�2,�g���԰{���z�Ȩ"��tZQQ�*��[��E(��8�dC�Hܕ���,�[���n�<�eNR�hR�4���ݲ̑�7aОͶ&�4a�󬑺 ��1Q����k}�k�-�����6��ZUI�U~�?�_�7���vGjj�t�'쬹�IɎ!`�'_�VҊ�CH�w0o��M�s��J���i�g������$Exq��k�ϧK�����ά9�Q�0IKN�������K�3%�;p���b�(�E%Y�](��`�)W�O�K�O0Q�s����>@r�0	�ҚC7�3$�Z���e�*�����
�Xj��_Un6�J1�!�^6�Q��%3��Ib��<>bg��W�PmD����@��<��VN�7Z����M�	�"a#��q��q��Y�rm�Q7��$�IB��$� �ի�9SV�J���$�%W�&�¥i靉%��`�A�&$9EfI�@Q���葬�*�;�mJ
�9�_���K�W����`Z3�&��sw���]7�Vj��*]����"�1�	0��������T4�c�����j��x�[¸�\�������̽ H:��VV���$�_>$<
߅�_I�k|���N�T>73e��fw#s��	=a���mg��ӗN�u��.�2��Y��*���Z��KT��]�E�;d}ҿJӜ�L��#�ђ�Tn���|'��r4�`)�ST)O�ϳ��=���aq�;��
R��9�B��$^��W����H-h[�rZ
�s�O>����t�Ǵ�4O_T�^UF\��25�0K��#V�fB� ��'bl��g���]ͷg���_Q������'��Wi�B��fӧ/$*�v?Qz��~��g��z�W�%��J�3����W�꺅��l���W�D XbZ���q�_�y�D�}_��Fr�W��<V'�h0��$�`��5��2�k�UQO����Z걜)�[A��InmiB�A���gmP�-v}��E�>�=ߜh��Ј2�&�DJ��2�Z���o���a}��4a��8�B �x2f���
'��Ka�+���Ԗ|cGɇ���pZ�g8#��U��-����,�۝|����x<��}�c���rY��x^��>Դ��gW�໋��\n�����{�qXdhc]�+�.�3��g{G[0ؓ�.&�})6��[ԫD�ڿ6 ${�G��&$E&9�y���:���۩�?��t]�gz�� u�H���Ģ~F�\L��t���c��ү��z�����c"V�3��v������K%ݹ��y����՛�	nI��Z�̯+�n�~�F��vY�b�_~]kvM��v�?lw��y%Xy�h�$�+�/���}�du��	��˱O��7�	���>E^i �<`��4�o�O�Ǟa�\�/E2�]_�q��.�`�#4�&�~��u۞o��~;��42����ӕ��lNl�6��*�nC��y���|�>]����O�]���G�
C7��\�з���T.C|G|���W���W3�/ë˿�H�_��YtϿ���5�Z�z[-�y�Q�F��c��p\�}����2�(l��[f�O?�*��kzu��(�ԇ%biJf��i����?�欎�sLg�b��r�Hk�4F�*&=�~S���U�fڒ����W��7}*5wK?�$��6�"�x�>7I_���}Â>i��j�H���zm��6����t�����O��9|)�m?�B�u��fٌ�^�Hq=����P��`��Tg/��6�
��Q�:����q�z�O�Kq��%_����:w���m�
�L�L&��<��'f��Zr�#����߸�}�R�Mʃ<�)�Y[љy�f=���E�"�b|������l��Jz.�t�k�m�����F�X�YgR�i�f�_�(;�����/+��j�O��H�:Z�`�i�>����l3'���O�p�r��x1���듺Vľӭ���W.�l��N���<�T_�ebſ�%�Kݪ�ӟ�:?[�����y���q���o4��#��;:�]%�v͙������s�WKN^������{�3i�_�i�G��ŏ��B�+.���C�\ѽ��{��������"U��Q��?����*�0y�jox���mi�s�zi���[(m�q7Ι?�ྜ�/]�����n,'��c&]+���*��w�2�&.�����.p���܀����I����_����@7���܍d�����
� k$ʴ����/ٿ��<�~�ߊ��;�b��q�(�7{����i��*�RP����DJ|�@6�ܮŶ��bui))���S��;��^��p�x�&M�Ih�p�n��.��]�c�����������->��=<�����{�֢0Ԯ����wx�+�_r�9�5�x�>��ޖ�
x�N��HoO�it��4��s����;,�ly�W	�	wa I����r$H�(��.@�р�a %��(��h G�$��9M�����y�}�N��ު:���:@T�*usO�~�ѵ�,�?��*;�*[x �o�� T6�0Pí� ��������;U��ZÜ�[�,��:��׉.��G�C���Do��Q�G�����R��q�tt� x�;�Pb���\F�B�L��s�;� ��]o^����|�d�c�L���g��'L���� 	 ��:o�^�3넞�����yUN	�Yy�� hE���ĺ|}�ɺ�;3H�roqۅ��bA�)c�yt�.-N;�P�U��[G��kfg��r�ׯ~N'ܡ�����
(�q`��K�2�':��=���p'@��+Z�)f9��Cu$�aQ������?9;=lIa��� ����{RӜ�3)���!����ˬ��"��9)֑�}��I�2Ȇf̭Q)��S�e���[�2+g�W�r�����n|/���v������_��x;�[A�����2dnb�<�a*�<G*`���Э|�F��L
���Tj$�)1����S_�����c7қ���aD�f���]�U�면țh�	���r،�
�����@9b�=2~�4D��j�Qvc!^��N��7�-fh�@5��l��.�b�ܺwRA6�獼-����|Cq��V�e���֒����$1� ��h��w�H��)�%�@�^B(4����k����;�7��"��DK�7��Á���*;~�#.�7����������s[�:Ve�Pn��F~�cH�����
>2�H�n 
��|����ϭ�pS�+���:�Jd��;3}�.M�� }�!q� N�6���w�*�;-_x��{Z���1����gЧۍ�i(�cZ��mc�;M���3�o��ꙋWu%a�g'8?֬y�\{~��lJ�Qi��	�(�/�=N�q��J�/�\�����Y�$�{���<O�Y�*�����.A;��Ytz���9�Kq������o'�����A���sO�$�[O�b���m`���?hTO���P/�S��[����[�ͪJA�*?�rP��T�'5���NtD����w����?�L��e�b+�<��V��дqr	&��r#�C0��3��i�6k����6�ͭ���Ke��.\H�jy;Y	��&p�G�}r�JjB��{����I	�������(V2��A��k�n�s�9��V>��M��ʴ���Iھ�Fa�;��	��6�i�Ň�1����5p�����z��ey�\@��M��q-J�y(�F��c���^a7Z���g��\�ŷl�w>z^�vr(�I0d6=->g�P���n�At.dSұ�GW��=�A̒���U�t��v2ׂb�o�0���?M
�mT��r���~�R�>�!��I+������j�ZY.Vw�Z�h`.��JS۹	�����+�s��]��t+痂Ÿ����\���#%39s0W���}����� G� eٌɱS��
6 D�ӽ?��C�F�tlb�.%B�E���jP��a-��
`����v��v��wʤ\r��/+���R؋��.΍5��c���c�|5�5;�6��K�� �{���!`b8�A��	ŗqc�W�!��3���O+��$Y��o�,~j�a��d�	�'��悩�t�nČ�~�Hu\c�;8��79� ��xU͸�&�g�Ip�I�Ӕ�Hv���m���4�Od�����Y&%�D4�U�*�h��h��z��<��c�hDX ��4.z��(��&�9���$���N_?�� �<kg�_�v�u4��h��r����\��u(d�2{�����;�ݭ� %�ƋAs��;��*�L2�~�5�r2���B��S;�}��0��<�yğ5�z�i��%�)Y.�s�Lh�PxN��8.��_�`�A
i�ދ�����X���o߄Mas��������L�[ɠE�wD�"��5��;x%��v�k`.�d��<�F��"q���2�V�S)��}`F��� �}��:�T����e�-��s>�Y|�̷��`=�Y�7.�6�} Ngf���0M��t�w�t0X��&�ϾZ)�"Ϛ/R�R�z:ő&���-1�Á��r�F��[-�o%���+��ߠ�`s4[������7Szۼ6��љU��Q���+�C�D"�N�Z�h������f(18m���:[��?�<�j.� ec����|P�(a�(���J
(��	��tC�3�[���6S��m3+�ZB��	�A�/Ո���*�#U�-:2l�-���g�qb��C�
tR��E�҄僁�ABU|Z│��i�b�D�����m�+ Y���.}RJ�x>����z�����Rb�4DI�F���?��l��:���`��y�6������8�����7��.�iWwق����ގ޸�K|����ދP��f� ��	Ɉg�K	��F�N�����FU�dYQ�q ��0��?�ѐ�q���<��r�CY3�K#v��S�6(�k2��&���:��F����o��s:ڡ�[a����m�;��rPUJ�mZ2�����m*��.�g>�y���9���dV�թ�����F���kxd.𐝯��G��o�V�7���H����z��="m�W���O��Ok�t��1`��Xs�6T{� �[�X�}]��t��F�s-"��DZ[��8i�>��q�nn|�;(�i!�5�r�n|�ج�TX^�6\��]<��(~U��%��c���LR�Y��MU���ٗ��5zv"z��?ƪڃ�� �~����һ\7�i%��'Ui'���m�iH�:�g)�����Y���7�# ������=�U��ϋ͝$\�^���ެx�گ���"�ZQ��bk�>�r�����@��6���!��3�iÊs�X(RRU��^|�"�=���!we�9�v������t.�xk��bk�Q�z�*?���"�Z��¢*|lE|ޓ_���ά��|���_��QJ�yJ�:׭MM��,�в���"��t�� �n��(i���֋j�b�CA��,I���Vy�A��|i�ib-	��KF>;)w.��ֶ�&��H�4?sۛ�$�Ȩ�����~�wP��?�N)���S�Tbŀ*���e�=g�&LISp�CQ 'ը���j�6��~���/[�������X�=���.q̅�$�>�����ԥ��
vw]����0_�+M:�$���x�t�g)-��c���Z\�1m�[ރ\9�
�h����7����Ag��r��mΨ+}�Y�s��J���Ѥ�	��8L�f�5�a�Y@����ǅ;���hc>Ș22-Ͱ�Z�9�b�u+f<��8 �|#��
[��-�{�h�z�ɒ{��o
�Q����`�V����?y�ކC�v�9?��&� ���p��
�i�7	m\�Ǒ<8���#t���<y�`u�I������8�(����Ҵe?���Y�譣,�)q�C�Zc��"��W����Z�A�A�E���a�K:S��CBd���	�Yo��w4�F��8	���|A���#o�wc�ޡ"��� 4���}JQ�������W|�Z�I���`�^/������za��k(��<][U?H�:�5`��K��������C@b�AZ�˰Lǭ�#�?�:+>pNj�?.��������S����-��f�99��aNK������Jb]��@J���y���\ ��[�a�ʣJGA^�Np3�G
oZ�#��/�3�,��XcF}�Tӕ�z
t�u�_O��Om������p�W;�O���Cd;SR8�[�~Y6BW
AZ-����5���iJ�M����h�����[|&.[��}���Ե+)E���{uh���4��MVJq�W,W�l�x=w���/���F�j�E���+�HH�QT�9`un\��{9Zcjm�]W ��ӗ0sQ5�-97�,
 F�k�l\��=U�"&P�'@�_��8郌���2�䐌x�|�6c6���ˁ�����{�KS	qQ�����t��('�T^P0�°S.T��&"h�55>ϡ˴�Ѳ��j��j+�|��P'WQ��.��O97��V��B �W ��_��/rU�G��2���3�,ɝY������
��)�bNtf�m���\�b��;Ԭ�IU q 4�di��񦣮�����Pv����EF�Y���ncb���څ�=]��0��]������FTN&���>�+�c��7r�TӾc�R�I÷�⛔o��͡�w��0��56��Mb[��i�o��,�$�3kȟY�^��[D뙔��=��ː֩�<�)6*���q��7�f7㮕��X�NxZ�}��������I��[S��+<3�z���La�x��&�wy촻�V�K|�!)����A�A�FQп�}�u	���V�y&��� AbS�y`���$���z� �P{����ܛ�O�C`�G�IW^Ć����C�E����V
�Ӻa��$�&���Ȳ�~%� z@,������(��G�z�I�S[Y&��.w�7�$���~�jY�=���t��h �EP|�g�6�5
C�#�B�g۾?12}����K �*b��9�����]:�ty��"��{�W�l�\b.�l��Z/�Y5��Ż"jf.w�����C'���靕h���)��蝄�Ût�+�z�D;�(��˛�j�X���Ȝ���c���
��|Q�t.�/���]����9
��I��lX$p#��l��:�f���*ķ�0���\�ֶ1����xT���c�t��(����Ǒ�_6����JUwz"U�g�ޞ"�r<B:*���b�Ý~�7V�)]U����ƏF��#X�b&&-`Z�Š�����克�p�2[���j�����`�LrMԲ��+/O6'���t�.9�A�] ����2Uv>���n;���XI�h[E�_7<��	���$̣T~	PF��"�Pv�� @�C#���-��l�A>�`m4b|��I��T�ZBKH���E��<s�pʷ�+�uLfg
�hz}�G�5C1�Cn��9?���N�m���$�n���ST<�̍j�!ΗsR�����H�t� ��Xnsb�{��BPyԾ��le�;�0H���p�g�T���>te �.TauδxFR��gq��X��b|N���**e捊����E�b��4F]:Ɨ7�tk�Q����r>��Ƕ�'B� %:��_M�Y,=���+�yWE�j�m5��<B(��K{��	u�2���Cb�<�QJ`�M  l��e����x��.��m���K)��˭a�F���}ݵ?�}g߽������'��ӊ�K�f����/�"�A��V�����ZϬ|��y3�T9�;Q[WY�v��V[P��Q�9}�?��tc-���I�jhlUFWڱ�|��GWP �turZ�b�+@e�����#�tn%��Q0�H$�#W�n��O�MhBH@��a�]"�ߒ���L2��㝏2�އ�VqS��1�EaŘ�SA�][�Fy�|$����B�h�Y�a��� �qk�q�ڣV�w���g�@�s�ܪ��3�N�~��4�	�k`e&�j���y�%P��
�r�e��u	����%�ǩM'T���ŌV���xz�ʅ5�L�*��ހ�tCVG�t3O��N��ZOb1Te�k5&�3����G���of��`<i �-.�9�mk�B�r ����
�U$��?8��ip�"���N��R�*V�ھ5�k���wS6>�-�k����3Qk\s4Y�/�a[W��1z��M�
w�.�{[��>�<�L���9��Z�G>{�������̇�&��Ε��߅� $��Kj6z��x�LT�,vd�nG��T�弾�-���O�k��.�n}PA�-Y��{;�V
�[xԡЎj�ۿ�(�݊ �]^���Ox�Z�44#�ё��Trb%̟�ڣ���?�k��k�+���T�;���F/	-���o�kY)w�z[^Q��HS|o����|E=j � �2(Ot�la�X�*�Q�K�!*�+���ՊX	pʢ
_ N^�9$=1O�`��l����tZ�U(Z���a��)�<}��z�ud�34FK�f�Ǜ�:��͍�`��x:B1w��Mq�K�mm����V ���<�2�?%����\�����<Z���#��'%�A��5P�o������/�BW���p���9����c)��A���咼D��皩Ϗ:ax�F����2_����3��I4�yi�rP��OpblW��/�p�|�(E��1�`�S�Nv'�g�EZ)��j2޼
�%@��sR�*��6�j��)t�A�h���;��f� Qy�N��z�i<'ds$���8������p4�hi܉ M��[RC���(�!�G��<��zƢ+m.�×�MN3�������z��Z�:��)/�GL8׺��\��{��m_j��c
�]3�S�}M@#��M�oޙn����~5AO�Qs����[j54eՕ#��+M�x���Dᕝz�|(�����Ö籧��
����}�����
j_.�_����WS�b��6ɵ���g��Q�E��΂MT	�]z`�@�>���F��#L&��BBg�V�P�׀TF-ע�/ݶ^xE���&j���~�����z"Tw������ m�x,��<���agN}k'�s~I�kc����2tŭ$���<,@�^4X��gsm��ڴ���6ir2Ci(�cy�]Y=���4,59M�s!M&�u�j��į�"e�˒��E�s�y3z��[g����JW�f�<�$Ԋ�P�O"����i �g�����d7�=G@�3�S��8-*��nQ㓔��j���H.���E�'cs�a�1��z�	%��:N�@7|����S���qP)2"N	۰��'���T+���D��P�W������j�!���V�#m��P��.i���Y����)����]�e����2'/�2QX���uTr�^�B_���l���|CGZ�o���(���9�t��4ڌ��KkA�0�\:��J�5�[����(�2�R��g�����k��we)OH̉Z�eT5n�V����\���܀����&�5�`y ����k�� ���/uG�l_�$޿ڙt؄}#tk��3�JFX�/�������Hxx83���&��,��9�"@c��đ�#�QCPT@��ϋO
���[@S�����g��r�
�:M���_Vv�* �q-U�hk��U���}U�����:�*����'��JrkG�),����p���OPHXC�� ��?��?�&>d<+}Ғ��,�r�}N����������$hz(��d�8�a��p9����3;4j{�l�N؄N�� "��[���n�6`�nV�����uq�k�����I�j�ZOc^Г+z�y�=w�خ�63/>�DN~@*���0��
�b>�:��i����/#o�yJ�ƻ���X�R
s�)�}a��Wl�?o��ZF��7=��E����T���
��!���ܾ̩���;~��<Q Ϭ�������B���cdq3f#_��yt�q-�A�3�[�� &�@,���Е��釾���<+�4�0F��ǤrZ׉'j{�|�6˖Nz3��;Y�ؤ�6���~�x�*<+1�>kW}�x���� ��;��* �QZ��!�
�ퟎAVg�}?�_�3}��}�o�k,k�����:���<�6�|y���^�D�G���i!zWv:����}Igޥ��޻��߻Ln�;V%�AW6M�=P�T��e1o�r�t�H�0���F˩��8�ƞ���}e���l�es`�����N4~"��~D3�p����i�r����Wֻe I;ɛ#�?�3h���`��B�<��xG靾�Y��i��S���t������������Ç��#��on\۸=ul�
���V�^yn�Υ��N�E�<�jN(}�����Z��|#�Iۉ��G�d�`P�|ƣKf��&&��m,E9 ���q�s�i�OB���})�f����ܓ�Y��¦~� �L���=kZdk��I̾E"p)�G&Eg�/u�Dr�r��o�2~�$���k�SY�,�X?��s<�����T�:�S9����~hzϖ��/t�2T�0��H0)�r<`���BT7���΄-J~h/���|Z��)X:��)� F~s��Q?� �j�E��pg�>\V������f�$�-"�AWj��ܒg{�5:!�굺CS����@�k�B{}���ͧ��uh]Do����;��	���[�k��꺱����,3O�U�y���Qh��p�"��bOvl@4��U�����^+MܾS���`8��L�NeI��D�&~!�ɺ"�_05��GcC���/�L��&J�~�����-?�S�o>���8|��] ������k+N��w0�׷�g��j�f�90(�:�0��T�Iқ�}:�lP���B4�_�wh�g�����Xv��� �Sw�8P���ߴ���}�����H�L�\)�O�Õ%���?��-�,���LH����ɥ��?h>��KxWc=���-����|�h�����c�z��X��W'�C��G\�!)kwFg4ɻ-є�,��-KQ�o��$�ۺd����{�`�όv����ȃ(1h��ӿ�"(&�7$����YH��=	�&�Z�k{Km=�ki�A�I�nY�y'gﲵ��P�.Y:�r�(C73�2V�(��Y��6Ֆ���M�) @BC�l�fySO����R��L�
w\�P�x���j>�ܫ�� �Su��*�/��ˡ�|�ȧx:��_�v��������g �}?��$*̽���df�&�p�fk���1.���ߡ��g���e.��-�'�F�e��xa�U G�&��{��e�Y��#O�F�����+?��l�x�ч�P|�O[~iWmj�d1�X
����:d��Y�W��#0�����u��}��������j�xZZ���a��LL���x�����/o�5� �N��sa#��濥} ���b;iM��2Y|�j�h9��ՠ�;�v7����9���F�ŋ�FP�ňM�"�X`��J�v��eh���E���2N��oޞ���|���l5�s�e̾�9�N�>~l����{�Sq��ktT�ڲ]�O�_�-uXw@Eҝ�n{'�
�;A�����sE�V
�ei0i��*��1䶢�cxM����E�x�* q���l"��Sϒ6�!�v~�d�\kҗ��F�Y@;L�.�����\"k獊�����o͕@�����]aVi��Ȱ%}P�:��v��#s�ҵ���%�{So;D�I:���W�b�M�
�@��� o� (��STF�s�#U/㺸g�6��n�B�}>a�����tF�Ү���"law6��Z���q �t�m���D0C�^�� �	��Լc= VF�D'c���?:b�ݓ�FU���8}H �;A'�	c��1|t 5VȔ�d��:�j� MTj�u*�qu��V�z�5sU%Ū�>�f�`����-g��\1T�F��K����{Yk˦E3y���@��V�V^XE�̓xw��ؠo����qH�"�����1�X#��Bȕ���?'��,%'&�,�e�S �MN��S�5�B2��Y$[��ϱ����������fpʿ��v�~��� ����h2UV���z��UQ�u#Y�k5��4yи �U�վ�8�R|U1� R�իrn�3v��qq��#���Q)+<�P�O�Ԡl@��׊��$X����}�
�*�X�J�+��;7�!�W��r����|��?wd�:��XB���X=� �Y��׵��EUW�NQ���\TX{`���ʺ��3*���v��j-_�Y�^���՘�|���e�<=�$�x��F�O7�͎'��:}�kE� �Ӭ�J�_�+�G����>���@�V;��� ��	e�k���PD��}�{�`K�%Co���N�=�YZ���E/��PJ���3�S���D�DF*|� �ל�u�����At������pb�u�T�s Fݲ�T���躴t�z��R�P���o:�����`�i�Ykؓ�S���x�L�����Z�2�f7J+��i�#S䷎�&��ǃ{ZP�L� ��$=��S���J�wc��{,�N�D]I����n�p��Ϋ���m<Vf��/^4��C<$�NR����i2b��J�� ��[J*��l�@���@�S����f)�ߒ�H.T��j: �f۾:�g���U�|e����:��瞾���e�%���ST��ݞ>�ڝ��?���y�ם��;a��������_�P3]?4T �8����OvC��R%�yr����U���x*�<�������!�,����m�,ѓ����d�[��.k5��J�/$�]��Ld|Ʋ���F! #	�����.�rφ��"�ӕsd㻟�j�k�N��tg�j�=M{�kS�޻���"�R��.�;'F�Ā�t�1VUKƥe��k�� `��W���0i��b$�nYZ��_���{ s�=�Ǿ�E�d�/�4��V=� �35��Rx����e�EȈ��(ŗަJS?f����~������_� .̛\�j���#d�t=�t@"���dO|TC�T]�b�"Kg�5��ŏ{4c�p���mb�;0Y�n҇v��JS+5�Ӽ�>k	���@���V)�� Y�c�'�Fl�I�S��07��1;�!#���~�'����FxB2�~��|~�����/�#	o��н@ad;�7K���?$��3�������;ܾ۠ ����a̾�F��P6�}�v�&
�7�mZ^ϻ�I��H�'!�3��S�O����gR`���E�9�?�A�"4�O��Gn������2LGC�5�n� ����fw���2�Q��"r.����Y�x��rVCr��(v1��&��H3°'�~�-�g;r��8�_ȕ���ڸ�Y�G�����bc�ul6S��l�:�h���~b���Ъ� )_v,��s4�S�� ���(G[IP%�|R�H��W���C+��f �Z��݋}t��!P���ꇹ�����x��@�˚�d{��z>�Ĵ����T�9�VL�Xp��+3�~����L�F����0�~l�G���� $��:��5��[�ڙ��%��>�1�ꜯ\x�hp�8u�F���R�1��͘�Ud�r
����𤃊R��s��ks0��%�6���p�L����d��CNU$��ڙiT�P������)�k�ݫ�ɖg'��8
	9��Sm�3�Ͻ&�+h�rL~�T�W�M���/�c�A12�%�!�U�s~��Nߢ�u,��"�>�Ƅ�h��ߖ۔�I`�؀��[�q�����Dm�r,��g�� @��W]*+�s;�����/�9ܲ��qI��k?{���A('I��u�_~[>�n��jP�}d��KP�62����8I�'Ȓņ�lɛ���y�AH�;ߜ1������F9��N�\������P���^7�}��-�p����4�jD�zM�A��A���|��c��d��U�C2c�4�CU3�y˵���.I��Ԇ	aJys��~�ct�F�R%�]&����)���Zo�5Kn�������L��z���3���מ�'�M\_&�.z\��)��%siÕNUc�d#�yS�Ut/E �ۗ�k�d�%��@4��X�i=��$�x��8E�*�$�ק���T�춄r*H&�v���l�&�?���Y���?��ťC��7�:Y�W�b��S�=��7�AO
�z�ZMƋj�����wܝE��1ݤӏ���\�ƾ�'GEJ���^��?�2���c`{P��ŧk�mh\�*�����1���ϛϜp-��_/���a�e�{7�5dc:dF
��&JiL�>�+<F`�|�F�;^�5Ӱ�a�!m����0�%h]�B9�Y|��w�TY2�27����"���Vf;���,��ǡ�f0��luhۍ�kXǀ�j&_��CC������g���E���$�8��KM��;6E��Ӏg�C��p1Z!�l��]���4�~.@����~�4�	�%�3}�h��aas���Ճq�u�x�U�6�N5q)��������,'N�rAG�=3�}K�ouQ���ں�0������n�v��+��h(8�+3�i�cjv�_��mȭ���LhL�6}��Nl��me��A�H������
Ŧ�]��­2ܪ��3Aˆ^�%����n<��F
�6w��F9�;Ц�����!�z����x�t�:�=G&>�,N������o�L��w�%��OAx��S�+�/��a���x	^7��t(W�k�_N`[<{���.w�ѥ��0�'�kᆬ�>Կ�'��z1�g��C= Pc��s��^���6GT�C���緖�۶&�v2�-%T6��y{A#^p���� �.��GU3�=��z��%l�Y�6[�h�f|�}׌i�B�^q�����,}�yB��G�mi�D��"����3\��><.�(-

)}mkn�]WD+��;6v�C�=�C���G�t:��& �ڝQ�`�����bgP)�_$.�n�-�;�ۗ�?��g�`g-�ץ���չ�\�{�Yit�a�Rn\ PX��9v�M��W.p`��-�2��C��a|m����2�*8P��,��N��s5�Y�Y��4��G헻 	OgI�T�#8�d��,`>mhY��; ���$�#����.��*���i��f�5������kT]k>JV�h��3���	 S��Y�{^�
��}��:tsm��ͤ8�0=f?C���n�L
0BǢ:Ty�b]:�X�0���CxZ��>{��%�vvܧ�s SŞs����)�!���y-�x�Uq���C�}O+s�':�t��w8J?��.�*.��Fu=tMM�r�yC�p�*С��"�(�B)O�{�b�߇o9�]�6z�]�� �N ������OA)��:9��e̺�"6a#@���^U��&ɛ7����=���,mk	HU	�u|�H-'��'uac?�D6(My�2�v�����<4.'8��, �Qm�u�h�� 8<u&�r1�_��������Y���U�農X͢�����=��A��z��6��<n����f 	p�� ��L��N��D	������i]48�C�]eh?�]_�uTi�X�����_�wE�j�}tm˜=���&�-�o7�`�AOE�T��k����h�	�~�}���`AO�h�꺁��S�f�֒ �����݄>tI%j���s�i[�Y�铷q	�%�U#��������.����ã��[W��l���@�
��t|B#�L���w���,���"\��]�?e�*'��޾�.����x>���p��]'6�3�#�z�
iA�;�Gχ;0�4��t@��|�]{zs1Vg)z���xق�X4G%�(��B\�#��q32g�C��Aͻy5���m#��BL��4t��?j*�%�	w`^d=F�XY�����m>�� �4ӊԸ�؆Ǐk{$����D�����Ro�NS��:RO]ݫt�����@5��h��)2��  ���jv3�������]�U#�k[�x� ��.za�E��ѣ�q�T3�A��^%�*(�;���vD�o��X�eI�ɪ� �tWQl����Zw�R�Py�%hQ�Ovs�ݠA>�K�P=�{�+{��Ɔ���۲���$ ��9���A�Ჷ�����	z�pdH�v�C����OǯD��=����Z��� >�\"\��0�X��"d2��*=�򫸂��ZM��2��^.�������TR� xI�ŗT����T���>���	��~����)�|��Ho9�4v�WW������T���(��z�\�����K��{�B �V�����.�j��B����JM	��<D9{���ă�b���Ϋ�?�s�7@��f;3&�OW�8�uJE	�Ԣ���ro�a��J��h��+�a-���o9e,\VOu�^�"�Ǿ��1��,�VW���ۃ���8�U����7��_�k�qޭq�ؘ�w�2�jzxh �v9�9��dǚ"[M�[�<0p�^��^w�������?��v�`�9R�?Z��Z��bC4��+���������S�F������K�9�cɀff^+"]��Ž5	���D3���c������¸L�u�/��E��!M�W���W	��_w�{�ǔ1$:�� ���k_x��v�4�8�v�ȅh9�n���������m]�z���Ɠ�ڋ��-ZI��L���T����L�1�1sk�W&�U������+��G+�q����1�B�N�ӵ�H�˜��Xt	�.@�]�4�2<J��Ƈ�l���U ��o�l{�?t��o�aW������?"��;Q1�Yx���� �$�FM�E�1:��
��S�� >�D��t�E{/~���.I'�C����j���'������\��]�"��!�A�V�M���[Um��5@$��u[a�1�j����e^-�,4!��1N#<���\C	���.���|]���fC�I^0���.��}���/g䪱%.U��Q�p��v���V.�:��:��J,ݣEn��6��}/5 uN�7rW�.�"��z��M�����ޅ|f�>XJ]��2�s���c�Cpo��2��6����>I���>�|�;�#zR���X�K����'$������1�B��$ŵ�&��3t��(�K�8S���q�������ޅ�ܕ��c�T��8B?̾Y��y�{���f|�,z}��8��M�"��Eq�>ݞ��z�~�gh�v���ͼ-tF�ZD�t�n
�g�$��U���c���Gy�l�zӢ�`��t�w7:�r{k ��8��W��>�s2����9h����%���M�ъ��F_��m$L��-�e˳�����z)��H��Q\A\��,�g?ǜ�7�i��s�(�etܒ�5�����)���l��F�DC5�{}��������1,�J��2���RG)j݌+x�F�0C�8;�)��+xn��p��(�Y��*��3x��,�]��A�'흝����O���(s��¿OV�W|�x�&��A.��ˡ��v?�1	7��s���'Q	wc=��LN��_���B�}�r�g�2Sz"a��͠��<�3Q�4[E�d3�hk��osO��Ϋ�A��ߓyQ1sx��~)z�������w�Y��ȧ���H���?tt�/@�(�@�oekH��N�`�4�4��
�Y
��;(g�O�Sy���j�����ST�!h���\	��H��gv�C���/��ǧL��#\A<	 ��Q9��%�d1�7 �%�wJyz��`�E|�o�� h����,��C�?1{Pb��
i�d��po�~���p; �s~��z�]\W� �]��owe�bmf��j��H��u�tu��X�ZҶ�Ƥ�Y0�Nj �]/T��}���`(G���C�_L�Ŀ�A���}B�T�]�Ʌ+Pl��lx��$��L�`�.fS1�^.��Ό�?�̍ρG\�^L��K==o4+(��W�`�]e�?��� � �'���\n=Xu��WO�M����(��`B��ms�!a�����a���GU�d]H�?�xk������7޹�o�6Mt���h��W��Z�e�/�7���v��&�n�&�£;4�sR�� �� �Z�Z4�:3�{��I������i�p"���c�# Z��W���9��P��D	�Z5�>)�1j�R�o��_�mi�>V�T�IJO�����o;���_�8��9�*�;�J���?��#�I�Yx�|ޠ��aqU�e�Qv���Zq �����0�Uz<�a2�j7��R��*~V�.��@�se�|J�5*����}*|��x�����'�R����ePs��̌���ypPo2����uj47+�#� �Ճ.'oG����~E���K����x{���(�L�9y��3 �ܾ��e���g��+>��l��m�[��U�����/bf��R���P�yI��1v�򵰏V�/1�v�slDB8�C��:�j�]*Ǜ�q�pK'z�҇�r�k��䵇�}ȟc)W��;��i缍[�l1�NG0��K��LF�[��pxi8���eEK;[���� �Jq{}�j�Ja����Ըt/&/�);��[	��-7��烓��@�G�G��j��`@�J�z'$M*d��YBW���߉���*���a�'�D��_�k���D'�h����ݨ;�����b�2�РNWp��,5�o�1՛}B({Ӿ��l����D��e�ш<|
�V�8@=yfk��$�'�S��
'�Y��WJ��s��P���jo���*��i��@r:�Ќ��O�<��t��� w��8vQ�X�4�� @�N���1�ZG�T���#��j���p-#O�[�q�I�3$�*�D�KuS��;qU�%��6�	 Vh�������U�.�R�`Kv��ҵ�#��^>#]:W�F�E�������b���0���x�Zw�oǋ�Wh�ӻhx����o F�s��H�����,��"�=ZwKR��C�\v%��� Y"8��-����M�E�ȾN6��E�T�2�I--�Dm�"s�*soЩYe������#�, �����Y������諫�ρ�-�Z�|�2�26*[X��5Y���@R�5�v֝��0���vj�h��eZAL��T�5�NRsZ����U�����1���%@��ꐹIe^Vr�+}W@�G�nV	.�NbwV]Ѭ�'e�=��  �$:���5~��7�LŬ��1"f ��y���h][;��w`G�>�� ��v�x�Y�d@�8r�H!��7��`}'��5s�g�;�q?��l�)��h���׊����7��W��ʷ�J��
�n%�1/�o��1q��[�����]W��v��M�{��O�ς`t�P�3����?�����tGP���'��rxz��o㥝���bx����x��|Q��M3y�� ��>��� o�?i?����C������ �^f�m��N�*�H6�_�0����,��2�H�-M��J�~A�\�M#�6z�!����,��?�ॹ�0�m0(@�Ö���{҆�E��2�k� a ׯE�0�����oA7����1��P)�&�&/vڰR���@�4L.���pW��+o��Q�	�=��Qu2�C�8������ȩ����l	�߇�u���O��+^�#.~b���	�80�����k����Q�w!���ʵ��PC�{(<r�e�5i����w��澋��f����#B�WA�����/��4�ek�&E�rzJv}�8n2��>��m���ڣ�.e�%^����BQ:�Ig5j�Hm�Y.קdz��ރ���%F��l�E|���3x/:?���?�A��L<�k1�)�_����C�!%�Ex;�L]��>{�z��V��k<L�~L��2$6JdӲ�	F�^�\|BrJ�p��M��[]`˴G�bA���U�"�M�Buq�N)�SO!� ���!�)�x�a5�x�̎_C�#�q���?�� �P{�YV�6o����!�s�t��RH��0\i8�;��u+ȕ�=(K�zyGM���9Rf�$=��I@�rm�ZԺTLJu�!~LWɶ�ӄ:F���!ɋ��C<����)P�������MȌ�	�U���A�@�N�����NlaBl�9�*7�k�Ϛ����.�k�^��׀��>D�x�I2_d7��lr�#�(M��m-���թ���ܓ}�z8�Q�@7bl4�5Fu�kQU�];ݟ=��0�H��b{��N"g���!{|���'*{Q�T�A<��J!Df Ou1�p�����;.��`m4߯�sy����{�B�PZ�Kl��d�]R�g�F\�T��y��I������@	�ѯ�����%���
g��;�g�:-G*�͸�t��&���� ����~l[~"���XN�pDHW6�M��x��?S(R�*��
��|��<��G��I���(��^��1��R���X�x@��W0�l~����+���w ��d?vɕ�j�R_8R���"���ú�������D,�0�$��	�,a�0D��T�nH�֖Ѹ�LQ��"�we�����)�Q	�lql�����BIr*zك��5�`3�( ���-"�z�/�1���L�7^d��O��&��B��j���p���FV��Ld� qP�k+��@Ԉ�Hę�������.�`�`&'�|�] HL/��h�cL
�ꈊ�+�AX��A=�'Z�`
N�9�����$��Iz0Vg(+V5�;ޏ]_�#��k���X�H X��8�ߑ�����Ü5n��i榞�ѐ��Iju��_��=X�EĀ�O��S+S�;��IȹX�H0�����~�J����.+��t�Px-���-�����n�z�ɔ��TJ�sl(�\�8�?/�\��ᶝ A!�Ny�� �q�Q�K�G�Y�XNOW_�kA9Y�^��^�g"��3��ް�uw�-K��w;���*m���C�ͩ���[oԄ�A�����|�Aj9)=yN&O�^��+��it:�8y��4�lM�|��uB��>���'/b�%@2���ς�~�����K��G�����/��v�R���~�e����3�^#.\Q�"=r�c>Y�2(������L�)�RZP��ӁY 5��]�QS�:�Ƞ�9��H��;�����K����P��iXF���ݍK��	�QY?���2���h�i��&.6�K<6?ę�R]9v� �!#X`e�鄘Y�-��"m����.�_��E��L]y T��Wn����M����J!B�� �}Ϛ}���e�ʒ*�ؗc0�dg$�m�[���{�,���ߙ�<���<�{�{R�Y�W�'�e`��_3ƨ2T�#��{Y�A�8G�8�(ѥW�}S>�<	?oJ���K��g������kod���}��'/g���O�.�"@������9V[�5`��M���2 �̄�e�\��Xߑn��r�O�n�o��R}�}4��n�g&+*j�3�\m\� .Ȋ�;x�P�'�M�������F=��*P���Y�)�L((�	�� ;!�l�b�+�W 4v9����1���;M��f:=74�XNw*�{X��?uC�U��$�GrobH]C1�Gw~Gf=��h�!�G�(>�n�>}�J#&4�2�o��v��,]�8d�S�?L�r\��gCլ�_�����S��:��h׋��	��e����v��S@V��C�}�������o-�U�W%�'T����v�юO�UĬ��_��E)��ۻG,^���g�w��6�y�	PL���6le_��R������"�w�)s�'i��kb��a��﬉��`���f�c��0������
�
qHD��Gt�M��.�k����3w�{�3�:��K1��.�2�ك�:B��z`�m�rS�(@:�0+����W�lI����n� ��>��u�S����5�t�k˟g��eÚo�]�,��ה7,�o�����zA:�(.<h�3��墣�E�_�>�������g��]�ډ[ty��_#S����my.�& i=` kh�\ս���BnۦO ]8	�IF<qg��还<-��VS8]c	����?�^����	0�� q2 $ׄ����Nx�ó~�Sp�O�9q�����h�_<gW�|�Bp{��%tbn�N�ȡ[�]�@Г����&'�u��D����������f�Dz;���O��<d6���~��1��T`��ob%���h�S�f�*��Y��̀@l��qn}	�?����?�t��'���1�n a�7����+o�N<�M��1苒!`���V-��o��՛o�T��캫8b!�n��6=���?V��0�*P	\c j��*���g�\5X�V|l0S��$��]:߹`E�������E}I�R�(4(������[��-c�y���"(�X҅�����E^î(�ѻK��+��_��������Lx��~�rk��N�0�䭁��;��6�_�/�< ^Ȗ��:|yK���Y��`Axp��&�?ua��4�pJQ�����	��@�p˺z-s�?-/���egt]�}�+��wf��Y�Mp!vg�/�jj�J6�15	1zg�����-�ٽ�<	b�?i�4�5^���U����`<�fy|��mP��U���6�0�	n׫Q�x��a�����1A����A
�H���B<Th'e�ډ;�t�?��GН/	ӿA;_sh����݇�;?}�[4��{'��k�1:z��
�"e�7�m���@D3�T���{�H�`
k
^՝� �'y�4<rwpu~Յ�`2{ uee���hg��|t�\�t����2�C�Ԑt�b
��^�D	�!y�.��p�{
��.g�R�cU�-������ۑ�y�#?�KM�Z2�駘��Z@J)V�\��=�{0(�ï�*�������Q���z�t���|�.?��ea]��p(�	�3[��:�Hh���	�[��(	�~�^�ⅴ��������Lg�H�6�a��kW��Ar5�-Y��L��y���FPp���f�nhɱ����T�Z��o��~^-!��Z�S��`UP�ϭ9�֡���K�&�������1���@xѮm1�n?�s����h;��� �J.�ܖ�O�l �z�5Y�8�u������0�?��Z�etN���i$�\�	�Nm����6�8x׉�BM�w�JѰ1`0�KW�:H4�Nlm7W~E{70�}O����0��	!in-�O��;�)	o��J�f�LR}z	/����4ޣ����(Eð6`'��E�0�S�㒥�]k��.��<�+_�$2�Mg����A��:K�+�x�@��G���q��-�'���%z:�t�(�>@ eiZ��nd���|j�8��z_g�/�i+Cr����4�(���<�&�3� �p!��kp>t]�P��#Q�
@Iç&�,k��p�T=�cP�=H*Y�$���P!�����U$s~�5e1e�Q&���Y���͙4����럿<��x���s5��O����G}9��{�����''�+����>����W��Y;'�&�8?��B��mɈ1��|7�P�p�_"C�6;���_{{��w����:N+Z���>L�?>�q�j�e=���a�z̴p�|�|�~��1>�g���>�xtr��	tu�S��?����:�P�k�|��l�c9�kS��I�;��dA-�n�>=i�=od��z�,�͖�1�j���\��8U�s��>��p��^�Ì!��:��|&t�LV�!\���ӴP�8��q�L��7,l4{���S��p9W4=k�WR7F����: t���Um�8y�뾧���0-߫u�9�jb�㏤®�M�A!)�"�i}���ۏ��x�&�i�38G�q㫨:�
�|�Ęf��q���О�*��AT��I�!��Όxbg٧~�l\ �|6{�@>!c{jpJ�U`=o7ae�'~��PPdx��@���� ��oo���L�
�D;����D5gٱ3��A�ί'�z�J} �FL{�9�)#cB�-i���E��AY��O��W�����������gB�s�mm88���a.�f̺��1<\_L����5���y�Q�������1�tl�9�q��� �%�:}f:��3(F�*.��i����;�Omr��M���LI-�� l�	���v_�C�N�u��B��0l�����O-��U��Ni�֛I�嚴#��c���>f�u��E^�>?��J��ar��o��"�QS'��Qm,�~��?c��D�~SU�C�eO��\1��Iiȟ��䞏�M=rVrȮ #q���������ͦ�M^���M�F���_gb��Ͼ��Tj�p��+��_�{@l���Gڥn��e;<�W͘O�����4��z"?�C��P�cU����ZgĜ/�����[�^�V�˶<[�X�<7T����Q���:�|��d��i	��Z�î�#��}f��=��9n��������{Fz�9Jg�����	�U�h���W��N��d�T_�x��jd&�̨-W����Ji�3i�%g��9�1�����6e<����t[I���,σ�n�釅@tY�co�˗���)�YL����yǢ�5i��Bx��@|+����'+ +#�̕�Yd7Z�*�Hg��L�د3+Ε��AH-�*��C9C_�t�cj�UB��'����1�=�% %�� �^��퐳\�_����M�}����T�]���+�"V��ES�$'���;*fB8���	�7|��:~M-V�������VN��O�!#+l��2�f�������:�a���,,r&{~a��b��gw��ȉ՞�z���z���@������%O�N� ��}�/�	D�! �M�d�/��~eǙ�Z�q�i�3�?�Ƕ�ݼ����V��U����@b��(�W�w/�/{�o"t���=�IQ���*8��+�
�-���#5$���oVlu3����U�����h��ح~�������gߊ�iٗq��ᩯ�5��jo|��4Y�}�e���L�t���M`�/�UѼ��N�<	f	��!�1 Fq�I���IK����:VXY��~u�v+?�&����V�.�נ��l
F=��i�5"M��/b� \)�+����S{�n�O���k�~�bZ&Y�����x]�o���۫?����Tbh��`�kZ*�@���4б���"��}�X��U��Y(���a�K�vU��8����X~��ɡ�:|�2�AV:�.�)�KJ�����+��QǘX��j��ט��B0�v�%ݔX����zI�����1�>I�*v��N:�T�S�>��}Fc��~�G�d��Q�U�,�m�O�,\ɯ}A>�My�r	4X��M�|��}�.~������䳎�UA\�/�>ԑ��w�v\��3$�֥%�3�Fa�%��tII�2��a�b��6���,�=?㱬r�-"22�#%�����m�.4�_�2���|e"����\_@/��������C�d��C���ȴ$�۵��{�8���Z��dx>����9����ۼ�;��2ۖb��HǬg����Mj��#���(lE�^pm_6��шL*�(40�W�ǯ�=�/�"K^����?Ȏ�Q}�i�rQ���r�Ja��pJ(E(�O�èˤ���?j��tɻ*1�3CQ�ǙV�f�Xe�7����4X�M��zm��N�;1A$��X��=�L����h$^'hB�j
 A���+%I�X��£}D/dl�,�j[tPRHB�N��u�9�l�����1����4�_����ev�o�D���P$�PXL���ZiJQL����Tr|�;���1Ӫ�e.�-�d��7�S�6�Tj�s#u`�a^Y	��o��va��<�5�~��Г�	�L�E�\�a�W�D���ݶ�M�g��P\c�,-�أX�ƚ)��`��!/\#���wC��Ċ ����eb=��<*�-cp
td�u?ɕvO�N���v�1�jgEmyE(���\��a��G�Ω_�Hˇ�v�
�X
n9�hj9�I��5Q�z�l��5���>�j��A}Q�0�j+�O��PjȆ����Ga�����#֑��s�5��$�7}C�"b&�Ol��'
�DՏC1�� �j��C�l�uGd��{����8x� ��z6	��nTc�ρ qr�k��ZJ�5X��A%�=)���}����ȩ� p�c�rn[�v�8n�j^�@���`^Y�3pxe}��ez�1����Bmi�֛q6���)�я�g���G�+j�}!���aixW 1�Vj��m��z��Ї���,)i�1��k�JdW�
;&��m�Ѯ�l_6KE���yX��x�v�����2�p�\�A潸��P�\˩��G}ɳ�Qli��m'��p�E��хGNj��f��e�j���1�fim�� �T8��O�E����˿�6П���B��q�='��������
!Q7E�4h�b��e�Qf�Sb��D	�� �J�m�hj�Ciq�����\�t�3���6��H�l�� V�c�m�DK���:�]�i>G�L��^��_Cy����v�L.�L~t�K��Ӈ�g�t�C2��!g��sdK�*j=3/�*1;L��<��=:�|��)m���4@�����"W\'h����-���{���c�y.�9��d��緋wTeM^H��Ik�m"{�����ph=Ym��ǩ~���yD���L#9Z[}�z�����y�W&CE��u�O����-�.�pð�/�N���HG��N�~�$r������%2 ��0o����C�B�|+ef���8��L�J ��7Yq���t��om^6�K}�>wO�X�jq�_(�z�X<�@"�C|5��d*�rl�E��[��ֵ����$���:C3��X�z�F��d�<Gy^'���L���
]]3Ɨ`1��GTo���2���w�e�hY�>/��^&����CGHA��1��&��9�.�e���B?mZ�cnS�����P��,ʮx�Gm�yMh���%��n�d�Q�,����/��h<q�ʹ�+nbO������1�L��e�-��|<4��a������@3�n5^w��o��PQ���f���ōt�?�s�:HKvf��y�2��M�1�$���ǝq2��qg����W��'lфTӇ���Ss�x��v9�cL>r��/S���W?��Ƕ��C�#�_=�G��;�=(&V�>={#�E¼�=Zb_�L}���UB��j��x��$����6A~�Q��K��ݩg[�dU�Si�9���w,4s�"�������D&�k�μ!�-�'����\ӾE%�.� FG*&�r?o6?��Jv��ު�3A����x��k��{4P?�ߝlm�T��.bF"��:F�L2�:�st�Q]���T)w���@S�T��u*H���//߁^�Ψ�@�b<�e1�>���F5�U��=C����p����+A5���bk���*��⯳�pn��H]۵���N"�;7��dq+Rܫ�6gM*���M�9�s�,�$�A�+�fW�_�-<�?���P��t�C�N�=�a��|�6i���׽�u�m�0>"["͔������Wvg�P=ƽC�L%�%7��G��Z�=��v��v�h�;;)�٤��0�T��C֬������᱁ý]ب�y���_�ɱ�ԯ͒�{�����[+=	���p�%�)����Q{��b{���F����c��&n6w��� AXZ9�]�ܝ^�p�}C}���.���}�$/BE��͊d�� �5ȟ7.ܩ��� Hʼ,��[��[C�-�(�P����QQ�)�G�#�UpqJų��s�����k9mI�^_�]�b�l�iz%h��]���)�BYH�[�X�ZɄ�o�Ou���/�"�"�����3��,��}'�����{`�u5��H}��"�ӽ���%��||��	.�C��	�3?��h`B>� "�5O�;4�����A�iiE��)D1|@�i�=�p�^_������̓[L-4��5�@��F�)���ZKm|3Pf�"�ƟR�q��8��!�V�*�� 9#���G}XQМ>��$j�^K��B�xh}b�g��B=���A�.�����Hi��������_�`���Fk�,��@�#w��c�m��ڴ�7}�2l�׽l�!eفY��$Z�>a��S�w B�nY!禱IY�qNw���c��HM�r��#S{�M��ų�Xj5�t�������Ƹ*��$"���B ��C�#-D��s��߉��h��0h� ��>�R�����>�Ǧ/ u�o+�%C��.�dD6�����ѕ��G��H�(�ٿ*��v�b����l�+R���W7�e�\���OC�>"���([j�|תM��+BN�յy�#�2�Nc���+S��q��0�3oS>�Wz�Ω��'�A�A�K�k��G�����6dۢ�_ H��n�W0�U��<�Ed���@�[��WJ![P����ق-=�����X���U�qd�X�Cg�؞a�}oӾ�;��ˀ7.��
v�t�v|_.�@�=b̆v_LJD:U�����mg��&�O�(��2S��UEEA��n�|���ǳ?I-ͯ/����ۘ}��ez״�ќ�����N4}�J&VH��f���jB���i%�a���4\5�����Y"[E*�V��v�Tr���36��/�����DB������P0�a?Ud	;U�%^��U���d���m�� ~��?i�&d��k��IHĩf���31t�P΀����[�Mb���ČeS�3�ڵ�~�}�4�xa��GbS���Դ��~��b\����QAվ;��Q�5Cu���9o��ۇ���C�~�5G'[����m�H�A���6�瘫!���ؿ�Z&ܸ��?-�B�ߧ���g��>9@���BJ}/3����D/�2�e����U3�f��Z��1^au�gO�i�B.:���[~
��;#�9i�Q!YN��ъ�U(�����K�r�/T�^���)��<���������V��[�����P�$^R�Z�{I@��p��jc1D�t�r�!i�8v�*�y������ït.u�;���!�� ��N�P�"vIqo=_f���qE�wZNI{�$�FP�C��[���y�l�K{=mտ�I���9J�"���G?z��}���Ї
v��2�F��\F�Л�9Ax�l �� ��Dñgg<�KwK���wv_@����n� �HL�c�]3���"���뭂�)}�bEHDo)��[�Ib$����X�uGsbg����<!rd����q�)u0��]w3�8��(�@����#�(w;��9v���Bz����X2;�8��7�6�� ��r n��T7-�˷�
��"U��Gdn,�x�ch"f��{3�>�Y��*}P�3�%���)Q'��JG�*ʢ`�/������M)�K; S,ӿ �a�[�����qo�>��x�A��K�gV��z��G
ެe9�_L>,���E�#����n��o���I�]h���ta}����Y�i�_5� %�ώI��Oj>�8G�=��6����_��C�By-D�6DoY�P��u�`��QԀ�'r��mE)��1����jn;����9|��@�b����3����M�,|�K1N�Gm~s�R�'2^�{�&�Ɋ>���&Z�0�k��t������C�g���G���QŗE�*v*!���ߟP8a�];H�<����섾^;�:$W+K�CzQ�!ȱGn�ʗ݄�vi�����}@�Ї)bh*1�h�����]#��p��1r`O"F�0K�b��ΠfHi2G|�Y�A�D��	Pg��p�����>�]-�Y�~��A����HI�t�9������}�Wq[gS	p�"/J,�k;�u/a��<.���������`1���� ՆNh����<�ne�\���D��C��
J����ں�N�/�v��AoL��LA�|]�R��ϋ�,�JK�j?�N���R�N�:���}W�h�- ye�������< ��m�$'+UYJj�e�=���ߨg��2�A7��R�����G��U ,b4:��A�+A�n� ]���W@S~Hi^�2�
�"��N�hS��2���"NAh4>�u�aS}˺�s:Z�XDN�7�$sq�w��
�Č0ƪ��;EB��"�oD[���leB�c̑�[�:�"�[��������ي8[F��ɐ�����٣mx�d���L����J�_�g�����1Ǆ������LG_-!:#}m"�+i�C��RMx�o5���=�'E�C(�.|�1�yDD6��Z0�����h!k��Mo�"��Q��Fj߷�������9�+�D��}�����e�^2dH�/�q�XW�U�횐�Q��:A�}���ŋBAp��$\���n�X����k�k�1y����"�s�"	�����	%���1�[y��@⛪�v�`�:�s*� �:J�\��s(�IF٪Э�1�#���Dg�1��x�KǄ�g��ԙ��	�I�b�	�-��2<�d�qu���J��ߧ;B�4\����،�!;���g7g�xa���%�_@[��w`^���
��Whji<�U�&#�m�5�&���Y���˼�tH�����!��w�(�뭢
.n����D(@�c�M~����z�c�>�$q��h�� ��	��a�gw�f/hy����$�B]��V����P$�����-_��)���b~��BYȬ�Q&��b�Ɲfs��R)�l�gg�^�����@����~S��=n�I�t[H���ǴP�R���-6K�#ᒋ-��S�i��v|4,~k;���M��6�Y����ce�rip�kT�����2�I���?�~���p2�}��^�Q���N�1-��s�Y늆��e@��{>��|���hN�"�E�bapH��NaL���:V�C�_x�U�^�$�'��!nw$�ЇQ7�J�a͞OJ��4���7���Dy�I�Slc�c�z�	��"�)�DԀl�]��'�����b?֤��O�*Iv�8	:}��\�&[&X�f<0�N���Y\��+��술VWip.�d�9�$��� 2��m9I_��ֲ8T"U��H�Yv��}���n��ͺ�č���$�������
��5b�_���aq)x�W�	���[�;�W[۶�a����(������t��-�
��:#��㡍�$���o�*�{��%�;'���i�V4��>&�h��������	-��e&�Xd�7?[R�V&1��!Z ��Ic5ez�f�u��	�R���j2�]lK#Я	=!\��Q���e~�����T�-\��!U�nף�}�y�qX)T�l��.X�V�4�@YI��4Ў�R+�nuqг�*�@��<V�1�a�KJP`Q�
�cyj>�k=�����~dC����.�A ٴ'���Ss5� �+C�˧r[����9�=�3힕�٘D ��κ�1���j6��ٚc�a�0��2(	1!K�g+ ��èYc�����q�"F6NBʎ�#�h�B�,!�[%/|+/)n[��ɿdAF����j���Xw��]�԰�Q��"|)*����L_��[t��p)�?o6kH��W	���1���ٖ���MS����|���B�QQ9�,R�|��j�g''����_C�m8��˿�Ėm�(튓��m����+�Ti��> ~7q�`0c��]1v��_fz�o���x��9CeT���W&�*���wc�ب�n�e�$f��2]�5���)]K�8�OX�7�r��xh@5q��&j1l����PR<�=O���_k q��B�����Ҋ/���J��q�=coC���kX�4h���0���U�CyK/�5I".vfr�p�X��V6��]��ʷt��|_h�/h[�%�	��آѢ�'�
�	����9���TP!}cU�r?g�B�RY �9�WR����!��i��������'�o��ٿ:��g�0,�,0����~���|N	�yC9{�*�ԝ��w��ƙ����l?yX\��y��H�vA�����`G��o$���a��)g�������^�pZX���+z�q�g�� ����۱ק+���u7����]ö�{�B�X>2bܑ�q>$?]e�<�<g������I�����ߊT��2�+�oj�(�}�����z\R����������K��q�=�A�I�~��*���s���ǪE��}2}����H��#��٧���/�W�r�)��6̵���}V�q�����% �����CJ{��RV��(X����b@#ʏ����F9�:�t����s��W�Ӏ����Y��HG��o��`E �Zz
��pɁqL؁H�ed���D>��򼅡�D�<Gkc��"��*~Η�k^�GI��J�VȂ��H���,����xO�}��������c m�%:6`7����Q6��BA����߃5v�C�~	8��7}i�F+��o�zI�vB�ڜo�XQ�=�;u:m���ӗ�'[�F	X�^�GL1�E���}�>>k~����M�W�2ϵ�tE���đ�Hz�i�:��ev@0HK��qiY��MP��Tx�c�I�ŀ���oǊ��n|_�ϩ�e"�".;�\(S-<m�!�$���h�DG�J�*����nY��K�N���3}͡0��=��D����)�Z��2�%eq�`��>�]0�Q��"���Sp�*��ZŘ��,F�'�ڙ�^i��b^����!,, X���] ��Y�S�;r��n���̵��B&��@jW�.���1�Y�i{��1ot#�~N�>gA��,Y|�k��ޣ�A�F�f�:i�Е���:�:�q߳ϣ�K�5�3�[:D��t��������������vC
擔L�%Z����-���N'�_�♟�Z\�S�� ?�P���	hb�i��������sdd������;���L�j(���gDT�d�%�q	-�����Ľ �1�vΥBS��T�/}{Hy]c�n��=��v#���%����6[>58#�  ڵ~B"�n��g��� �܄c�r,����
C/�pR:�L�V�j��p��V �=V�Ozɺ��C/?��Q��By�\��|ؑ��_R�rYk���b���GS�u����J�_�����_Ĥ�K=�����:ǃƶ��{[��-������Vgق���d��w �$m'�(�����P��d&�*�+ŵ.t���^I�ZUü��5�!�*�A>�U���>�ƅ��U�vLCh�G��)�הּ����9_�۝�8�_�@��u�ݚ���s�}�&�0�k�w��#E�4���_�� ����.w�K*���?��޽=S�aϽ�#�(�թe���Uآ������|~u��ؓ��F(��+0�����a�F�o��cJ^�ǳ�N te�;�g9(��� ��R�b�N.��u?�7�N���C��T���F�k|�r�X1���_�?��"�L�P��*/|,[d%������#p�s��k��D�s�rSÔ�(����7a�Q���לk��%$N,�Ś�r�Gw��!/�Y�i�>��Oճal-��h��\ާnG���#��qk���2s%��;kg��y~�R��&d�+��n�������;~D�6�\0���Gɧ`���ʴ,�����2�A�����9Z�,>��{��w� ���Uh�mK6�P�v�[�Bg�cS<���K{�j,�4/�}��0������cbJ�6q˓"����^/�i;�m�%B�[\� C�XD�a\�݉d�NUܱ2��4یM�ݵ�L���P0��jD�F���Bht���s�0'��v�bwp�qẵ��o�*��Fd���|c�H�u�uF�rvzW�5�YSp#�Z�qXM��?	0V�>Hx��;]Q���A�(��R�~�5^��I�6J"���Ä ���> u'x�Re�[I�C���Z��P��՘�*Ҕ��2�u-y�7ETR��D�����b!
�}�a:�9���@
�D���m���=yM�^�0>�lϽul���^�B�ږ��iC]��wE�Uz��Q��5�S�g�������n^���)��"b�N��cY͊�
0��k��/o�̉�9Y�L3��L�W�|}��I9�-Ő�������M>�n� �
L�y�O�d����e�Pt��S`����>��F�	��*'v`%�k���#<Y(e T��:!.]��{�v���굜��|�\{��	m.��$�1Y�e3r
򢏶�N�Z�t����0²���%G#f�v��_�*�$.ޞ�s����ZMŔ���f�l�?6�{?��p�U0����B3�#TUD��l�>����� ���s (�8.��%
YZ���4z̟�=��-it��`���ANA���J������Z�!�^G�|E>�J{�q%�F=�sX��a�3���ǯ DWT��}h2����8C�f�X�g���A`��=l��8�ȫH�����L������Z������@��ǆ)�,K�E�zU��
���r�f�WP���Mڅ�*�9����t5��#�t���X�� ;7�oӶ�j��B����#��7�ƃ�X݂���(B~CVR�����=����JnFO��?/y� �=�W����I��)hu�4�[�K�m��r�{Z�HM�$����$���e��.s�\˰��Z_@Y7@�����-�(�,�Ro���ۼ��T+��G�{d���]�xzv����8Q�A��}cX>�H��OO�Ee�6E"�67���	Nw�~�ٵYKG޶���iA�ǬU���e��\�b�?�X!5�VFl�S��_p;8�O=IK���l2\-#V��Tƥ�:�rtb�^q \�l��s�0C^�Z��J{� ?�"�$=���7��77Zo�U�I��+ϮC�M��a�k�6J�������-�,u>�"pE�	�H�۠¥h�,���v�qG��`�iU�~î�"��s�ۦ�8ϕB�5X�Z'����jϞ����J@S���"��S�������@ˌ������[ȋLg�:M��u��a��d�Kk���6`]��3����	X�Ut�_���]X�����7�4��#:��n98L(j�Ű���M��5�����Z�w�A��bh��5�!	o��yެ(m�� �1�S�8�$�1UB�(� G@�ܫ�ո0��;��,�h�dT+>J�L!���C6�ѭ>K�*r��`���b%�<I�\�/�����s�'NQ� �3z�38��=ӣ���oM�%?l��+��Kڏ=,ԗ�fls0l��g�lw��_ �v��
"�Zy��b���,��r�6q�p�n��� q#�Ǧ�xWeӱ,`����aRt���z�Ei�w�1!e(V P�t�Z;�ah��Ҽo5~FL��l�P
���Z��t�W6�$/㈶3��D���Y��`2��r��|���=J(�f��i�m�B���ew�+p-xN����4y\��+kV1��(��6l�*��+��Z��6;X�H��Kx�<G!n�B��2aW1]�v�1]q[�a�D5G��Ɉ�9��ĥ6�{��)�˺�� �����'<a������>f�i!D�L+��®��ԝt(/�Gsn� �'���7� B�3��e��2���uu�o��Ob�pki���CQ�Od�b�viN�ͺ�;�/+��;�_Z���u�H���܀��]���Q��#�f�j�[�3����8U˸�u�'S�
o�7�� xӻS�}��G��"q}�O���_<�,D��Łg�踞蘾���k�]E����*pbE>PZ &�bF�����<��FN�8M7�`u��hX�N�r���xpp�Yaǯ�=�Il{{o��cS�k�)öp��>��:�)�<�Vo4�s^A�!&n����{��AR.���b��94��/�
�w���յy@��B����^ML� ��kN3N?���0I<�L䖡��pc�+ ��k�W\m��еelE��Z^IP�XWoPRr�������#ׅ?�f���v�'����B�q�Y����7��W'���@;�w��.'G�s�j�E��4T���mi���[�d�1e[���~�j(K`W'�����?�j�@��!T��]d���gk�E��I]F���MJ:��o�`Ϧ+M�WQDg�7H��� +{v�i�8��]z��QE�b��ם�E�~x�[ �q��<�=���L�fY�7���}�t 
A�:A�-h����RM�B8�����}̔�%R���<��"Vܯ$x�1t�@ē^d`6��L�7|~W�V^���Ěݎ?Nu�� W�b�����"��
�g/����W����_?��Z���<��+���xqR-��v�����*aZ<N ��|VM+�w�� �Z;�Xc�%>����d�yu�k�|��/������3ٛ����=�g�GD����KB'l��y������d��^p!v��9��c���y��Y�
�&�=�RaGr�"$=׃S:ғ����>
L_�)�U1�W�m�<n����1'��%����$�������c�M�J�G�L�IOF]S�s�Վ�ή�C_����Z��NH�	� ,Y}�~.�w>
�haς-U�_ۣ�E׼a��3��P��D]dz������	<��W-�}O���ٺ�ū�����v;���.��M�j�G��z��p���vKH�����̈́6!H��rt��g����>e��!�{n=�jj	����Y�z�ќ_�Ni���l��I�w>6���f�޶�a	Y��{@��ݖ���oK���w������h�<~-ZZ'~��Ǐ#�1�r\˥7E%�]�r0�۹M���Y����r� N�z_Z���՘�*�+��!��M�u�.�fԿ��G�U\d�p�P�r'��������O���9�Z{�p8�u7��x���0���5�ϰ�B�ݿ���wuH)�6�a������٢G�mԨ.�kB���J,e`	�5�,�;z#0^�G%�YX��)��]�����vAX�Y��e�0��F�V22c�Pq�:Kg��+2�����#���G�O��'���?F�8�G*)Pn����%�qv>�-�lz�ױ�u��9v�h���tٍ��C߉�r�[�������v�\��35HB;
����>�ȹ {�kŁ�7d�>d��T	��T��$]ϓ۩�;/��p��WæWS�zm�"�$S>Q%B���_Ѵ�9��C"%Z� w`�ԡ�o�ߗ�&E�岅��	��2��JZ���*_�����;^���"�.�Vr�ʛ��"���>�	��8������P�@o���O�#:��!�7,t�ΣL�Đ*(�Q&*�����j�1?�/����t��<�`����`�!9]���E���y�G��oDy��xJ>�v{%�c���`3RZ�����c#{Q+��]�~��%ܒ�v��ݏ��n�T�B�^���p3�
K��2�v��V��d�)&���ծpA==�G?�
�sC��i��T��F>Z��NΆاr�=W[3���m��:a9vň�E�i�0�Mc��u[����ʽP�*�XM:�Pk�-���_�8E"w\��B�F*�n���b�!w�l�=�����w*b�ekD�B��|[��ey�E|M)8��7�G*�BDʨ��ĭ<���?�
F���p�*��k+�)St�U��t:|(�6��m)�O��E��Q+��o�H���\�����a]vkv.���W��n�危S��>�B�����F�%5�*��j�v�˳G�(��$E��P��0+{�Z��H�~5dϖ,��V@Tv?�v9}��UK�~�X�F�H�0��V���2Yb��*�#��@�:�_�Rx��^��7t������j��0|[��:���BC�evxʦ�D�r��� 6���kR��k"�ބ�M�������E�ŧk2��8Ŭ���6���\N.e6�D���[������u�\|E+�>��*o�V�k#s�8��WQ;�i�}h���j��\����s�UX*MT�ԿVm�rσ��1h���|�R�lz�G�F0��R]��ȴ��U#� sM�l����ل�2�~Z1�w0��T_��2g���8���(Ε;* *��_�.�jhR���D	��Ƌ��SX4����!�݈�=�c��#���y��S��k�}[�`O�>����!�=��W`N?��h��H/��V�Q�����Z"�ҥA �%/�|����A�x=�Y���^Z�zB��ZQE���d�#n��L~S����*T1t�ȼ��^��,��r,>?3q�ݧ4@����1���C�Ae��q�^����z>���~֛@�A�t��?�
DM�_ԙ�G�\�P��u�dg��m���óS��"��+d@��j?5�������˝������I��=�5a��2n��E��L�I��]u�W1�&m�ބQ���ա��R�Ϩ0���{�Ǭ$>(!��Я�Ɂt�O�<���.ZN�ui�5�::4LƆ���M/6i�`��s�u>��,ۯ����M:�N��W�`v!�К�8���Kat�ϣ� ,Z�~Ls�P��Dj��T�$��U��*}�As.���dI��hP�0�nx̝�V��$�bi��i�'�,�H@\�2��BhC��9�QjW[nqA�g������Ꝇ����m���Ra���y�":Ʉ�����3�a�y�ʽ�X/Q�n��b�sxD�P#�H4p�_���?��Ը�W���9����˭�)�T{�Q��N�4.x|�� �����Z�m14�炦�3 �J]�����(CŰ�=��]�V��;
�'΍���L��aE��(�ě��5?������j]fTk]�׸�M���N�����霿�X~�H�]�b��P�Y���$SP|�r4�2�[V�Q��[��܃|�7���P-������3��V�%�I�[0r�"-py�0�Gh�?Sm�(Ug ��1����þ���P�8S|I"��N��tS��:�j��{ R�~+K��]�n�ވ������7��Y���8O��"ﱘ��#u�<��Dܳ[�.���mmQ�;���\r�@B!��8�rV��[�|��|"�����5e؂s�S�m��	��܅j'�u��� 0�mo2.�l?���Q0��ћ/��rў��|�f�ݘgg)����~r�'h���kv�/��>����Rn^w'lL�:�G�ێ�g
��0)p�ͣǒ��ۼ:a!ʵw��M�<���$`��̻���ǜ�DfQ��Z@b4���焪�]y/���6�~᷅��0����Y����.�������aM�q�0���� AB���Fi%�%���"�5L@EEZ@@@B�ѣk�tw�Rb�6z4�k����7�q�Rw���'��y�, �A�'�d� 0��Euef3�ۏT��5x+�2_S�7�X�}77Wv�+���ϣ��8� ;TZ�r[�!�D�ʠ= �Q�����߂p'�޲BZ.�bCG�30ۖӖ9�ؚEb�j��F��	Z'ʅEG�8V{r7�O�W��We�Ǎ�O屚����p'Un�7Xi�u���Q(���
�n��&�}����b���h�?Ka�N��a��ɲ�5U~'Z��׻����M%��`L����見�pt#����ʏ����;�:�׈�Z��'��fO���1֨d������,�/��E��䷟cq���9�8�N���,��,�����7l���:�.P�f�S��ɗ��Hl=����G\	�x��a[�����?*#E]G��.�l���4�� �C��W����Z��y��G��.��.I�olZ�H����p�N#�c4QX���7(������P��667Q);4�I2�h���f(Z��5N����OI�f[y�����/m/]Z�"d7��4��$�7�E�<W�!o����G&�Y��]Eڣ�H���7�����2��+�V|�|N{(c]I'[GL��)���4l7��F}Ĳ|s���ϟɸ���7|�o��m�njT�ʋ��<$�xs�� K�2�{YIe�Η��r\PJ��G�t0�0i���\��%kv�9����b%��c b9�،ryA'{����͚-��[�N����R��]'�@f�vK��b��Ǥ�2о����ą	^�e	+����nE�v��$�6���V�����E����ƼT�У.��4�u���:[1�������C�㐛[^|�!H�)'G�E$�D.�����Yo������'�hRq(�.����鱣�q���\[6 H5/��Z{���6���@���PP�ˮ�~��Nt^̈���/���=�n��Y��L����ו�*yͥ�;�p�y��6��}��45�²�O�����]w�}����x6�Fk�����0+�L��i���h�}L?��4�i���V]ǀ|I���� Y����&&���noQ�)��x.]��ktj\K�:�g3�%�v( �~[��#y��	!�z/i�u-(7;��d8��8������;�׮_�c@9t��k��au~  ��_�~�&�/���F+�C�c _3��JqG��x���߻ͼ2���H/|y�	qy��zM�ʬ�	Er
k�e��N�'�iZu��S҄R�ٵI;\m����\�-����}(@%dc�R%��u�B����2Gj���/��O��R�2=����7�Q<�l��d>��n��I��[�� O�u�P]_bh34�N�s�'����w�Ls��a�Z�M.+�*�qV
1a��:�܉4��
@��jpWN����e������{Y.�I������ķ��@ꉓ���\j�N�ЩsKg�$[b�L*��P�����Q*�
ͩ�+�G�,�V�[WkU�F����z �Y�I��1E_$���X�9^�S��gRW� �%�H%dw�NG�,���O
��/g�2���y���h�P8�(��7�me���<����P�/ܽ�_�o54ЧW3n��������)R�߈!�CFA���X7N�5~
>2���/]A�N�Gw�m\����}ƙ�Hż���M9�mE��<Ù���%�n���]�z
�y�?d��u)N����p&�H/������a���;�o@��m�^0=���\`G
 �|hN�o� \3YQ,6��8�s�c$脸���@ƥ01I��^�0hԜ�X( í{�y�t�g��d_q��e����M�:�- �K�`�s��-N �d���Yp���]�����j��%>z�۔�@�_�&y��}��o��k֌���(���L&Q:���b��0�A���r���
��o�o��`s+�B�2�ʬH4���}�Υ����z!�e�����[�[��"���1����o蚵[I�N�R۝�n��e�R�Ӷ�X�tY1�ת�nf.҅%��v?����$^��L �� &@�̐�����*o��<�cJ�$�C��<�sA��`ho��)�ad��(B����-Z�13�> dv�_<Ox�OpA�
��3��]�a-�&��1%nya���\v���m��r�kYe�M��0�y\�ύ��=> ^��	hMO���z|��&�oIsV���>� 4$�FJR4��x̴8an�×�s6��AfO��Aqg������9:��z�T�$P�u��t9Ώ��i���Օ������a<]��ZW���K�L_s>����n,i��M��ҁ�[g_EB�_~&0�ˬqZצּjM�W����Fꦻo��~�:��ښ̳GF�C-{��A��?����X��xI
����2�K��ޱ/#�8+��B3�NB�4d�{��HU�C����z��	!��v�E@�(_{7q}��}nӷV��^��7�|�Lז-��4AML��3b��f�1V���s��Լ��d���,+�S1�I�p^_����+�c6X����GI���W ��c�71Z��q�|�0h�G�lÛBY����4^.e]����z��,�='��5Kb֢E���+~�Q�b�)�|Ҕ! 
�*6#��<=��X��i��9H��d��T�Q�����9����*��N�e��U`~��L�+������*t�x5l����]R�l��@Z�+�M����#%GW x��Բ������� ֽ$��"]���]0nkd����qYDcn�Ƃ��q��\ ����)�YUs���	��ly��^w�3Δ4�j�T�&�s'�L�f<5����,Ǿl���i�Ahn�[�ڭ)����.L�H[��5�/tfveo��Z��rqq�C���/2����3�:lv��!ɘ?��:C�
�t��d#76��'TCUR�N��Q��ܺ���餙R�6�֔17��ַ���P�%�M���inO���{�ي���'���	��3#����1V������0����2	��������O��˼(|�犙]F�m�ǖ�+���9�B��/�e��Y�.夏Q�vɯ����<�VwҒs�!�z� �]�ԯo�x�h-�[^a-q�4˚�on�ѧ����P�t�5��Z��&��g�Vb�G�FO̙��nY�v�Z�.�_�������q[]�%ճ���O-:� 43M�b�'����/4�%	��cc:��WF�i*H�п
�Rn�����?UX�I��S$%&��ݚ������<��;Ah�"� ْ��9�ka��ܠvw�)3{p�~�B�1�t���lI(`<���_m�Xr&2$:��-�A�zG�k֓0�<�Қ7G8N�%��lW`�ޙX(��H@�6�kP�j8��wRdtZ�ʺ�i��������%!R��idM��g�r{fۊ%1P�[�����V��c�VZݭ�e�����r0Г��y�hٽ����?t9<>��������GV��A8&0�[����`�j����볇<"�p{I�J ���g3�u&��������G�L��	��JV瀄�$zT�5��ޤ�E;�����K@�ON��`���AzP��q�c���}�W|���_|Z�1 �]���S�LFV�vT.J��o+����V�c�������-J}� ��2���-$?&�I� ܬ\���>�B�}�I�N���۽po�y�h��-��V��Qn��꜅R�#�+�ݠ���En��#b��K�����Zw�f��}cWrK�/D7k�(���[ķ���c���#��$��8:�N�X�LB��b�D`r�=�_�4=���̍�����w�\��].�100�E�i��J󅹢^Ӣ�c����=�,��m%��Vp(��xR��֒���OzY̋b�O�K+��|����t'4���*n� ��=n!���0�����(.Sq�S/���ˇ|�PXZ�d�k&��[�oہ-�5�~%��sY��� ��đ1�Wn9�F/t�j��F�����R�i���s-���0,��2�V��6�-Fiq��_����m5sE\g�D�eךq[�r��`MG��X�}#P����*��ԅ�Sr���*W�i��Cӳ� z�_`�}�PC�I�h��`.tz+�|��|��3?�F\/�(���}��������
jfQ	(%e�*�m��?(��@�$��Om�g�7j��u
��Gz.=�ta|2.P��v�Ί��::����"� �01�]g���R<����f�i�}+� ��W�	?3ӜXny�	�n�v�<��R$�"[<���x�W߲)�7����ʼN��7'L��H�]OY��;�Q�$hm�~�o��R�n/ǩb���]KD����%�~���ߐ��^��~��j%��Y���ڙ�ė^�Jѩ��A��Z�L#�$��w�C�;�$��8���x�h�-C�	Cͻ�����4> ����ٿ�����Y��म��e�󻓔I��i�8z�~��f_tLzϗb a�v��+���]��1+�s��6V���V@Q�-��<�ԣl]�|P��������B&[��%M+X:;;��O�<��E�z�,Eʿ�O<,��w�\(Π�[=�� �[�m�?����Y���k����n�G�}( aK�?���,2�Md�/
�o��&6,��X����(l�L�SYэ��h#�S��&}%B.漐�ч� ��O�[��ԯ2Q���OS��,���J�A�&�'+p�BbR(�>� ����|��$�\�m��x
�Q�,;ܷ�������j��c0d�l &�eg����l�s�^�l�d!��(�����5��U;2�H�FT��F�!O���-�WʝA#G�d��H�����B�WY����4�.��`=�d�="�y�*����$~<�Vd:ώLV�!��xb,��Mn������1'L��Q=L�9�דϱڑ�n*ja�a&=�_+4�.P$L��1%�	���5 
+��Y�l?2&�J]����ղ�;H��2wR�l�����X���� �������U� ��]�K�b��j�R� �O�fP�BHsJ��
˫p}*��C?d%���ߚ41��v
��w��	��B0� ����[5�V�)T-��
�w��K�eOG��$7�JT�ʚ�
J�YQ��ٹ�>���ϧ��]��q���}]�0�S�&ѽW���Ʀ�ye��DJ*7�a��߹݉�	��G����(�0�դ˖+/�@s*:���o)�X�'���bo�=�e]z֜�h�]����ų�R�Ν [y�F�pO�í;������;*6&r)X]6\�~��"&��ɭ[�f���ZsK1@��\$�٣%��t.��S��-�P5��*D������|�q5��z���<Lq���ۿ1Z2����?{��??��?��?m�3���?��&�O���w09go���vU����Z�4@1��^8���C�kd�M�hosJzdԴ�h��פ�v��"���8u#~I�'���7ˣ���Q�وl8w\�Q�	Wb�kk�q*�*�IqR�Å�O�8�i��w
��"�z ���t�E���zᵄ�BiW�|T�l\*S�����^|zv`�)�I:D��lF�Ccc��FY�D	���N���7~�a�¼��P�|
#`H��y/I���g�&��/�1O؇%��{��&󌢓dqO��wjaX�2.+���q�u c>��}��MGHOO���B^���	�F]�6��?P~���ˏ�}������������ū�/���*̈j��N�;��S5��Wi�U�h�I����%��)o$�X�'����x�^�Nj����6�Nw�;���wڼ�o�!�e�R	R�/�	zY�P��3<�Mi��5?v����J@o�\����&���n���K]��yi�w�s��Gȩ�����xj�n:	����Q�������!�ĽB���e�WuL��C����ֈ�M���Z�ư�H4�@�b�hg���g8ū��~7�V��^-#������Y#��J����q�$�:5�'z��nyL�yV�s���.�����<!�MW�I�q�g}%^�l_�65?!m)&t��=�5�^�ЉH���|9z8}��!Y��i||����㥕�+>����
�|��Ǭ��Fg���$ŉ��M��d�Kj��(���d�	�_��߇�+��xi]�5��������'h����mi/����;+E:����;d6}�s�XB���X���ǅm'�2�ʘ��5"��>�2��5�]S]k��V
�ʖ����G��<n�?{�z}6H��m����^!�v:�r^z��6kz��o{f����������Z��uf}�{�n�eXn&wSg�ɬ�-�����ߛ�U�m�Bb� �q��VW���0���)���_B����Q�l��_W6��B���^�\�@ؘ)�-���TM����]5a��g���¢�?�������4F�g4����;�3�s�2�F��0�M29���p��g���d#	L0
�ZJ�z�v�(�m-�](I�(]d��I?�y�ڨ�s+������r}J/��`
_�Fڳ���Ò�C��9'OFݪ:_O.�u�w����k��Ĉ�wk�B�n��j]�`܍�移����(������JF�\i���1Lպ/j'�G�H� �R�jXu�G�pPP��x�&U3Y�/��~�Y3	�Ǩ�.��5@���}n�RQR=�X5"���M���afzz�*G�^<�me��w�dWݎސ�C|�;�����F'Ů{�0��w�O����?l+��ZcËC�mO��Ƕi>���A�mY!��^c%Y���C����;�S��پen�\	��H�閑�;Y_J2�X���E��TG��#\������V[D���a-�&�m5g���u�O����
ɓ�x�y��N��Y�Ě%��n�|��ɕ(��� ?���*&Щ�>c��N}���~%>~�A�vy�i�	�L5�������'����YbM���\��XEe0�@�銕�I�Y���"�$<ݵ"F0 ��_����R�
�tEFDn>��f�M�L=M=�_�'į�@u���"���vv;+�&�`��Q���/�h�>!�7���Ք��ƣ*�����s�Qq<��%�U���1];2?����s=3ٻr�qn�(;���n��DH���m��"�:L=�0������w61"�-�����Jt����������8��d;<����~��i�Kn9Ϟ�[[~�ͻ��@Y�:it���D����'�:N6kw���
� P-
����w���io<�� DD��s�J�n���,��R�A?">n�����w.��9��?�S�/H��Y;Eo��ڌ���H �	���'��%��*++M���`=��`o���u��TF㶐0���Vꑗ���9)U�C�^ 㝰�ۢ35�W����9Hk�d�AO�B/��s�n=m�/j��mc��/�M�2u�\]���N��R=�Y�h?}��&v<�����x�N�.���hJ5f�/o�Z=� ���BM����z!J51i;!ȎeQ+���zi�CާGĒ�(F2���4D`�t˱!���З���|�3SU4B�t���w��K� d�nVڣ/�.{i��5	��K:���H�u4�x�n􎽛����O<��Y����=|�Ϧ|+���
��O��b�gC���-�9@��U7I�R�Y(� �^����!��䯺P�e�y\S�%�x�G<��8�zlydtnEd�&�4��T53 k�e5'>䓥�>�c����ǈ��e��V������m������^P�M���_f�a��1�ⰶ_�Ny]��L6r���ن<G;?|ć� n�`nЍ�~�頋�I.�+C���l��R�pPf�������g��<5'I2'
�c�)an�Ӝ����pW�b��~YV�<��2O��z&?��S�єQC-�CL�N�W[LXf`
����߈��>��&�N�ƒ�"�*�HD��%4���'-��o"��yOޢ���@��2qj����Ù�Bi�h�Zb6Y�sB�	@�����U���,���dW�R6Ά��P��7T��;�,=�I'�ꏭgl'3��ݺ�����WHYs��[��a��@��Eܼ4��{c�	�+�M��cN'��y�&u�%-�����Y�{ߊ�Y�{k����8^�o�=�A6�CT�d���P�7:s���
!��	���1ʐxu���X���9��wyו��*�6~������꟝�.s��G�\1:0� ��E�	��Ց$�	�0�2�����ɔX���6x�q����	UF��%�8������W�Wq.-W�Y����>�g�P���] w��>,��.�v�RU9�_��{��� �x`P���Bwc���P!_^R���]��k!�nrSD��*�=���.O>��߉�Ъ�6�L���۴BJ�-�%�m� �Z�T�5R���P��݈NU
P�T䇄>�	ںR@H"zq�^�č� \�>����^e�1+c��XK��#}� iXR��G3�V
MO�f��z�T'u��Ub�U��ah����bdp�D�b��@��'��R����C�O�5s���۾��|�c��}��j��6(�q)BT��+�+ �:�^V}S���7��$�G��ɞ�7�n��W�z�7j_��@(�6K{w�|�M��B�u��Tc+�d��v����r�<U�$�Di�׾��
����[��z�\��7i#3k�2|u�7� �@:��[wI�D�N�Ƿ(��ijNq�v�s�vh������W-����}�+׋ee�T���8�=y:�wFgFw�yK#�-�F����ǋO|�~��V�[,Õ!\�U�;/֙�@eWg� �}u���|���T0A]�����I�3��SE�n����b ���@�N/��Rq���A����^��j��8��H�1j���ݕd�fę�!^�H�%������a!,�#4ޏ`=��v���IW���[��|��4M�%�+S�թ	���7���>�H��z�'�7T�z�����-�(}F�N=��1��r�����-O��t<���v��p�LH0&�'��rמ����Z3�)�Qٻ���x��ʟ��q�d�K�>�i�5kO<�ȯ6u���{|�a��R�Nl��n�S+��@�N���� ��� ���Pҝ���ϐsX^yJEJw���.<�V3�:<a-C���U�Yȹ�S��י��vׯF�����<�N���W|�+��^P�J�����8{���r������ZAI-3��#<C��`r�tsep��O�p����)�BvFi�# q�H���i��h8YŠ��@?,ئ����_h4���u18h���d��r�)(e��8lU�9Z�H�}�WOl@=��|��������z!"ǳ�2t���P�T�k�v�B~��Y�ϗ����������(z��g�<�K�Od3��%�E��d��*_˜(���J��&Օ�OL����+���}�Le&��^��M��a� u Y7�����ȉ%U��W� R$�����-8�0���~d1ډ�X���.O�SQM{���}�CeH�ih�\���+����L;���g/�į�D��ao_�f�aK���������;m	<W"L���Vl��eK���[%iA�^��c#�4��B5f�L�r�� ���Xa�
���>��z��6_�r��hT%?�w.(��+�����[,�b~�Qf/�S��2{�l���XP������s�lQ9��ʿ���b���Uk�<>A͐hߕAٺ�3���X�V15OK��v�e�|7l��!���]Q��e��q�#��h/I�(
�ʳ��v8h7�&뾵��M��m��ҩ[O��%>�}c6)\���ڇ�o(�� J��ԇ�[��i��;P0���������fa�t����������z>�H*xĳ�
v�}����t�U1�ʛ(r���ؙg��2��<�4���w��C ��4������ظ?h�v��{6����q�t� �v�>��=o������pB��V�L�(Q��0���-m
�!T����<��K�M�3�s*_����ٽYI��+�h�-��>e"���!�
H�+$>$�G�*��$�2�3mJD�	P*z�D+��~wSs(2Ll\�Ob��o%����T��^�[N����):�#t&rC�k�y8��l�!i�,X���jl�p�:���/⥬W�֕&�]92�WH���С�������ʯ��1��fz��Gt�a���d���td<w'SN�-e��쫓��+c���0�?�́�?u�B���6Iv~�)<�b(.\���7}G��J$x�Q�4���͌+�v|��A����l���<1͸}�T�2��F�ke
 � �"���6��W�r�V�����~,�vZA���T���㇃?��գ%y��+V^>�-����H���Iq��a6���i׈8���rDs.Q f"Av�~�9�b��Y��R���� �D�d�i����^6�ꇜ_�Ĵ(��V�V]!���ʀ\�M�n
�<,��w#aBs��"�Sd�V���۫��<��!j��D���Uuԭ�k�:ϖ�F����]�Qv�/ʎ��Y��е_����'�d���p�ԕ���� -���}��RR1�r��z	���WH�!nᬺV��E$��sd��t2�����	$ͧ�'�����O���y��N���q�YߍY�&r���*�	��;�Hx�����XH�1�h��=��74��D=\����ưNȄ0K�Uu�$%�g��_)�T�fci8�E*�m��:��c,�^�PhLa���l��W9?�?�����2�8.?������ WNX�:E�W#2�Iyf��-`���8�Q���(��"'d;�.��ʍ�	�R'�P-Dq��7���6�ֲg|�t�����:.k�������z����"ɉ��S�u�5���^Z�Ffĩ���^�./��ҷ��M��H.�h|��0v/����F�j�.�����E���G�#����M"��J���B���qj��r�[�谄������'�5F�]�����>d���wo��6��u��z�M�@K��9�s�f����\D̘hqg*x�ü��Nd��P�n&��`�<�
��+Xq:�zY��U�؄GX�ˡߑ�+߈h���,J���f�1'F�Gx�H�Y��r���3������_�qs�t��o���RǠ�����G����Xm7�)���ߡA9M�h	,c���	4~�8���2��y��� `PV#���ZE �E����_�M#Mhq�1݈�����i~��$�,�!�j�����9_� ������y_�h�FG]�~Y�3�0J�=�7�q �'Y���W$������8�q%�0=�fPV�P����&��>��̚�iɛ|�W 'f�%/��V��0�g� �C��u1]P��ЗC���&�|ǹd�	w��Ɍ��xc'ٷ�>�0|z0*;sXu�������GXPX�8�e�i�]>9Rm�>(3!���{(UB�VJVMh��|��Ç
���7�����ml'��F���Ѷ�7�mT�"ؙ��p��O=�"�-�H���&��ec#��������?خ6�^F��6�9��4b&-	��>�$M�<����=rCf�P�FW�������p�c�����K�|	�}C?�"����y��PR�u"����?C�?C0
҉�d����un����{�-	�x�����o������%���9�q�p�9�i��'k��҂�s ]��H��% �چ�嗨��i*:�[��O��z��H}��a&�L%]iIW�*i`���]��Po��W)r�R�����d�a�}iO1��])E�����ϴf:�H�ry�iY�PԼ�gm���T�H-�z}�)�LW�Bv���4E��	@��"�*��_�.�����Y�aL���#��.f��9 �􎶰�T5q���! ���̵�U��Ab��: a�N={8G�Ӳ���*����e#��E���{}P~2x�}d/�4�-�,g;ԨR��]z��H�^�O�[C9s��N�}u��J�}Cƨ��UqiO%j� :f���0ᨤ�I�f��.)��%	e+m�i�Co�R~�涍s�8�S���dj�v�����Θ����W�N������D&�2v�Y�8�;�2{&63
�I�D���2��儐�,>�_G��9�z�k_F>�Q�.jk6T�,?��>c(���L�8
�E�b��ρe��/��;L�6w�15� �l����d��h��Glh/%:���;�k]Pk�eq�\|�'f�֦��iS0�����Ę�F� F�BT{����C����k�����і:��o�~.��\����0(���)<<:�UBڼ���C8�#v|u��h&6ˁ)�S�śo2���6����� Z}�r��mc��__	���G�_dN���cX�+'kj�B�ڹ�qҐ��C�p*�W���wM�*z?gWV� c�mm�Z�5:
8�`9�(�:B^Nc��]�C�Z��/e,S{�S�$f��oq��t'��Y@OǨgY֦�;�N﷟1�-3�+`<?5ew5���f{Y`�u]?}�*D٤7j2{����4�p_ٟ�^�T3������
�����b6뙏Y��LJ��E����?�*�ݰI�.��>|gӹ���3,b���A��"�W��?�l��nuў?�9�i���?i=��8kM黤`%�4�
� ѐ��#
���v���O㏗���L�,��lM�A�����>sIU��@!�*N)�j�6�(��Pl�I��į�u������̚:���A���K|��nj4����׾�����~��?��r�,8����Ė�%ę�R�v�����#�k�]�Z	����ᙡ5ΓP����D�ӧK��ok,|���#@oӎ 'X�Ϛ���t;�T�̗���l��$�#�+=�0�f6H��U�R�e# �������tm���q��X��v8c.�0�Q����Y�)&�*��i�XFY17ђW(�Z��{���Ͽ"f[{Qa����^4����V?�D�Tu���l�S�U��A���=#D~J�,��ĝ*���uL�'v�5{�1v8�'E �й2�<�)"b�m��ܲ;A�M6��Ӄ���u�d��b8��$A���P�u�$Rg�/z��Qy��sx���� t3�X4W��@ar.@넕-�G��o����N�+$��W��Ye;\O��`ɨ8���{�6V
�{���8��V�� E��8��4p��䥯*���CV�x���ȏ@�}pn�|�9��u?I�&]�BElCc΋Qb�Ү�u�{ŭDa�7�`@��������λ
 )���,��_
*7�����5�b-���ں�qGEO"#��h ���Zό��{��딕��.��5���kVg4x_!��$E�v.]v��
�+y��
����g����k$�e���Ws5���k���K��4x�P�ə�<�H��Gbq*zZ�9<ľՋqTW�ШBN}12Z�G|��k {�wՇK� �KC�m(V�/�7�n��ns�q.���d���x�=-��hd]�����d��h�B�zl����ߴ����8�Ei������ͭ,GR�)e�xU�N�mnOx�FoۮM�02�ڋWr�'�4��Īg��ǟ%rnZ��`�I�C��E7�9a͇���2����b/��ل+�~�Ò���"�}1���HB��U'�تP*56���d(��r��&�q'8/#u�\���g�$�D=�AD4�&57�3���s���w5o}S�90����P��*%�m�k||��&��L��|G����x묦���}��tz-ũ��oT�@�1�<0=�2u�S>�,�	4-���辚��%��,G�Q�(���t}�*&��P뗑�I���ȅ���u$���p< g��[&8�,� �O��7#�{u��)yr���\��C0>����{om����*��
���+�%߉��'�8���-+�]= z7R����ɑ?z�}h��n�k�^�u+gHeϳ�J��jL�ρR�&w����}9>���)��9'ǽ�Υ�R��>S���,/��q嶭l����ݭ���f�����
{8��?#����{�d_pŨm��S>V] ������"�J��cb���d��O���ΚAIra�a�E���犉^�.HS���7�+���*�p�;��ʦ�g�Z�j���',�T�K|ީ�|A�2�I�y��OVYV�o"y��X[�IQ���c0%��U2�����N%7M$�����j�9$��Ӳ���J�1I��\� JC*~'p&�"\:2�L=}�l����o�Wxޕc7��+�}j	�����g�W�9z�)�M�c?��.�� 7����.Cw����LO�|�����ܹ�*78�;(��=��;0�I���d�@��d�X���Aꮌ.�.j2�%ŖQOCC�Քr����� ����0�׺,����F�t��'�:�Qa�li��|H=[�v�T�9^F�Y����jH`sV�zye�c���*L�{K���zh�a��y�b�xpHg����ͨ[�{F�,��խ��S��P�X����j.�b :ޕ�φYj�� u[#\���]5�ȑ���n���<�绘��g3z��ң��
i�
�H����^��w.ֻ.��/��G����p �U����$�ϡ�W��`�+SoDdݴ�q�����᫰b�����{�,\���_�>ջ�\�4Wյ���[@Iߡ�2](y��+�kiڴ�:�Z/�?��gW��;��T�6���I�Cl^������X�x����E 7#*Y&�OZ��U[��$��·gd,m��C3�8��:n��hEѠzfh/,+>>Y��c��Gyk���z��q\`5���7]Wt�=L�]��%��@N�!����=� �J����^�Q����صci�����X�xE��m���2��TRt����hK~�S~��UMܯ�]����螺����NWO~8��u�{��o��BX�zf���%�J���6�����_�p�W��#w5.h�}���������j�XtWᄍv���n�ᱵ}��E_��?15��>4��������V�M8JKS������m��O�]TN��C�'��s>��M"�b��������ꌖ�e=7����-��5+4�1��}<f��`��n$�B��l�^�X�PYR�g
�6U���Do��5���W��ڼ�w&�U>� A��~J�g��H���%ʳ(+�l3�ҝ��y.�P���F���2S�sk�����W���J]㓜jL�*���+oM���O&]F?�|ĕ:8d�g�hQV����FU��m�tE{�gB�?ݾ�Jį�Uf���i
��;N�v��̥���YN�x����s�ak��[['��}_��z+z����wu��SD|.��<]p���/��It_,@��̕��l��`&Α��a"O���m�}arj�@7a�����)!Q�]��M�M(*�����k CtE�z'�(v|�]�-�(%b{�U�T�aCA#/���7��+����%�lĸ�ɍ�v��_������.
���^~�f��7��_�����J�(�/�ư����Bw�����2 K��_���bF�F^x���\�({~ȩ��7
��)�66�o���W	7��NU��
��^Z�Fr���e��]Y�^Y����:��F	HWW��Z$Tu�kVV��dn�xG�r�LL�=���K�f9&��䝏p?2;\�d���d�Z,���EiJ�$��+�E���-z�鳍�	=��+����f��;�W���W��j��=��Pe�"�ᔯ�F~R48e$�����*_QO���4j �iG�UΨy�7e�� ��]��d�*F
�C��\.ZY����3���[53W廬�0��8�Α��쵤w�"= �'�Q�n@�h�p���Y,W����G��z�L!ȫ���t.�Ͽ���!�k. :E��U�7_ T�����P��6�ࡤ�b�W~CI���K�������t��X�K<��\54U ��ި�{:;�T��X�,g�d"{!��O���^R#M��}�W�
YN� T��R�4'��2��d<�O8U;Fz��(=Pp���`L7��{K�{���[V��c<��/Z��L�s+{/v�_T)���T�X�Fl�:Y�z��sX��O*�ϼ��
�a/.s�R�@�����X��#�;)��<x���~��qg�"�:W�Ȱ��x���pB����� � 0��>%ӧc��������/�3���X���D^�-T�t��/�t���U���ڵ@��,gzj��W��O�unE��k2:9��(-y��p'�{͆�4J���_�^�Yn���I�vԳ�����Kb�)8�ȗٱ:�f"<+,d��Q���iL8AF֍˾c	x��O}�ʥ���j��K��o�Z�=�s#��]Ȫ�j��ײ?ǻ�o��������S�giy��T��.2lmfze��Q�涚��F+���X�.�*�|��T_G��X2[�n?��U�����F-�'�fz0���=Q ��ͦ�E�R9/���u�~&���2	*���q}���)���ȅ�sx
\ Ns�8vVU��6@��oa�]J邭l��)#�8�$�����.M9Jۅ�IH�o���\~��+/~��Y����ta�j���ҳTn'���8y�d�x�ռ����,uu`t��F��`�R��ZM[gSN*'al�#��]g���rj��ϕqS5~��MK�4;�:�;Px��Ƥ��L��z�L>)�����,���R7Ss}�z��R��͝B˒�6@wP�+��������0N�eb��#dK`�M��I}E��Lvgm����*Yz���?�Y�py�
�{ź�u��/O�*�ܢ>k��+�#�PA�wLyJ@5��,�|KWc5��V�-��{��z�LO�N�Ֆ��T=�{��l�����מ�\Y��K�O4>U�^�V�N����<^�-	,�������K&6�<2�+�zL�1\/jM~��ܩ��0��Y������y�������z�2y�����M�em�6�Z����GU1MK��U�Jx7m���u��3����@���`q�_}�BI
����U+p��Kb�R6rY��^#�v�͞��8`7��7�Կ�.����L�e�ߥ7��땂�n�f�UR��*s��pu?�ω������)����`T�WOS���}?QoөM�X��G�[GE�}o��VP)��RRQD	AZ:�c�!UDA@��D�T��n��y� ���]�Z�Z,�?��s�~���}�9wR�W�,�ˠۛ��&����G�"`�P� �>�Cw����>�[���^36���W����y����F�afRO�i����Xj�3I�o��lu����0��{`ڋ�zj��>�I�͑EN��+���7�&��Iw�Nɉ�B��~�o�|t�-_?戄�v��e��HH��d�e�U_����ӕwB�U�eH\�tU����D%v�0�EH������,��7=g_X}0�n�	[��C�B����S�'�{�2
A0"-h��]v�����m����E�6�Q���p�U��	���a���������r�1�ₖP�l�;�y���1~�bI�b��Z�X+��­~�M���%�t]��iv���v/���?|�ǲ�k��}0}�/����&O '�u�œ�<�l�#�R�G7����y���_Σ_����#�LCi��ܕe1K�Fl�5��3�*��L27���9QZ��+�L�RŁ�>��0�:�5��4��6-I^W2�I��"���+�/�1�%߿���c�G�������!�x���N�f��Q��ؙ��=��/<��b�-!5����.�p0�~p���*-�C��V`��8���`�C����Γ�������z��_�A������.��K���޳�V�w
�A��Vя*���p���2�s�%�6�a�ز�ӡw�~�WÄ�����?*5)�7<1?������d�P���x����dw(��T�� ��,X���$}���~�<�?�q=�7�Ӆ�/�IN��09,�_�?���߁�9�@�A����U�^�Zr�}����E��G1�n���@�'�;�8�o�!�����_ʃD�͋�@V]iߔ:DZ�-͆�v��b� L�8�$K��:j�;�Tȭ�R����9���?muH�
�"~�[��"4���Hq;�82J� p���ڶC���P�$�}k^'���ݓ��<5}"�W��W2��uf�^Uq��|�N��4=�&�gp��h�+Vo��V9�ٵ(�I���+�];�)��?]*���'�_\�Y�<�K[�}w�F���(��A����%�b�3���ʠ$��;�5�"_*A�(���Ε�[q-�%zS�Xe���P�o5}�o�7�crq�;��D���`���)Ef�o�kt�������:T��?���%6j��LP;u�WVB��q��K��9ȭ�Y��\?�J)M���c%�{�],"Pl�M��n,�%V'�z��OTU��_W�V���H�?rH��'
�T8#��3qq5T�{���ͫٞ"d�A�t�����*N�QS�Hc~�n��\���	� ���X=�1��xg}F����(��.��;;�DrXBz�u8@z(0<���̓:y�H���9Kf��>���~���r	h���[�*�~�����(�J��J戛�
��������&94����Nڪ}����Z.:��7x�pd�9:��zX��0dDKz���~C�˚�G��U�GȽo���Q�g�?v�&��[R�}x�����s���̵��c�/�{��������ݚ���1����v��_&"�|���+5I����_�-J��i����2��Ǉp�	V9}xO�5=�X5��pl�}"����|�)p�(f�{cX��/��5_|s����N�-�[�ooa�v:�;!�I{\#[�N�P��LoSm�0@/)/'�I	��Ȥ܏����:�*�Я�j��L}��@cM1��1��S�FK@/��&X@W,�œ#j�{.�"�$�Jɰ#r��omy�/���	+u׆�:ҋ�?��5蔿^S���
fJ���Ͼ��s��*Y�b�b�0m,T�S 5�����N
���@ORG�XO��9i���0���G΂*�7">,����֑v��������@�����r5����}��K���ͨ�?,��[Y�0|*�z��s��u��O�{H�^�e������ �5l"��\,���e-=qa�7��|�]��+����J��XL�0a����R�n���-�C(.2J)�� �7m������>c��g�^�'n�b"׼s�ɚ�c��3��7]P����=ZyȌ{F��/ɧu�S�We@ڝĚ�i52��'�=Q��maQߙ$x�Xo}_yK�dW�v|��o"ν�_���jE��ܠ�Q��GZ���:�pc�,�]����BRJ�I��B謄ui�s��F4�
v�������0z(�4��rқk��"�:A��I ��YI?�-8\��c����YH �27+yL�z�|�h��7��z�rD������_��S#Dɓ=�{�4Y�u��?������*�j����w A���w�
YG������g�¸8_؇��{+��P�w̐3�Iq��k'5��چ�W��CW^�1��rP2CP:�Q��X&:���Q�G�<U~I�_�K���������E�<pzs��S��<a�m6,&������U	������RM1�ֽ8a�8��q8^M�xh�D�CR5�$W~��W���?!��V���fy5*��)�~L�KuSRn�Oؓ����R��H�t~Z=AnW��)��S&i�d�6sk��h���1N�'#Vë��$�54��WƵ���(Т��M#����w�{��Ί�����Q�OO��z������e><���x(�H<0C^nT@�k>}��`�l�@�����V {tKQ �VQ`z�X缦��-ߢ�ҷ����M�>�p���:,HۻF�;y*�1<����B���޽��g"b>Y���0<?Y��{N��"�U��y������O�2M�Gu�V��)�����~}d����:[��7(?	�T��C��R��@�t���ڰ������}��́2�2�|�[_�+��~���5��8$��M謎��Qe�;�q����!��1b��r��O�F(}��}xeܟE�d�y���/QV�$6a�=�����_yxU���ە��bz�.G�tBi���
�W�XݴGߤ[�"`�EB8�~J��k�h�?��ghX�Q��!Ng�3��Nٱ��U.���U~Y�fO���з�:��h�!Xg�5_�1P�LA<�}�˩�!���F/�uL����`�gI���S��X�j�����5ź{ ��HC V�ȓ�ޥ�N�hǥ�h,� ���Y?�Ey�^������ۍ�	���lZ��u��S��zӛ^�8�v��:�_ƽ���@Sb�oNWRA����i|�蕎x�7����W��R2+�]����@����Bɶ���x1k�*�������x�:v���'�Nw{k��j����:���	�R~���K� ����1k0(z�!,D�)��w���<��"�7��J\׊�L~����s��B����@p��I��uL�63�T�h�+�"��h�I*'i���kR�s����xo�a�R`Q|�&���V�)�41��l>5A�yޜw/R:�F�1�S����N�vR�HC��t\��y��VE|[��
|t�����o[���#=�)PKh��,��&F���� �Μ�f��O��(9�'��[Oz�����5'��C3_�d��f��eߝJ%�����Z�Xެ˸�R�����@�x���Q���
0dkS`ޑf���ݾm�S�s��%A^g�c��2�1�meV�"�1�qf�v����j,�f���F�%b��)���8<���HS+CLVoC���_f�Mo�74���T$�ݛUxR����;$w�mx���\v��C��G�3?�v�#3��A. �x)t��_$Z�@3c0 ������9�������4���A'�@���܀dz��}�Y�7�*7��L7Ĩ"�;�e�J��F�:Eg�4�v���S+��Q�T,x��tv+��,��Ӊ��[�f���9\n��Ŗ�����DG��W�0����f��<���O:�F�J�p�$G0�:lM�	�M!��r�JzY��wAῥ���<�ڼ���"~A	��u:�VB*}���m껨�g�	/�Go4��ՉG��E\�?`��wd4V
�C)-���x�0I��K�eB<Ü�#���$��ώ������?_�w3`��Ƕ�(%�&���=K<��������h٫��/vew��_�u�|7���Yb��-�<|�a4�1�)�m�
��/���f�x[������p��
�ı�]������_�y��0�)3Jx���C?6�[��ޑ�q��
����n[Z��8��o��:�	��h����ȏ��K��ֶf,o�W����5J/��ٛ��u�?^���p!�,_-T�@~�N;/pK��>��^���l�BtP��[O1���(�v���,��9����y��9:1r2?=��[�)�'��+uٜ1��e�2C�{la�v�ߟX��Z�y-�YT�󺺇�[x�q�珠=���b����)�a6���j�R���
T��e��C�F5�9�Vw�NQ�ɪ���1.Ƽұ��Y�B<v>����q��S/�(�����}�~c&��;��"�O��� �g�~p�l��X�"y�Jü�^`�w��4�p��M�N���AI~��#s\ڸ"c�m~z����H���"E$e=w{����dQ���Cl��[qm��ݥXI��W�����X�VuI�X�V�u��m[�9�&�e��;W�?&>���h��?��_�*I�78=e>�|���s�	�B�8�9�� 1�g�s�u5�Aѡk���j�#��N	^��.���L�P����c�+�:#�6K,��^ޖڮO��"�"��[���1��Z6�s�0����"��:m'͇�j2�/68b����`�����](�9�#�#s4ڸ�UX'�����ee��qE~�zc��网cP-�����}>ъVn���N�`i41�n���.ԹXW�H�+��0>�O���_Iܵ��k�,�.���9cp�o�׬y�Z��V>]NlexE�
�X�}bW�O-YB���a�-�L�P���V�+�󭎩�!@�����=���U�����*�]`jM����ў
��wu��ĢR�H�j>���ʛ{3�Q��;֦�w�8Jo���:5�ɖ�k+�]�7��9�p��5��ŗyYQ��7�xe���J��*+��T�)�1���U�/G�{:iE�YJ/�3�V����e�5Y��C/a3"�,����%�ߐ3>m�BM�D�wD~��[�IG{��������[Smd~1��E��T�07/&�kS@#}��Ӄ����ra������f�O����i���K�AuÓ5�2�^�V>�����������F-�!�G6g�|������EG��jP�1mPTӞ�&,���y�{���94�Ԡ�jl?����s7�|�v'緈���掃4���9YRj��)��_E1�%���g��eTd65W��~�	W���]���͜窩>�rvg1˖�V��ޭ> @�]�B[]�Z�S3�O}�� -��7�\?��q�'G{4Ѝ ��y���>W��6��#ϧ�J�(��� �`�I��*h!P���ޙJ!��p��;)��Wk>��eЇ��W^�apn�l���D�{�ܜl\���fP_�h��Vsy-j��"X���_�L�Z� �h�9�{=VP��@T�2=�s��}��wz����Hg�������Z���2M�����9~�
��U����4�ߘH*0�'H���0����Y3ܴB1W�!��^�÷��砒�1����e�3ы-��OmS�C8�[�~�p-�Z�RR��wϡ�����rǡ%�G������|Z�=@>�e�����6��ig�0�[�c��RT��fw%���,P>�+����^[7V9�R��UIP`�}�x2�=Vbu\չ�}���*`���Xh�~`m�b,�
z���''.��>oh�;��Wϥf�XpzbR<�������\Z�D ��,��c�����l�3#��y�N�g5�.�y�vqE� XmT�M���9Yb�ƌ�;��h�HJ|E"�y�Z���$b[qr2z�5)�$`���x�wWk%����&���é�9 �0~�/}�(X+��gh#�P5��di�@����5�Oy��8����f����t���Rb�rKcѷ� ����>�hؤ���jȥA��+~U��<*g'Ն��0���*�6��NB�]���.���_,��5��}�� �'z�l_xu�ָ�-MY�������W��PH�h�����>5b?@sf��]����ٗ�i�J=AM�N�S�>n�$ӡ$�R(���ICąs`nwL����*��R�:c/^82�gaA��O��:MqM�eA�.$��J�P����0�K���z���`f�� r��˿d�u��	L��f� ^���a�e�#
�u%��>phYYBGU�&V�
ڢ�n?���u�nP)Ծ�yI��|}���Sy�l�)��8�u�毲/A�O!�Z_��-v�a�FI'�R�fڭ���:D�{>x���������Z3}д���3��wNab�i������_]ޅ-��:[ʮj�c!{��Q�L�A��zs�۷lc��D������Wա��(Ekh�p�Εq������:�� �N}�Ӽ�%GW��ق&��F�J`Z2��Y+s�pu��|�R����\i3�?jD�d%1s�&���O� �7ۨ�m'�U;�ټ���%�4�D���64ّ^�g�e�E���T�����{�L�^�3c��S������'Cb�2����d@���rdC�fx�����e,w�|	��Y���.Io��9Xp<)�lp��wb�r��n�Gl`�e<X��n)����-� 龜ص�w2�_qF����K4�7N�x�� ��b���8��8�C�'���H/�� =�m��k����Ӌ{s�? ��_��S��ヨ՞�í��n��TQZ��:�~�3��>c�=	H_����}o��q��҅*^+ٰ��U�ܱDl�y>��O��g��UlC1�ݱ��e�ZgM�&�H4L�x>�嚛5��ѿ��4�S`�����nl��S*��f�>}��wt��]���36�"#�yO�fsk!!�6ٗ�*��h�=9��[��-���^,7E�������������&�H�z�������,��|tr,2�]kŦ����R��<^���U�!�x@̲I��I�3YQ߬Q��5x�:ܰ�m����^HJΝU�ȘO�# �G);�]|����Z��L���-E[m�v�A��w	��v���EI&�V���^b�1��+)�g3)޷Um�Ӂ-=�E�+>3�.o��B�o-i�޵E!k吵� ż��y^da����~�2��f)���Z����������s�KN�e����w��s �Z�0�X,*(A@�y�����u��&�����)h���<�p���*�`u�,OM�X(�-�{���D8�D��jS#L2I�a��$�?r� ��Ԑv�l�H��;t�ϓ<�����^(l�;D�����@�2���Li�"���L��
*ڡ��~z"�)��b�Ƒ���%G��].P������&a<<kM���}�5cЎ}g�1��*�%6��>q#R�5��)���!�����E$t+i���k�p���7�o�}�*AݻQ'��'�G���K�j���9���Z3[̚I�X<�=�XA�����-�����_>���K�D�S����?��[�*�5s=����&~�IFW
��j�{��p��s�����Q ���Lγ\QrZ������{ Tb�K�y�ɴѡI.,��F�VxdbY%�t'�����]���ED ��1A~��)��QG���ϯ�-*�'��e%vJQ��ԡ�! 
�k�'x����/���š�FQ̒����(���3�@�?{��0���w�����Y���am[y(�8,w�#8�|�:Ȁ&�g�Vv���pr��i��5"�� ��_��P>W���&D���G���:��H:�|�/�4g:�/F)���K�v�����l֜ĭ!T
��W�9�٬�!>O.��|�;���׼Oz��.�d�"��:S�{�g+Tv�@{s�Sĭmoq�*U�\�� %)Gb���^?��e��!,g)��=��¯K�#�5T@P� %]�I��-پ3`3����2�|^��7�a�}��Jܡ�Y���!׀�دL�R���jU��lG��2�����N�F��u�|Ľ�@n|̷>V�y���L_��^Uh��X���j(��:�n}�d{�)��t<���l��H�#�g�z���ţ�V�{�B�/�Gݖ�j�uB���!�r���Xl��~�ֱ��=_ג�8V�,n���?���Xֳ�?MF'���t,�o��'80��-�u�1ԑ����SzF���1��M�2�;E��|�2�5B�2���L$�D��LOh��Wb���N��C!�b((�0>Oy�mH���5��L;���^D��_�����c���h�%���ύ���1h/򺇦���`zc�v�PѦ�{��Y2��C��|d�5e2�� M4h��!�fy3>�Mq���q�֑v�mގe�=��VV;/�sH�rBr����:�$!�Y��~�Z��h�TO(�1���a�wov��x������_����zI�	ڋ,�=-V�v]L�̄�zl(`��Y�C���Rנ��<��0qS�!-����db�r�ҫ�G���
Tc�Zׄ���j}�3�m@����vr�.buK�8� ��@���')�ΉI�C�_83��f�D�يN��|�E�
$T�;ʾ;�z��B��aߙF�R:Y�����F�2)x�|�I;�����kc^qR�$�~4x�ZKj���a�Q�6�����$�����x=���fT�'�����r�p 8�ݞ���X�'�At\|��$��7c��F��`�����lk8���6����U��v�&X��-q�4(k�I_&
�g?�~�W:��e�|��g���1?���^��"���]��9϶�U0>��ؾ���F�@v�k���Ov����^��b�Za�����@�e��ۑ�/��cD��G���%Yc��T#�h+�ͲA���3fƀ�ĉ%�@O2�f�(�U��v��ZL9��n��vNy�Bl@�M��I�ݽ�ޓIIr��3;��3��bD0HS��ط�N��6�(���P{�\������fj+}Le�զY�����k\�����uZ5'z4�<�[R`�o��t5�B����᳭��M�Y�>u$D+�L$�-*rB�G�O�H��	���o�O�#)R�Œ}����]m2Kf����
[�W�j�g�Vn)ۧ�8�\���؍
�(	�A��kٞQ8�  ��zt���%n�RQm^v�݄O��#QBd/��w�K��.�	�e9{��Dz<w�S<�%�_�Ր�	�v���C_�+/A�A��t����/���:NLd��+:���W�<S?NN|����ʄ�}c=��31vS-���[�e,��K֖�V6-��Jgk�b��sF0�x� hΓ��Uo�Ks���n�Bd�Ϲ%:6������W�Dh�Rx+�4X0\^�T<XL�l� u�}��[�,Y�E[r`(��,X:��N_�p���ɳ�a��O��ݻ>��.-����,o���L������Y��=.l�\��>^F}��D�tq�`���%$���ΩPQ��Z��]��E��1�"�7SDi|��UH�|�GY�:P(	�0N���\<�gip��t��b��E-`3��X���g*1G�I[�Ү�9'��E��!�pSX�j����f�h���`��� �������BU�tK�0-��`'{��G*�so03^�E���_�ꆮ��>ڕ�����TP��?q�?�X�JQ��F$a�h�#�Η��.����8F��_��3p����SK�Qʈ��C׭�my K�0I�=V�0��_�� �F�����Y N��Fov����K5����jF�U�m|,���	�pse�Ԩ?�z���Q���h���0����<,�|��=�4��mٳy��SG�����щi �`b�3s4�L�R����:��!k�2���)^D�si�%�]��9?%�u�?�@ �6���o�ke�����gȭ�6��h�?�0E���$E<`��0vy�B��] ��ۇ�M�>�Fh-※�Ia�a�zO�-8�(}���/����#�F�tS��X�)����J)A��y:p:� �1��)F5�7I���
���������g�ptíTE��{h'Í�T�Po����<O��{Y􉂑h�脳�dA���kZk�{��e}VH
|_^-�t�|uR,q>�(4{i�e�/�&�=K�:<�v�܅�U%N$^P��x�S1�F�Q4OvϻϨ!�Ake#��U�b�c���&�3+)�F����e;�s��j�[/ZX���ܵZU]�9żF�����nc�Ջ�'���[�J�g�&�"ZO��ٕV�WfτM�L�Z��uܮ�e_6�U2fqu}��Cz�&���K�hy�r���k�E�		ے5+Lh�MÑ��e��Y =�;�$��Q�?������?��|��49 \�m{V6ʮߨ���~$�%R�o�����o��Y��P���ӕ@����T��zC��f��Ͻ/����5-P��X�dBf~>��u�~w{\�s��P�½Rђ�yQ����IЩG�Y��|�7'����e3Ǟ4Q�T/
�ݚ��F����i �
0�ʣƳ�nqϑσ�d�1�%t��/���7��]��i8�b<�X+k �4z3g��'�Ɍ�E�����Y�Q�$�_]�`����2��꣹��˷�<���b a�mi��Qm'�A�����b��a�Ϗ��w�g��QqXr��T��s_ �����c/ஃ!=�W�ܼ\�"70vy��3���0�g�ٸ$���������d�Sϛ�:��-c�Uf�,���C�:����������|W;I��{�i{�������g�n���$~�/�G�?Eo�������ˮ��tg"@��^JHyEY�]���K�*��\��5����l�}[-�ϖ<l��J\>05�/�\k��-�����؝���䠐Թ�]�s�4�5Ņ�kh;=+¡��^�G��nu��N�D�T��~��~����7�z.�dF�qL&j���R�
��,T���k7�KG#:2@g���}&�z�5�x�U�m�i�	&`�l
����efa������+�]Y��1a�qiIv��^��7��u��$H�¡�xʁ7�;�8)E�V�E+������T�i�^�
βŻ^�&K�b&ׅ,r�$U_�`=�Q\�S��=KM�>6��h�EnB_����{ұ��W�uԡ��~��\��d�u%�Fz�v��v�HU���?�`��Y������ƁQP��F�������S��W��#qe����\/�����D}n�����*�37d7�ʕ�x�uj����ݤ|�P���O�ub_���[Q���r�n��Õ���]B��jH�;ގ>ߪ�L6�y��i}��s����f�G�Y��{���6�'�T�q��çvo ~��\:;y����cqEd��f�bz�B�p1��U���{Y�}YZ,)�M�H�y�7�cRo���sD�q��"��z�q�x�� ���?����h�V��{�]4���D*��G��������) ��e�Ϋ	�ل*ɒ����ؿ+Y�*L1�H�/�Q�O�9�_�@{U���1�޳\��&�����a����}0���� `������4�LX��#<E��EK{he��(-�S2Wj��B���[��>�#l���ߔJVB��ׅ]V�)�FD4j���ጾ���T��^��kw$d���4�:���_��	�83�4�5B<Z�up����,���1�9LQ(r�^MV�WY�)P�j���>b��;d�[���T65�� 2JV�K�3���8<��H]>���r�1/ ?n�O�ر.�����Nzt����R���O����W�Pn3S����m��]]���w�&��?���3*������%�5@��ñ�Pe�%���a���Z�5���� "��O����5C�E�B_a ��-rZ'��zMuH*Ƶ�=+�:K����j�y��g�o+��у=����iB��I�a@s����hϏ��Ƥ4��v<Ky��Θwۻ꧓��z�Fp����|Y>"������zn-Y���WIw��+�c�g\ _Ť�rLY�k{���8�B�����������d�z�Kc?�$��[R(Z��9R=zz��Bww6�B^l�\�!��U�� �;�y�O��w˛�?��<H�e�W�v8�K��BZ�A�wtf�;�@eem�����_�O9�.}01�*
�RÌ�,Wj�sJ�YJ��К���)��]L�~��]=�����w�}���Ώ�O�FW�}-���L�����\rpH�2��ր��+�O&����y7zC��> +ȃ���g�&��V�HV{������p�'yU'Q}�k�t�r?�}T7|[&���P��$�$��>L�'�<��
�(_��߯�S��KS_z)�ȇ�GP%FOߴ"�PF ��_�H3l�K��[�I��p{�%�n��.2��p�����١8� �t��E����c��"��ú(�mhW���--�TԎB�@j�����0�W1	�����x�:���n�-� 1�U͡��!�iYЮ$���ڱM0���X�����h=�
@�~�{�jf3}�w]"1��j�((��D�~#n^�R�|Oڠ�=C��9���Qꌕ0��+"�z����'3sd}��Xb���?����I9�u0[̸z ����d�����������өP�i��ux��R�a��O�[��
�񾺖�w*�z�
�?%v�qL�Ƕ�DP������B�,i��E���>����k�Y"q����?Kó4���E��5��I^�8���^��.2��ho<���ʞ|�Q�r8�hem�7M�zͬ��zl	u�������M�ǳ�u�d+V1���"*��ec�p$�����d8�348eyH��J����J5<ֽ�jrk����<�Ӓ�	��U[�t���M���Tߺɖ��A���k���(2�p(<�	@�ee��I�M+�����(���_F�,���0�p84з�R�e�t��)6a��3|yK�y�o�J����b��#����,����@�?�k�2lО�_�O���-��w�բ��u��$.-��⾓&a�o>C�/���>0��p�o� +*i�F��ҍ�"�0��B�~m��i���+*�#n<uc��&��ߗ�楒����//�A�wXR0��w��c܄��=�Q͇
�A�����A��w�XcX���+������������V<�n�t���7 ����X����s2=���BK�,y����h�l�0�sզW�����C��Ä���/�t�R��+0g��lar�gկ��eiӽ����O�q�mk���v�<�<�%�<�hy*-�}Mk��!�V��0�!��ֻ������k� A�eM����<�?�!�>3��Gg�.��X�&Pr���l�'l#U"vt�Ɍ���^(]�N�`)�����oJ_ѝ�����`�Bn��{�9j��c��T24x��L���-FX3R<���^�C_������0�Ӕ[���9�f�Gy�78�2��7�k!4�Z��酆�Gi�Ҝ�e?��/� ���޽����`��y�(-����h�ٟ)�L<��0��]�8]��f��U@�J��˦�~�d���o��ԟa��)T ���}a�w-��3���F��L�A��]�yo�Q~Cl���Y#��x��S��h�\%�ً;+r:,d4�*
X�tM�
�tP�Қ�\)�
��d��l���Ʀ���/k@a�<���p<_�l�NV�l�B[�
%J�����
�x�tz��n�o4�`��FϚX�)ZʶO�34֮��
=�~�e��t��r�u?.Epܣ�خ�P���U��Q��<�N���;w�\�ą��a������A�~�������NaTW���T��p�샳Ǡ�a��6�/�gI?(yf�yOV�ZD}����Cy��ݜ�I�����5n����e(����*V��ѹRɐ��2�rFg�s��ߤ?q)�	g�;���0�2a��&'�g>>�ٯ��S������C����(�;��=�ҡ����~./]�r/�'td(���^~�y�a��$6���!'���(x��n�8נ�������m���8␝"kje��Q�z�$���UR8��L?���}U;u�f�|��'�	5��,>ڒFy�L�{��hIJGu%E�06t	/Y'0�]���ݻ���D?Q�Lhu���=�g�8����<��ey4�3���B*����	��d.�[��������66l+��������-D��j�}���h;��X^��3㽹�#c$6����͔��U��<��~쵘~��ߤ��C���q�q��q
�l{�%l#�������猻�R؁�ԩb��~F�¨�A_@֯JOK�6"AZ�m���'�q��u�Ou��Z��?^�>�l�=(6���Ƚ��S�#/���F-�qȚ˰��/� ��w�,��{~�,�Z;�!�����(s�K�pv��� �?wI�A(n�1��8�M��d��\���P����v�W�G���0ه���jyz���fF{�I�M�dB�p�/�����"+2.��L�ͳ������{#����t�φ!<�cl�w�T0��X���h~��-��n\1nM �t�]p�~ YTgs�F�1�b�'������h�J�<za �0}�� �-dru}��e(Mw$l��M��F�:��$�|���qQ(�`�v�Fӏ�'L�O�ʣ�����p����mh)��ign��<�7��٫ҌF�Z_�4"Lb�,��
C�����u����3��9:t�Z�BP��h���Õ�2	�=h�Y^F�R��5�޲�	�ݫ�l�<���Mҥʻ���|�O��cK�!���sUe�T�_@w��
�H��G7c��V;r�7GЇ�PH����(��T�
��E#��"��7/4P)"��;E��q\H��z��K�e��u(���ti����Y��b��?�ɸ�c4g��\��o�ބ���L�n[4�<l���(=J��B��Z#���	��>�<[V���QY��9e�x\_�h
�_�8�ФzO�{�\>&k\7�ǥ�8/�FK�=:.�%�?0l����=N�/|��s�,��F���kZ���拫-���1�Ay��Y��ppT��G{��)ǭ�2O��w���'$�����D��u0�Ro��F���`���5{G�c���}�|�F��s"C��S���	#גs�R��Y��	9E䲲--��������38a�&����;�e �#���L݀�� ��j��n1�g�s~(`�
���L�>,��ѷ��E�'G��}��!��!`��;'o���_��]λ����Z嗵�5@��ſκ���.�NGLt�g��ͼT�`iݍ�=��xٚK�T�-�	d$�Rv��������`�W�J�����+R�~N��o�]n�<Z���g�����x����@�r�fe���̉I	ј�it�Y6���Y6_cOy��`��Q�����1�f���ᎏq/(��$1P>vc���O�����C��p�.Ӱ4���Pŀ ����"�#�in���F<�ү<����H�m�����}\�������
߅�H��Wq��kx�N�3O�t�i��6<��7���r���/O� ��5H����D������vS��M�Iq�y��P���l�9d�����p���,)�Xޤ�ﱡ�s��c<�I�Po)]Pk���
L�J��{�^t�y7*Yv�#u/��(��_|U�N!%�)KJ� ��g�UZ�{A�j��M12�_�8%�?f
��ԗ8S&c�D�i�@�*�Z��M��V�b��_'�7S����PY�3ӛ0�ú�I�;m���!�f
e��S���#�x5��%�~��P ��� +>&�oX�\_M�L4��{
	ޒ�Eܲ��� -���sV��V����N��j�g������[��X��s^���o���ը���{sw� �<��(ǉ<F5;" `c)V��`a-��pZ	C�fyWD=@װ���� U��9�&�x�OR�|��*�!~틄�s/�Ү���4�g3�
��9-ұ�F�-����h�B�v]�g�)�v��Ȫ���3���}��)�L�h�L��K��_g�{'�8w�{��q�}hR�?���Y�H�����VC����+M���I�vߡ;�ɭ�2l����|�rХ�|6T�J	���2�!i��w��������b�pqC�BU�2q�x�/����~2��N��Ca�3����S}�� q��{��,�����0f��B+1��Q�<��*�N f��1�U�yj��>���sl$z�@�*������i�h5�}��m��<�x�/u��h���)t��9����
�t���b���d�3EF9$S���c�ISxR4E�pH9n�����2ʑ��8r�PK\�����<�aխ[�E�9��� -|�1�&J��p_C5Lԟwh�ݙ�X����i���8axS^��k��]���`c#�Fp����'�VΈ&���>��b O������㱝��OdƎk�[l�����q��O���?駶�k��`�#H����p�o�������-�S��HDa�`=��S�����]�zw��l��;�p�JL���,Lwr�(���X������LЍ��O���3��ih�t��%BM���L����{"�ຍ�z
�~��OKʊ|5���+��Z��}��[�b������^�zz8��WREF=ػi�`}�q|]�|�����"�w�cO��E�o@�����7�c�S��}�73���_F0q����.�(��ge�}^�U�+|�Jn�v��rZ��!8ꟹ�Da�ގ��p�ΪD���;�I<������1�"��v�T�L���qM��.J����x���:<����^M�]�q���QaT�� �HA�n�HWi�T�5���
"MzJ�JP)�Ez�$@�B�=�2����޵d-��$'���{�'�	M�_XM(1>�� =T:�{3��m3������$���G�v������2E�����0c�-�[�C#�rӅ�R�_�[���/��I5٪�x!�d�&�Ύ)ah��M ;H�ޑ���Sۡ���/-\����߈�9�R�p}-R�1P2�[��%u�p�C�#�D��J~��B+��VMf�(�H��s|{0����/�.�m2W��3#f^H=?=qH0o<Ua��L��[������⻌��*�f}��<h��.����$n�M��5��T�QL��]�����}p��և�K<Z�ɼ�&��]�J�اT����^7���qz7Π��\]R�C��D�#K���p��I{���2H��<BG	߃��á)�:�����aIó��j���|�zh��ղ��R�v#���4��o���|�9��'�.�d�`�a��D�h�۩)�������[6�ߖ��}Ѯ�^�%]+�� �+O���=�����o�X��v��?|�ƪ�)�����!���S!�oFo+��&]u5_$>�׷�}ߓ��`o����i�^d��4y{ڜS��y�
$����G���ѓ&�C�Bg�3
e9�el�L�:_l��>����^�5�?��q��f� ��$�_a�ߞ��n�5)��~c�>�Ѫ'��U��J����ѥ;q􊐎;5vhR�J�by	�N�4(\X���`��I;�I�]@܂%Md���T�3�2jE�ij2����/��pV����!v)�O%"��eRA�É��e�iu0F���HW�U��M�7|Kܩ�G*���+�����5�����^:{	0NY�qC&
?qyo|���׈GWb�iAsz��=����臙�����T���F�i5�W!�y�mr�> ᤿sa�g�M�me�&��V���N�I��y���W�%�zG������?E3_k�ܙ�J-%�Җ[��[{��Y0T�E�2�3P�┌U�i�C�9�|, �;��_�n&}G��S|��`�w�i���p3ǭ)T7R��MUuB߃���c��6E�?H������B������_�x[h
�Ȑ)I�Ǩ
P��U��xz��s*|��ы���m:#>���/>���T���}5*ݧN�L\��|�C���%�0��))*/w�Yt����#���B��B�2�=u�G�v��T,�0�D����?bN�?��O�CG޸'?>
�˭�жh$[�Y�4:Zr�B��_`�EDi׹���ѝ����/_Np�LŊJ�M�h;�]�������o�Ve��6������H�'Ӿ�B�#����[zw��4�j|��У�� V�F�P`�H��R�i���s��lg�ZM6�0D5��Yp�0l�rv�咫z�0�E��W�?�Ƴ�V���8{\��n<歅u�.�<�]]w�H�)\�"���@U�?���!��x*1e34�K��V�R�z�-P�j��������Z�g�܇��}���52|P�3[Vj���G;6���h��[��{�-%%m���ΓIߕ?ԃ�fr�Bj�]���C��-���@��e��j���4d����b��߆RGK�_l�}��٠YN��^6����؍��I��'����������{.�F�g�3/��{;\��Ү�C��(�x+���N3��z�;��e� �x��^� �T�k5�~"b�D]i�'W�&�y�c��5��ª�O��[wbǆ��0+�kꝄ�F*"
,�W1ˠ�NxX��v��0��:*4#�UU1F~��<ǂh7=�A�zh1%"��3;���ݦ��i�#���W23���3�oy���d�f
��և
�E�F�
�/�/P��Q�����Ƀ(jBQ~�̔�`����h��f�2�gx�O\�s��Ja��RK��򊳒��	01Qѡ#�#u`b*db�+�_ͨ�t������C�
�H@fu�B����eYv�*s��kNn�t]������G(���%e�	���[owE��6R������R�`gz�9���ֹ�w8	Ɂoi�+�����?�#�p$H]w� s�{o:@-,�W V��W?��SF6��5c99���	���C2�	�@�>���2u5ժ�ϼɲ��8^�W�݈�On��=46TZ�Dg9)�Ε�Ӑ���#M���Z(���`5lTK˟���m������s�)�<��y#��.�:q�':kD'�ų�%�=p�:�B:]���������?�V���5�	4O�9W�a7�ﹹ9�e _���ɂ�����W���J��t˄8��b��n�=_���g4�yMK�W���DdZ�]��Qnntr�����A�T��f��	
�>��3Tga�hܷ
��o˴Z�� ���@�k���Ew�}|Z����l)��FJ��7H]�o�`�/�]zM���([zJ���d�����1\�E���7�H��DB�h���ϫ��{�֩ސ}�
����M	����Ѣ|�Й3h��NF��؛���YW���ɯg5���썢��
���V�Ţ|� |!�o�K��ؾL��ה�}�ᢵ_&�������dR��)��Y�h` ��f,�	w_t �T�J�PT�T&�b�I�g�X�,<����_+쌨�R(�5?a���o@v��
��u���r]�bG4���G"=F�]K[��28^r�k�X�V�bۭ��2���^�@��#�(J�eڀ%5��[�륍.ҩ��l^�!k_/[�^*Ȫ���x�1�݇��9�����?�!���20�͗�\�V�\�'m��WIώd�KS�I�uN?�x��u2�aXf[�FY�`���'�8ot,^BL��xɿ���\#~�K���n�Vj�E�!g��Ɠ�L�j�S�^E�^y������~k�.(C�y)���.��A">��ލ�(��,�3P�}�v���o@��W]��U9���ۦ�Uf�I�0[W�:--��W�9�g�>��!a(�<~���xR.K��M����2������ʇ�G}5���;����C{Z�~�G����t��%ԋ�
��rzߍ�t2�
��Q b��<�t��.ˍFD?�}�gzW�����٥��f��f^D��9R�:I���Jo�4h�n��'�S�,�����1�� ���$g�-��w"��`'Ҥ�ٸݝC�{�IUS=�\H�P.,4v���$�EE� �{�4E�������I�pL�����h��5��@?A�֋��xx�І�s���J������+!�o�t�K`+١ӣ�^t:�%$�3����^��z��Nwy3|:f�\Y�2�Yh�y2a�f؁�y���-Y��VJ��J�-����X}���EN]�g�[�7��K�>R������� ��Run��m�E�+�uN���7�	�24�zM�{Jڅ�<s�0Ev�-�V(G�4�t��`���n7K��HN=8^�S�ZE*����"��̕��}��N�O�A+B:֌nC�/�A	��������h_�Bgcц�E-͙�hkG*#/Ln�t=(��Q//:PnTN��S4���$Y��L1���y�.�0�_���X
ʞ��H�/��'�����v=�H���p|q�GP��jD��Z=��Ym;t���`~;��qH��z�ߗ-!?�Z1�0bS��2�J��v��9��>�P~�#�0�6�&�#��4jav��Yg�!k�7���$�t�Zy����羫��t�0!���M?�7���*��h����A����L|-�3&)�z���!Ǹ���֮�fC��AA�^A!,Y<В�"�R[h�6�M�� ���{�$�9cCy�f�߈�<x`ad�ꏞ���>f}e�;9��0�e<2�~w���K�>�V��L0�dC{u%�4���FU:2/����S��-�-*�i�]��<�u��[J���#Lj���aX���9q�(�
���`|�P�����ށ�ε�J���(I�e��Vg�ԞS9�x>�h�L�,3�u�|.�'�-'�vE�Á��<\uCU��<���%E8�4։��k9V4�,�3�.C��&�����Bڝ�S}���}�f���V�w/_^����q|��~�����Vm�o����8�Dp�z�o�x�:4u=umبb�߮Wq�� Uf#&�a9o۶�/��^JD�*;�ӽ���̈́ݰ�4�;�z�g��@@�;��"z�w�HK�@9����Ex�~9f��R.b�ژ'������ca����f���u�wN�BF����J|�J�w��M�+��#�Bh��/�4_��mESa�G� �_RT��T�"��&�e��|���F�I�����N����902S���[ƣ\��x� 2*��\�|�	/���n,�lkʰ;�S��e!=�m+��e떚��%���N�1�]����2@m��P����Ҩu�Y*�h����e^\��vL���r�b�Z�CA��j����{�/��7��4}Yar� GzASg�c3��^�Ϣ����Iq���
M����]�~90�4K<�yT�����4��nz���d��I��	���\���I�uӘ�߁���g��	3O\^�g֪�T��RB
�c:�A���`+`~��.�WɆ>���=pO�Z��k�gM�)0۸T
�WB�Hx��ݗ�1���M��AH˰!�xM{���]|o�*��Te��O����IlG�R��f	�l���)`̞k������KxY��SI���6��@~M��e��� �	�z㩘������7�_��1U��g ���8P�{IӽQh��.��%W=����A's�d`��_^�$�ἴ1��*�@�>Ogj��l��� ��yx�r�E5�z��3�����3.����������l�R�������4�m�n�{��tw�R��hb�i)�1-3/���(�H��λ��q�������U=�m���p�s�3���f;+[�_��qH��� n��q�:���e@��쎺 )GUj�՗tq���%>H��f9H�R��:7�����̌tNT�=�9���aer�IϿ�����Y>� �����o��@�4i.8/<�/�N%|�4����k�*�d!��[���\��d�V�>��~_MZ�i��{K�=��;9CD]�V]��M�|��N���,��`��9�\��rF��lk��
��BL��� #o����nW2D#v���#��Lm���Qf�ќt��qP��X��K\kQ� ��f�h�g8�|�@�]�W���v�q���|r�"��f烒
43�JGZ��َA�>�J��N�>oqWih�+s��Q���`uY��xg�(љE�� ��3l*f�9j�=G�J�w����66Yij�a�t���zs�dcl��;%���d��c':�G"�M��:(y�������͍/~�x�8f[SI@�[�8��دr��3O��Κ<0T��,�Gq7�)=�;�  ܩ`�V�X3��(իK
%��0f��2ᬾS�oP��>��^ܑ�U4,�	-ዼ�-��r�u]����b[[G/��6�b�E��MA�K$m�O؄�lc��)	�?J���X皀�BAO��E��o��;����b�Ө(ic�hW�3��u�_��4������<����w�Za�9C�}<��1COo��W�uZ�C_������cF?=�Z;OˤMwH`���EL1ui�"|Q M�Nк�Υr�i����S�C�A� 	�{o3�ݺ��bl����E�F��p~��h+��=���0��i&,�S37���X��mEN0���M:�b2�28@���� �չ���M!9�7��ϕ.W�;��#,-��et� ������h��\��يv��@H3�������ϱ�f.2��"3����)e�[W��D�H�`�<�e0���JDE^��`9ϱ�Jt$#%� �~��q��`�6&���=�k�V&G�tf�b� -�o�[Y@[�_^�}l�C�
i�-��}���X��g���gm�.�K m��l��]#k�W�.@�A�|�N������`��s>c��N�>�G��oF����@�� ��3٢�R�&E
b#?�[��[����� h,��f5G���� �9��y����9��b�SG���B�۸J1��Ui'�(׼=�ӥpn���r�Μ{M�y ����1��}�����4**bx8�*����%`��~hb`�Xz�� >^C��� ?����n^��@��~ ��ϭ���|�ix�~�����є�L�+Bjxa�b`ty�I�����萺�)yp5͋�����Z��̱k����_��}�T�'���5�3,ɤ���/I<c��|4��V�ݿ�ecK[ӈ����@�Te���L)�$)Zz;��D�:r���u)�ݾD�1�2)���}+��Dɴ e��{Q��e_�|m�̦|Nx8�U�r�B�5'E���˵��뎣0ѐ�o�Ѧ�#��p��m�vG���I���?MF� k��~��0���\s��4� �:"�-��i00� ������ ��vb^�����������(qW@�O�!��쪁v��m9\��S�]��e����0j�.�\ߤ�����֕� �zp</+�������$1�`���q�ps����+o��Z��߀	�c��@9#'c�8���i\ۮ 捾+$�P�-�Y��p~�E
�ݮ��mE�}�Z���.���J�ɀ�{IY���G&'������>{̕��@�{��P�Ց8����0[���0�C5��A�nd�Em����J�3ٞΧ�Hefui�)��K�˕� 򃛉�!���ݎ������88$��$P�������v�i(��$�r�(tE�d	�_��F�\����Phow.e)4�
���+����.����լ�2uvI�]F-' ]�����0��&�r�y'#������� E_��b����Ũ���� �� �ؠ[�����}�Ϙ�J�ĳ����]X���Į]%�@%=��w6�ץ�B~�Ěf6m�O�!�1��G"w�2���( �Q�6j�{���F�\ls|� K=�~f��T�s�;��27�(�uQm� ��l�]����}��q�@�h���\�$E�%�L�5G��)�&"��W���,l�5���pSz�(�252�@��]+�ny�!�Q��{֫�B�Xs��Ԗ�,��x[�x�hIk9�'0V��̬H�I[�&�I��.22g}
�ccL��M��l�/[a�0C�H��̎�}[W�����;-/��^�y��h�mM��$&�! #o�H���w��5�J����X_����!��ii�Lo4���¾<S���A��z:|�i�M3lz��49v�TL�J��{˝Q���?fS�b��Lإ��Q�h<���6�W��h�R<�+�%�\
ۉ�|5p�o����Ӈ7n���NsԨ6?؅z3N�J���<0�+���wVC����҇�©u%9Qs8׿�!I@�twl����5�Ԛ@����6���?��x�Ixcɓ)��n�Ɂ�����@���3h%���(^,�VL������x�UHl��PBkBƑ��a�sb�OM�P�5H�8=ݩ|Ҹ��R1V��\�S��6�Y����hP-�tѢ9|���X��I���C
4��I⯗	y�莩,��$���ߪ�&s�7�=�!OL��ݠ�v�S�Y�ň�.�f)��EL��,N�3��u���gij�����+�ʎp��yd�QU8�+��=����<��H�f'���@��6ZdT�^t¾z9P_RH�[*\�+CA]��9�>����x\jfwy%p����eͣy�UYam>���r'L|����Կ�,�d��7��d� ��X�G��;����t�V`'�����i��ȉ�Rb㘬ѫwo��!��h�wmT����R�$�@�+�6�������MŅ�؁3x���/����6SA��;vu����F)�p�Hb<�r��0�O~�S�d�U���H����J����{3�TfZ�i�
(l�Bv^w��2m�yۏ���� :׊�h�����d��bYLgju��k�6֜����G�U��L;:�W�M��}�*��FMlP�4*��U��eD��Ao��^��Vڱ��?�&?����!�����i����̙^�rY7d1$u���h�J	T��@-0�jn)�۪;�����V	�s�s )^?|+�h���N���W�Q�ٻ`�v�H��N�`T^�����v�i.�ÓJ��E�"~`:L�0��:��n�@��a&6�p�s�u��ڠ7�j�a��[��bGٺ�9���� ܈8���E�e����q�k��{�B�o P}�׾QgEN=c�"\⡺(��(3�V�b=���[�|+�8{p�h���m���*m�N��0w��0�UL=��f�^ی�9����!�9/9��m�'�[�p��u@���{]w�Uo���9��8�}��1�r��K�?�z�N�0b)��B+�z�M~����3k�{�z���tg��gŅT���T����L��HX�]���Đ�NJ0�<��Ɣ6��j4�	�ȋS���?�^��[.�]�g���� \�P%XX���V�	6�E0`pP��`���#�j
�L��4���x�Z���lgB�,9[l��w�f#xN��`LI��s��9�ڽ��'�C�����1d��y�m)gXr���ǫ.�I1���-��.�=�	���4�-E���:�+�,�<�V��Kq^�-��|��)~���=>E��~��P�.������M]�$�qd��ӯ�O�!w�_����E�"z������,���L��ϣ"h��w�J��ï��D)�dJ����e��uo|[<v֛>��0J�#���k�?dC�T��%wB��C/G1i�=w��3�d�;[�p��I���U78D�]�[�,�t��k���*M������ Fgef���c�1'�^]�����u����7��;w�˹�� ���'����BOy�������p���	�%)�w2�<t�#g*6�+�h�?>{냯ϸ�1�m��f�i�@cë���E������0v�6(ɔ�l4>U:Q���{�H���|!%Ui�����ks���n��4�_�L��'-�����B�QO�eۼEA��*kk�/<���yϽ�
�P\�
fm�yϋSr+�e%�z�rJ!���u�O2��QUP����{+��5x�-]�����~�'h`�2E�5T>��HX���Jq��3Tc@f}�\R���6�̒��`�E���J�`�w żyvA��H�\(.��zF��S\{����� ���fx߷��G���%�x�+�V�D�v��MX�� !y�2�$j��rr�[ )��SR�����6�2g��vC���[����B�+��]��C�'��:�����;��S��7� E�x+�oP��R�ߎjw_�Tќ����8��K�x+;J�r���lv�}_��!t�
6l����3Q�@"�v�Q�@���U�E��{<vr�˒���`?��/���_�m��`Ñ�FG���OIh����D�_ ��gP����[�<�4׽���^�]Ҹ	�žbd�:G�^z�m-m�.���������Ƣ|����%#r�ZCPq�	�X�@��Ѡ�������K���1v.�����!p��S)@�^w�����H��O6x����J�V���70�l)�R�[����cP� ư�,��&n����>�,܆���3�:O>����G�W��.5���(ے �,r�v�
NX�a�QZE|q�W��?�.Zڇnl���l�O�\e��SSe7� /�zGb���[�8��8�a)��	 �A��/�*N^�]}��zOiw!�<�W����$�#��|��]ï���'d���s�dN�Q4�v Wj��*yMM'<5\�6a� E�Gq���0���Ygl��<�©w�Z�°,�\.�BQ&������S�����5���7�/5h"��S�drO�=������7Վ=�z?yc�p,D�_õ~%�H�)�ͺ��U���B3� ��ƻ�^�P���{�P�Z����Rg}c��j"^�Op[%M-��L�v⮻�^+j�7.S�9Q�����}��ݏ�څĦ�.��@�e��g������I��VHг���Ȋ��rk����.�ԟ��b�jDN�ښ�3���X�?�&w���g�Db�Q��Lt�ju�2F������M���"����Ӛٻ	��@v�Al�2�"���7�+�*0Nq�=��-�f2�b�`���ޜ6H����
���'��]�u��O����\t��?YE!c.E�lIH�OM�{��X��Q!���%�p���l���ZS
���ۀF�9�WtlS̴�^��lL%)gp�kU����u���(�x���fYE��k��T�����l�A��r"���*~�'Csz}�)�<48g�ĥ�E!��g��E��e�����f�<�6�Vgژ�L��I���c�K�:W�YV���n�uo�������.���i,]�'��	�>ϥ����&��>0���"�b+Pp9=wt�F�`����-�k*��wQ��S+"sW?��ɥ���V�'yAqƊI��lM�,2���l����h�c���ʧ��p)�Ť��~��~�d��w`����)Ƴ������)~���5N?h6����o�Z=�a�WY��k����,��5�˰��ɑ�����gI=�vB];��<EARb��ō`��1�٭��
Y猨�-U�D��>��̜m� �M��ܾ<�r��J�����Bv4"��� �$���
a_A�̦̳S�L���HA��k�f�%�h���yn�T���G����^�chc��I0��SLc��6	��i�wz=�Zơ#��&-9JR��:@�V;��S$�?�0J1�0՞�u�i��WO�߇�E����hKjд�&w��e%Bf}����j�Sm[oyl#V�{�	�#�Q�;}��VC����I���<i	T�E%e��f[�����傑�J��(�U���)|ޘ
��{ "���n\����[�����!+a�b�:����RH2ä��7�]�� ��DX�V�&��Ɣ�:��e2�9���!��ȿ2��&y)v`D?�4�Z*��\ccm��B^@��x��!0�����я1BڌX���Ff�<Z�CcQ���gu�沬	���\uB������p�칑�����)�W�^�����W
�i�VO���U�ec�ٝI=��C��X��1Қ�G���J'a1����ŵ��A<~�$<L�ř��r�c����_�����t��QR�S֋���2-踹gaI�EH��&d�����l+���	߮���a��x���ͅ�๿�~:�G��_G�Ck.ZA_H�~��@��x��G�QY�Q<:L��΢�<�)�~�T�!ݼTu���:i�3���R�@�6�@�k)融�iX���ik���V0��=?,5в2\��Êc�הbV�H�=���zb�ϭm�A�奢��b��������8g�Ҹ�����)`=ᔢ&�Y��EM�w�6W�`i#�K��<�l��|�0.�����1>�	���J"��kTs��[p}�Z��T�B>n��}�.A�M�E��?!�4�)�H�^pߠ��d�N�H���H6�VM���#�gP����.E���ڝ�]ħ>E�u@�m��pX7D !n��3S�Z\#Ӹ+" *L�����s��\/VR��x� ��"�R�C����C%7@������gt��ʜ��Y�/�͟�%�����:I������ǀK#��&$�]����"�m{/Oas���Q��7!�l~�lKYԁ�_oOތt-�&dY�!و���L�^��8q6�Ǔ�+�/�1�V�FF$�������y^����:���E˚�[@k��� ��7�1 �r<�0�jl��AYqr���f�L�sP���UJɋ�R�)0G%I����3+�f0��� ִPI,2?x���O7�Ht�"ĬgQw�ND�n̖�O���1�X`���l���y�d�Im�)K3Ӷ�
1C����Ff�@Z���v����
Xyh��C5"S-���d����7�p�h�릵��C���Ӷ��`�u�B�r5-�Xͥ7��xN,1�Aӛk������o�5��j
w�E��nW�|f�:�$��%�C D+gF�ӻ�S�,�3��B��?0 ,����.�as�چ-���
9������.��d.�`�yBb�,����䳌B��z������Ŋ���FF�?��5&�N�Z�Ī;��EC���p&� !���D��IGM0��u�[�h!�q\��̀�T���[
�Y��W�܏ XZZzK'e~�jW���E��5i��j�Y����@
()&D���G�E����iӛ����BI���r@�j?KKԷ�k�Rz@vC�-�Ƶ�	��ǧk��Voy� �����y�� &8I"�qk�ύ�����z�q1!Lo�l[��l�'jƚԘJV|5�*ԙ�ؽ�䆱K��4��q3Ԑ�G�Ǳ��f�x�����F;�E��t�6.�u_PS܋rwe�c��rq�-���¼�����ߥ��:��&S��e���%ʴmt��X)6^�7�5q���S*�BW`��;2;7������ ��K���I�9����<��YKZM6�N(�$�l��-����G�d�Hvu��+a���(�G&u�9��^,B2��i�rM�JЅ_͋T�����5%K��D�����NH��{)DN<JY�J��� �]���$�Ku��vsa� �m���J��|Mdw��'v���u���iW����4�g������䞂�����l)݈k�I��pcC�6���&T�k�hWEV/�,�4���Ո(�Mm���~���\z�L�i_*%[�:�!����a�pg)�y/`�@���	�8~�&0�QiR�G�_$F-�xIFh2�����/��nY�x�Y'ֆe�_��������h���k�=�Ƒ���\����;���N�Bo`m��D�F���	<t�ݚ�5U�]${��m����kl0v;��v�O͸MΩ	�j��D���&�O����!�S�l��Y�Ԗ�q|�%���˄��VAw�KY<f2=9z�~n����z	!�"l����m�QQ��ޠ�+4ù.���_�L�Gٯ;�E4�;�`�9''A�"�$ݿ%[Ppi�QXx�s�U��	+˜S�GBr⺚��;��-Z�m��֊A�}���`���'���a��~]q6���Y�VRzI�b�&L�#g�K�� ��u˵�C�d�Ǥ?�ZK�mR�H7��Z\M��%�śQ?�H*�yJ�a��"&!"�g,�Z�ӓz2�g�������&3���GN���n�7�.�P��v%{�A���/u�kU���y9�� 76}>x�����	��]��v�ô�m�Ȇ,�ֶ5��6����fu����Gt�\ϋN%�B��b���{�j��ݼ_(,�)6����]�&��bp�},߅�N���#ؐ��������c����qQ+8���a��PŃ�s��؋��1ѩܤ,�Ȗ?A��#z����\�
�.[sg�Buv�������D˿},����c�5��f��1{M�0Y]`X�X1ݪ��*Ks�Bڧ�UD�/<�miHh#��*�T",��fjz��(4�70�|���TE�D�����m��h�}����F�,FcE%����F�/r� �e�Nd�h��0ę6�J���L�7���}��=�Cs*��,�C�F���G<��m�xh��%CE�|J`C�Uu���{�M���Q�m$?H������RSMp:--�3�b�¹A=7O}���'����������u��.
�,
]͵�'�̿{
�l_Q�b���f<TZ��4�y�]�F&���Ĵ�<eAQ��p�S2����r�k��q3�*��3[t���93ٗܖaxu}�y�$��>�c�y��ٍm��c(�^rxXC�ޛv�ʛP��k�`�0㚑�M(�Ƌ�����+�"�೵ZT^a8�쬏3l�x����aYb�*�����=���FD���"sB]��z��p�|�L+c���W�<��@GyJ�ڎe������OU��&QNƤ�Z>*��'����lp��ڃ�ԫ�(�LN2�g����L����_u���/������V[tbs-�����8tS&���&ͼ!����s���P�Q�i����������sǏZ�N����mep������m��͙,�K��﹪��($�2���^�}�ìbc����ɨ��\���G�e.�b�M��FZ�Sf�r������>��S�0ӯ";��M�v��ڀ#���#��;A)�/��6�]'�D����!�Qwv�����mYzn+Gs̝�J�u�,,Kpj�I��^9:(�[��`pin���{֑�*�nIC�5	n��1m��O��U���B���i�Z���ք(���Ֆ8��Q�ַ�!M��jV5�0�ײ}뇧iuŠ$+Նb��=��g�P�v9�'s���^��{�W�{�
�#�#�:Y��-]X������Es��u�e����I��(/�86��D��$�cRo��a�B�a�����D��7��1bի�aꏧ;�O�dSPU����6��6�������u�j���j����8W17���}���և�:n�R�fTG�d
�t�w��d�åֳ���ܱ
eڭ�.���r^�7���}ϊ�vb�!O|g�'�hJmլ�0M��:��,�}��QB�_�'m;�[�<8y�{=9�L��_�<�^4�Z�u�2�K1^Ȭ|�e"n^1�ΠOA?�Ro����n�WnFL�]>�bU�1�Ǻu͋��U/KRh��u+���(��l:����o̘�_9�����˛H�O�6��3K�0�M�tOi��n�PzJ�XhޜҀ�[���g�۫��=5u����c'�2}�:���f�x�;�7#\���}�j����zV6��n��y7�|��ʽIί���j��I��3b��U��z�:I�&�jO,!S�p�Q���n��ξ}h�=�>:3�,]�,IRYRA��<�usч�wC6�
#�
����
�W�����vi�����I#�Y��w�_�g����G�U�.�ޘF3{Z�^����Hߨ' Sw'm���Ч:�z9v0��>��ѥ�$��
=K�X7B[G��g�+6팷�����fw����L[>��2?��l9�B�^�����_?�i���������O������4M���'h���ץ���ژ�����8�������o?����E.�sџ��\��?��u�qj�����yY���=���_�����ϫ�W?�~^���y�����ϫ�W?�~^���y����ݫ�g���#��!����2Ō"��XrBvL�R��������z7�a�M{�C'9;?qg����y���V@�$t��<Ӿ��W�����Ϣ��j�Vz�>	i��y�鸖Ք���_1?��'k"���xc�۫�c.���qC��"��lj\��foN��>�ܯ���g��?_����^:�"�p�+k��=^c|�]�}�(�-��/[[(�gԢE��|��MȀ>WϿ���ԓ��Z��{�T�U���_"o�@�<j�7*���3��";������+�]f�p'�����7��0Ȭ}Gv�/��>j�Ӹ��N�����h2A5�f(��Ɔ*M��싽��F��^\9{d���ǎ<�S��G��h�ʌ��G{��e��d���9�,t�E�恻D�ŉ�4�B��%H!��hK��/�A�5�ۑ���ص!<�Բ#uO]����tt�h�ڷ��O��/+�h�Z�D"�q�4�� (��X���4v
����.D���i6�:�3{����?�����������@�_S���^���x� �B�m!@�e��xt���:k�����{7g�)A~�ٳ���7	<z��q:�?O��n\�eǎ�+����{(T��ީ/|�x���6t/,W���2�-�.��?����C��,��b��]��---r�hn�����蹑�hw<�5� �NЦ��v�W���!���f�NP��~@Ӝ�@�d�-������4Fkg�Ǐ�w�	ٗ�欣C��y1���#B�_w�h���O-�s�����3���3��P<ǃ���SU�B��h^o�ױ����B�\0�+�x"z�2��˗�hz� �Wn�&!�ko�st�T�ϓ+6���_��иi�6@K4WJ������N�����ʀ��˖����K �6����u���
��˗v��n}�L.����V-��B���4c7$׳�	�S�$Mss���_h~�w9�(X~�J�
�wo_�^:���v5��׉9����~��I炔���0p��#ݣl@2n±\���]�9j�r� `��΁^����v�D^^^�8}m7�pH��(mY���e��������I�srr*�oC���=+z�`^��h>���N��ksw�<�<��0z1���9���o{Fgc��F��^������2wss�s����G�Nt�,���{�N��Jhؕ*��!�����֓�k���SGg�ę$��tws��=�+.*�z�Ҟ���ny��E�wWrfff�i(o�eO��g��~w�ݺkԇQ�P�&�?0��p��.�l����w���Ԏ� 剿����u�S .�=V�W\H@����야]����(�u��^8��f���w�%��C�'
�m܀ҾVt7�n;���f0�����py�n_��+ X��A���ce:���s0 ���O�7Q��-�O?�ض�7�<6,چ��L�]t�h���	qC�nn>C�}u�ޫ%|���Z*���ސ��ׇ���S�Q���>3�AF;(�A1Vc5��(����3�m.[�YG��J���=���0E�|�� ���n^|K�r]{A��Ƌ/��������-,��*�$���YK%�8ǲ��hS t,��R�Z�:x�eb�@N�x�h��1�P`���;2zg������_�j5{��U1#��G	ͼ셯@q�|E[���ŵ�.D��9�'i@Z\BV	ьf�_���.���HÞҥ�4|�G���3@y񽯢o�8���պk�:/r�1��k�c�Pn���4-������ U�\����\'�K���{:b�I2W�I�p����ݹ��
t�Z��"�!���.�:u�!�k��s{�S�\�L�q�7`�GN'��v� �����׼nFiM�%�u$d�Tb��;��{��� U3V\B��AB}�?%�
�;z����Tj0d�K��d�U�l9S�L�X*+��z�4����{*�K�
�!���ج���t�-^<��=4>;��0�R�6>�� `�Zϵ����Зhܕ��\k	L���s�S�bF�QpppG�c��^�����f�+g�K����xUcOU��q͢6�t�����斁�
� ��+GUx������s���+�!I5;{�) ��W���F+>?���)��b�E�����.�Ɏ�G3:j�_��ɪ*�h е��Ȫ�D> y�w#/������z�6�ubIXԣ=3���bdx1ۅ@��Q�x9$iה!�مSuuzR���}�h����P�J8~�� X�!^�K���~�����):LG�|�W�/�IY\8����@�[���忴U�?ީ@�{cq�ͨ��*���)�^�yv��[����0ὠT��wC��@����D�!r��M�Rs;�%"�7�#��:XZ�CszΞ�� ����>2���H롍4m��y�� ���(U^�@����{�W� f�������Rjg�q�ǽ�����&��&�L~����+x�T:!�ڹ���(���O���|�Dc���2ю����:r�Hi��f	9�+h�\��s�`�{ (��� K:�h��h=��]QW��?FFcfgeݦB�w�4��C<�s��o��?(߀�N�נ���u4u}���V۪��VPQ�PG�BZQ	(���� dD�Rdoٴ�+��(�� ��^��B
2�)�Y"���G��O�ͽ��9�s�}�����Ԏ�:s|'�u |0�+/��P�@���b�t
�!a�O֞H��+y���kB��*�H���y��CCC��}
��h�#��NC5'	?t'b�<q��Tx���UM���K����!��5�J�QBg��2b���߉l���4�	��K����d��=i�B�脄�{wQ����U^)�6��:?�~P^�~��KM�18a1l<-c��s��B�֢M��`�O08�4k4%����'{�҃��<�&Ҁ��$�G�E����Bm��0M�byP�}�s���چ��5����/�Y���$�j��A-�c�87>�yP��ƉT0�W�b��ZJv�K�zB8ʽE-�̂�$����j	0}8yqee��<�S^�ްu��ya�k�v�� ��t��,��~9���љ����|�;Z�=7�{%�\��lI:�cVou�K�r�NP�z�:}!�8@lM�P�ߏ~�����TȓC�sK���(~�ܢ���zU�6C(������8ޫH�*�(=���hɿ�h9<\gH���&������S|lG"��_����z�,�׏/�{�f�`�Do�G��3��sIr8gOI�����LR?�C�XqvZZZ���|XY��a&��1�_㿑��c�G|v�0����̷^��! ��b�6P�LD��p{q��p�j���p���]v66��(�7��E�A������JRD]�>j*`��Z|Y���ZA�����:�e� ,[q��l����˗/�f*�H�������]{���D�۷og*��C-��Dݘ�
4��,����շbB�������1~JT!G�4��Ign�~(UsI*\�Z��>��sn���z�~p'��O�)mo��:b�w�Yd9K�A�uY�
������i�/c�/��P�z�s$�r���k�Vj%+yi�qC=A�V� ӕ	�˩��_K�mS<�n����	]L��_���r����Y�w=��s�^Z�'.���(ԣ�l��q$"�Z�ɞ��s]tՋ؊Y��,XK,��~��]������8P�&��g�*\�{�KjU�˚�E>4� ����/ 
��٭?�eu��h���/�����_9A�b>-|�;�zӥ��Q�b�)m���]��k��L�ݺu+��n�}�&�t�9�j楫O�2P�|~��
ग़��{�z��(��fR@���Ʊ6 7���Q�s�����v,�b���ήH��Gm�Rh�gP3�%�Ɨ@ܿ��Xp��^*fE��)�g�b�Og,BQ*c�V�a]V�}�ZT��
௮|���{aQ�H�7
s�Q�=�kOӏ���Nī�B�$2�e$O�"�#�J$�5�ķ.�SKR�J]�IQ�:�+m���ŽHZg��^��sS�ǗJ�>���*�F����Y�? ����)S�:����&E�����Vdu�-��u��`��8��7��DD݉��EB�,
Th`�~JK����#&�k���C�c��IE�Y^�S�n�Yȿ��1���"�B��ɉ�٭���R�{\�PW׮�@m��h�B��2������g<@6t����p>QVշ�k�{Rs�1;!ٲ힕Up�cL�����>�X_�#����m=�O��,�L��y?�qh�D ����x�Ȣ���J4^7���$2�3��y�� ��.Sf�s�*�^Ut��T�|	�$� Ԓ�H��Pd�U��k{{@�Yi6 �%��]q�Q�c���R��ϝ(#e撰������	���������ڴ���1z�r���=U��dH���ێ�>�	s�@���!��-���3+Zِ$�a��bQ���i�ROR50�]]],}���ϻ����ފ[��W%:��M��u�]��f@�~]V��m��#��;��y���J���i���mE�#65}�WQZ���!�F�JD52p�������*}���M�H��h6 f�u�rnh�K��Q�T���Ce��R��/gK� ����Ku���s��}��(�Q�˵�"O�t�O(o�&��;��E�] /;��ٝ�%A]�V(Z���ǇN���é��l$0|,��pL��GD��Jzv�FE]����YV��i5^UUe�N&��-o,^�߮��������?���O?��s��ӻ��o�0������[��m�O�*RRd�I����t��x��1�o'>�sݟ���[��ݚ'����V�8��������g�V�6`��n����-��;o��pa�2P������Vp�|��%T]��'���28��n׮�ݐN�U_��b�Ӹr��v1�o��|�-�k��Я�>T>��tP���� p�}�.*&�&�g�1��{�Z͖��v���e�}Z��-�P�إxz�z��<��;]b^�$'�^����l�AN��a\yx����߃�2;��{���A�Y�/.�2����cc��t�R˨��\�6��]�+�cnn��ś�`8T�l�|]wA(oԧM�6�����Y>���	P�(��#9��rVH.�5�a)+�u_������J�]-��]��Nŉ-�
��{��?�)ͦ����	W ���rC�E�Ы�x8�η���{��c�������m�]�֝���K�}�_\Т��{w�X���]@ለ�X'Eka��JVJ��#n����M݆��ޜ�*_􏀳#\�=�����7��,g���(����%�ٶv!�qOd��H��R5f�ϙ��Ǆu�0�z�)~T_@a�b�/�o����Y-3P,�u0g�΃ؔ�o��U���p�]�*ځ+�^��W�돤%'w�Zu�*��9�ϖ�%�m�=Au�y?ڐt������'W��Y��y��mQ�0�It\`GxǪCԄ5i��K�� ��G^��.�o"�n�Q�?9[UU;RkLYj��/�sK#[DmՂϖ���3s�;Kq�o���E�R��=��^�b[ب`�DTq����ڪjk�<��FUr�!\��#
dܳ�m� ����;���?O�6-4�����Sf�]�����T�s�Vm��^m���߼�߄4�`�B�q���w'���V���9P��!� �`>��M

;�(2x��`�b�'�Q+��>�АPᩖUɕ7��Hg�����F�����dCh�]K$�~H��c#�K�w4ݥF��7����'q�+��ii!����.P��}���;-xi���>}�t�i�x��8u�t��ԙE+Y�Z��EK�A�{��Q�gA����0{J�;���e��j�(h1�&�P��}�^�LcC�.�����	��G�v�F�Z�V;�Z�.�*��ҷ��-��Q�]�ioP���E^�cLvgSq�F��H�@���?��3��Ө���6��c�t���T�G�G��s�[�&�G8�zb	Lܠj�8��ꔀ��#%ȸ�6���º�11y����QN(x��ݼ�,P���2�5�b^�!��QG���\Ȳۉs�8+�y��O��m�7;oN���N>څ�?l��d^lb��\�GΉ�6�fbj:�B0^�t���Zr�)��z��X!Wp�nÕ+V��w�T�p	WUF����_�h�pP�㓑g������H~N]'�xT__�R�Ȼ����c�������Zń�ꪠ�"��8���`͖��k.��.�S�U���4�����75�<XJ0��ڂ��U���M��Q����u�{��$��$��q���*`hv]!@�&��'�}J�I6����!R�=��t��>>}+�=5D��6.�јӧO��u*T?�l��+����G��dge�>����T_�2�,H��ī�;��=��X�8@��@��n7h�M�f�vJTQhɯ�(����(5�)�N�x�g�N���]��8Mfˡ"z�k�|�pa6�G���ݶ5Q۬VZ��7)S#��ͳ��%�!�9���~��r���^�?�ª�F%�,Q��� ����HZ{���]�*�l�`�-��J4�f��y��0�j�L��˓D�hY��/�A��M����2��I�|߆Ϙ�B0�@�@eʡ�*�`32�T�uÖ_��9�#z@V��+��c��f�N*��fk�h�7rE^�yiMY���%{����vd׭����.�����/���5��>��!����27���ťK�"���è��S��ۘ=GP4���������WH��R�{2L����]��՘�gP�́c�ȕ��e�
�Tg�֨��7t63�(��{�����"by�W�7Ko1=L�hBcE8�B���WdT��6��f���Bmbх @	���|<۰�ɢ�`}��d yGҍ�+di�/��x������66A~��BL"�C9Q]�Eݾ���[�k�/Š�0�X�^�'�S5[��W06 �4�h�i�M�/��4�E
�F0W۲X"�j��"0+����q\�Q��"5��N�s�&��s��7�̝��r!��J6�6����:f9�.�T(�+�]�G�Q$�<0�kkk7e�]ܑ)w���I���eCǉ����S�t��%VU��վ[�]�o;��~MM�ac�@h���O�~?�$Q�*3Y��� T��/�If�ަ��Sk��& ?Nx[
UF�kJ1�t[Y�b4�ڏlɴ�����ɗ*��_II�g��k�Y�98.�`T���y�d�.Z�W��]!�y1=��{�<Nx�����eBN7 �|p���9/fϞmp�+d':�o�ْyQg�, d#L_ɼ�-�ȶ�F�_����WZ�b���M��w��6|��!��s�ہJ�Q7g ��Ǆ�����'OYʭ�L�	�Q�<a"�-I ��)[b������}�)zO�$���-�h�T�_�N{n(n*ޅq���@���Ċ�s	���"�;1�Gۚ&�p�Q{ ��:놀��LAM�~8 ���+���mJ��D>�\!_�?2\�Y�,�����:�0ݐ�q��1k�GƒH�����A�~�/���g�Y^����m1	U��T|1��r�d�y1{��h[�Y�P���ʷb���Ԣ&~�%���"��)�v�u%m�B�kC��ac3�S�e�3�g����t5�,'�r�$e����[�x�����4)�S���ԏ��dԈL�kz���HB�9fT�)[�lY}���=ᠼb9���k<u[{^^Z�62�5��ko��Ŭxf;�q�3���1F����TJ� =V�-�<�%M'���׽�=}\�_�H�n��������M9��g,JA��=I�⢒c�9ׯ��"�}N+��k�(s���E�ˆ.u���>����:n�q��ER�gk�+�'�@����8�c����Y�ui�� @������NTTT���VJ-p!��{�B7c��*�OeK�D8�o�fއH�P»>i��U$��N]$2��)�ϴwδ6\�@��/S�9���XY�����n��@!�ϻw?3�2����]뷳	g��%'��t�	�l���e�F�����6��b�����������:v�P���*$���455.p�YAH��YJ܋v�O/�^F��  *�D��W$&o�Ci�>W������G��� g��+�b�g�sR�q�+�;��d?rK8�#̑�6>�s��Դ?  ����)
͒z���
B���
���ԥ��b�$�}�����8����:�rEe����+o�@K��w�<e�1��w��F�H�[K]'���iklū�A�w�?�3��J�4�n��8�ɖ����V��mx�`�/uo�뱿<n`f{{{y����S��366�$�,c>%d����<�y�o:�I��̺N�e�چEdV���|u1K�{�33(�5\c^�%���S�\�[�;�nζ݆���U��b�^�� e*���V|vw����l1g}���E���v�eD�/(�f<�t����,��(�����g�����4�HkM(=�>Ė�^`���MU�dE)M�M�d'�)�Dlʮs�Ri?�*�o�<e��O��xrMnG��n���A���ӡ��ָ�M*`]w����u<o,�?e2#(H�ڿ��G�w"v%U>���ƶ�:O��5��΃�$Pt�1���q���$<lg2=ȆnRe������G+�C�
�%�d�B������6�`w��6+�$�5@�,!%�	��|�����dTw����<�L�P�������K���ҒK� �>�P%C�P�N���x���
K��7� 99��M�T�"�@�d�㤚�������,�ʎD�.u�UP��pߒ�zѬ2�ۙ��^�oN�3�r 磷nݚ��t�.��ؘ=vGTq|,d�<�_u�;cd[?�� YJ���7N����з�o�N��dk�ק��8l(9�S�Ʉb���n�0v%''����X�W��ُSy �Ѿ�ϋTZ��܇���q���6��u�,-����D��A�tU�o~�K���1a(\L:���*��n��Q��Aʫ:�3�����ġ���M��=�_+��B
�C6��X��V��J}��X�D�1����m�.��hZ&B�T��O����STY�d���G(o�� Ld}@{��n/�g��Qv����[˄]x'�{=�������Z��å��/����^�UdJҸ�����J���M�LQ����؍��ח������ �l(/�q|=�F0J���Nu�޽��j�$ֳLj%D�M��Q���c]{��h|/�'���Y�`!�����)�<����.��+1�ʰ�,�sf�@@a���g+r�Y��p����;�2�0����ƊɨĆ���	h`����D7r����B]}V5F��܂���x��̻p3j3����=
���Ҋ�)��S�>_���x�� ������7S�.]:@rA�*��^����ƴ���Tuuu�Ν;s����)Uk��l�A����0̀(5}h84���^��bɻj�d��u���DEiʧF��"��#�u�B�p0����,��p�c)p9��N~�zuvH��U^�iܭ�_��2(��<y�V��*u��{s.[�N�k����۷�$>/Po��m��
nE��G
��ћ�R5<�!��yͿN��1߼�;�sY��z$�o{F9X�up��J��^P����[,q�9�Q/}C��F$��U�.ģ"(�V�)oޣ����: ��ǅ�$��Bܷ煬���Z
3��U4�®\��x�&�]�jYG$|}��R�d<� CO�z�+�KP�BTyUT1͌�*��}�63�N�t�[(耱��s^I'5�=Æ��E���;�G�U!r���}�Cy| 	�Rj뷷Aq��o+jKp7�n����#G�MO��W�rr���yw>��g7��!G]��.hJkŶ_��e"NTu�KV302v��K7�8L`�M�r#���}�U�����Dj��[���p}��n�%[���Ե����tf�嘨� �u�T�d��T�
:���Kz�ަ�%)@=IH�e֥��m�+$����C��� fF&�\U��]���D��������^�wQ8MNWҏ
�����
�#�j����US�a�5����5�+���7�"Bh��>,!�@Ԥ �x�=��F����Y-|l�I����l�|^y�eQI"-�п_�Zm굛찗z,�A}}���ׯ�y!�ø�/�)yi��"�Z��ϰOJN�������R�,Wp�nWM�B+�'�`�߻E�i�/_�����7S�}���������?���L䋠l.��xN�P���&L�*�i�kթ�jX>�� ��?��|����q�0sQ���)��="[�[&?v12�]>{���6e㮹�ڰ�-ܰ,N����]��5���{{��΁��(�3�ȑN!{�����n�oaT!����Rp�l��ۦ��wf5�S!�NK�-��Z�|����m�ի��ғ���k��Ny��p������h��
^��l��Ч��8����*O�����-����:o<�L������W����v9ٔ��qz]�[��k?�	��+���P�� an(F�|�M��ꗓ����@L��Bסg5�Џ�Q����U��q��CNQgΘ6AY�h�Jw}no�f�|��#P����h�Mr��9���---�X-5|�K�����,0�Q�IgC&�}CI:��^O�����������x`�*��w,����kQ���+����o���;R��tr�=�$0}�
8�?��4���"�PKWB�{�T��$���� ���t�Jcb�V�C7����Z��ͨ�ZNkO8�	�ޘb�_�)ڽ�Ly�Q
vQ{��բ�&���C�4�[��ǅߣ��zq]����(8�Tqϕo�0Νp�t��������7�%Ӭ�|��:���IϦ����z�yP��yGv]�ɻQ��V�,�5������z���~���_�����}��m��H�%����:C8��z/_8\��t
(l<��)͡pR�RB�Ƽb�k^���6a;�g"�1�SL�]���X��L{��~�e%L6�T�o�E!_�G�I6���@�.P!oF��%<���i�7�CX�A���e����=T����
�j1�Ğ��W���������_p��Ř�;44T>�ب$�.�z�C���N����N�t���%ʽ��XQ��F�/ch���F���bz�U��yp���#����?����m�Z�Z^#V8߽Y]Scx��a[(^�ٓ��u���M*�tom+++5�F��S�5��o�S�^A�bh4�[��}�a����I߯k�>������Ǐ�ƻ�&d[��m9������%�	����d7�&'�Ȝ��E5O\�K�?c�w�xDl�'����o��k��%����.��9];>=��z�jӓ�x;|<���>n��Q���w�6;�KᗟL_�D���������Տ?���b����MI�V��}��g�4prCo���~zqq\y�]�>^�q�~���P&u��yς��֮'W��Hk=�S�c��Q�hr"/-ʂߠ�v��`(�5=%5:�{o���?d�ip����+:��а]�
=��]M9۹�d�(�� ^6��׮]�~:��o;���1&�b^!��W�A�Z6��kM2\�G�5[ʄ�{�V���5u�c�i�'�ne5��'^�� ��"�8Ա\p	uwC��V���Nߑo�=��b�X������	�B�&������q{ł��:j���*�3U-���7�ݖҗ�lM�[�r��8jkR����$.y����)�-�5 ��E͠.>07��dw5O|��%�Kq^!cP�<ǒ@����h�J��������*b���\�꾑�;HS���K��0��K6F��Bq� ��{��������P5>�r�A�]U2���?bl�.�b������%�J2H��=8&�Fo�����#��o~q����PwZ$�����v�q�B��o��+2��{,�IULy'˵a��)-w?!ݗ�&(��b]g�r�h���COf7��u�B9whSr�K��&
�āG�|��s8���'$�W�M���6�� ~^1�Q<f]i�w�P\x=V���#Vb�W��wdKf-���vttXI4��젶���U?4�<�p���B�Ԡ5�2UHiQX,��U^;eHw?)
)I���ZDf�]�6]�L�3=amL"X��n��Sb�L�W(�f6ct�R[V?	��	�:ګъl*J�toNx�F���]��鳐�b~���"�C���1:��הK��-^Ê��9�lb�.`63 ޙh�fwZ>����Q��2����|�&r ���fw]z���PC7��e��%�*�aR�����K0��PR�l������c��S�4��+$t�i��{�����ii�XܻE���\�;��V:��w��8ө&-�e3{Ɖ>�E���&𡜥���P�JĽO�=�q�˵�'U&G9���lw���óٮX۫���ϗ��
F��1�!�h˃H�Ȓ��\ID\	��/c�V�^�L�6[.є	V�!>anT[`����
[�*�sTvi��^د8��Q��q�#��g�T�=<���ᙟ�J��i�s�=��.fff���`B�Q��h�	��-̞��l�᫾�Ř�Ը̀	O!Z.QѢbg��Rg�,N�K��eq	��ϱ��U��~������v.��=���B��#�"E�̳����z�~'��$�1���K��JDi��W_�Ut��!KXխ���s���N_U��t�ҹ�ր�Y6��w�
.���mO��ɸ�!��kI�R�M{��P#�G
�H?�	��~�#a�&�W[�,lk�]3�Z��8�Dcj���BDQ�� MA��g�G�!��r��!u.ٝN1�ɥ�EQ�H�ݻ�������e5ڣ����g�N.�5�(����\�5���Ib34Jڵ���Sؕ�5}�P���م�d����Q'/h�s.+/O�ыS}!��R��j�����Mv;���m>q苢�y�a�ڏR�;����*�P��Z�w@*H�e��`�u���� ��Ѱ�7R���z�I��t��o$�.��r��C����v����Q��l��x���cǎ%��IJ`��1�CqS�u|��9uLv43?�w���x|��wX��D8���E���ܾm۶�h� 2�4D��S"��)�"�K����6�����x>)z�U��ʽt�1k�DԞ��ڳ�7}��sa䅸)ϯ�1�AP@=�
���Ak^=����Zo{*��G�leU�t8OQ�p����:��	���zf��N\�:��;���������ٓ^�A����r0T�n��T��C�^�0��Spir���%{5[\[�7<� o0�
ތ�5���R�־K��e��k��f����ɩ����+L�+Z����|����aެXc_���Ǵ�v�{�(�?���&'���kW���V�_��[���*���)��H�G�J�=/���	J���F�9,�1�[�nL��k�-�my!���ՖS;��	5~J�<ByP��L(̦8S�#�0���-����b��5����K�M�������Rw��5��Nÿŉ";���8h�3��*�+��fW꤀r��IPU\�r�{R��Rp-���ݚ�+��6*��<�%��7}�D*��G����X�0�KV�Ă ;�hCV܁�+��!,p�UU>�%op�^}u�� E�@z7a�Ժ��{\y$���>�ە����C�#G�*SRR"�Ʌ����n!�篢?���KC�_�]��ܨd�sNԻ��$:����+{�t%�{ʢN�3u�Ļ|���*N��\y�֘������K�y�fS;����`�~�w��З�x�ak���l	)|�=(�}x��yL�M��Y�I5
=���{孧�sv�ᆊQ� �����(>�����(�_�jD�!���52��S�u|/=�U��v�}�Z;������\�:ȥcg�V��� �Δ�%_�\������� �i���Ww�ګ3�5��ț��	Р2�����{����:YT�(�_���J	o"2��íڑ]l)
W�za{� :�PHΠ���s�5/���5���0���đ˩�cf�:��&�٭��U,*G*> �r}���P��CV̠QP0o����T�r'7��2�N!c�N(��._^�P�B�{���T�����L+/cם�Y�L��������Q�;G���F�9�"���L}����u��?M��^�	p�����M���G�G�$xpE�4ژ��0p��o���M����,wq��
�����ׯ_�K/~����\��
�U�&��&�cؒ�5���G���YM*u�}�U_*��K�����,D�#����4�ݱT�>��e�O�am�3�E�6ox襔;a�os"7�;�7�%�;���i���?`K�l(�c����z�t-�!��a���	ԌQ��m}�@�����A[j���E�l�����a������d���w4��h�_-�F/��]0[RC�U>E�{�߉���wL	/j��rK�޳�|r�Co���"�=o{�j�ʙ.��+��(\��݁6��.��%�R5G�($��;4��=_nrr#�f1���c��ΧJ:]L��cTMA^�p�p���9K�=.����S��4�J�l�]�v����+��wSݸ����Z��r_�9��<\���ˬ:EvH،57/Ѻ ۬�~��	�"%�-]�rd;Ⳕ^t�m8�4��9���G�}ZK���N��ZY�=%ō�9l�g�����>��J��S�4E���Sܔ1��|l��=>����0�*>?`иL�FH���t����c��*Z����P�Ol�̥���K��չ����n��V\y�&������̣��]oo����K�0kr��?<e>��YxM���dx+�CX�$�`TԻ��Jrp=�� U���n�P�X�x�l�0��\`b��U�D�#���ό�A.�ߌe0\X�Zy1ќ)��0��Q$L���w�$����OY��y�T��+ߎ��L.�hgʹ1_ߵ�[O�U	{��I��2y�}¢��v5["W���
��"���_��aDp彚-K�x�m�S�x���J%ͮ@�����%�r�u�6�^�K�u���!w���dC�P~U�����Iz�H��<f�qa�l3���\�Rzѹ���}�����-5[V���g�I�<Z�����؄���y��L��B�HW9�F��ֈ�6�*+f�;eq��oUEE�L⚟ӳm���z9Ӄ��D�����5�~z��5΍�u��)U[�R��
�C|L/����{<���PK>ڈ��m����֣n�Ѻ �\\k�������X=���CU߷#����@�@F��#�4Bx�az9p0���,_����������)�E�e�R��!C�!t��Ԡb��v�7�i�@F��"22�JN��v��/
�_(�����w9ò�/����ɬ������Ya�W�i��K�Z<��5a.SJGf�w^%�3a�;v	����`P�.cK��q_���%�8�ig�+�u�R�+�(26Y�%N��O�c�>��lieG����$F%K�v�԰߹s'�(8Z�NLW��)�g�� ���Y� �W~u��*��w{ ���PP����Ӈ����3>���r�l�UX���f����/����|M��Wrr�v�x��w'-����q���?ƒ���b��C�?7�t�W�B?��Ç��>���X	�3��wym�{�ҟG�܋��r.P� 2��〢'��'zBQ^�[Cq��,V�����^,�3�cH��Y�~_�z	���#�H!��&�H�Z�|l3:}�����U��Qq�>�+R�%0��V�x�O�(�~��*i@,���zy��"���%�X8�������h��\ya�]`�y%�k�lP�-�͑��:���i1��\g@�|C[�ʣNߦ�2eǄ�Dz�F�]vv�7�K/�p������a�"lQ�,�c�l�_�}�ї߀ĉ���Q(���j��]��xs�7?�5�
��]8��)}-�кn��Z���q��T�H� ��vL5���T��ܣ%s�OԽ�،W�O�˹\�ސ\�~O����9���y���o��F�p�pG�<�'��~l�y�EQ|S,<�}LOV��>|�+�E�F|�/�އs}69 ��C(܍��.
�����O �he5��nJ�̵	C�D)ަ�I�/`f�t?��w�M3q���Fe�kh0G�'�/�{�:�xM�W�o�K���H���,ta�?>H��&�|beU���8�u��g�S�
�s2������*�	T�G�-��D�)�X�x���|�Vԃ��+J������I���$X��;�
P�W+M��~�0ѹ��%�i<��u�]��e�'v͜�ξ����6���hk���~ژ=�`є�W�4t�@����������Ŭq7���C+V� E����q]�S�vO��W��IT���(���`�M���a¿���1���Ht��>R\�B�&�jP%R�b#^=��m��)Ӷ��qG�裱����Y��j�j��%�;K��k.��
���+�%d�d2��U-�@���	��f��,���j�����c��}Fs�q���>3���1����9�1M�V�+[Ҵ����*��
��Ԡ��7�^�!p�XX�&ܣ��Ɇ�{HE�}�kX5~Ёf�R&�sX��Q$��U�UP�� ]N��1��''����r���]��j��jN��
�����\v
�~�����n�
��(}��p#�P9rs��zcQ�>�JgL����E� ^����ü����� ����}�~D����v�l�|�Ԯ�v�'���N�;�Bx��ǫ2�����4��ܦ��T��&��dac9�}m�K�{�F+�`w�g�"L��w-z9DD��� ��ki��þ`�#m0I`�I��|�q���*G��LKk� �;=�fl��ڞ�Y��E�/h?�q��$9��S��K����hqW�v���l�/�|2�ri��6~�$����5��IK�*K�e\�������璓#�J�ٜ��̘r�#N������G�?�m��w�C̙���8�-����#!�:�ad܃���ӧ���;�Q�K�洽mʿGl�.��y�-�!8e�Q�� �p�fZ�O��}����0�z�^��P�Dq�
���/4wM>���0*hK�������.�����.mN�� ��hm���ҟ��k�K�GA�?(��l<�-�pʴLRE�r���MÄP?i*&�q���E,�MҞ�������5�9HP��P<G�Æ�(D�Sl�wSff�1,N�VO�w='g���� ^^|'�V֞x��y�C���9�VU5y}��';�X���a�J��C7<#/��P]�����H_�������f3Vs`���bʡ�h��ct�����:�+O①������dD濫L���0����|���ޭ�?����h��}| 3^�,2�M�:0f��-͕JHuK�A��k�z~ۇ��=�l��_�x�lԘ؃
;�>q���$$+t�YZY5�1ˏN `�����!�愨"$���[-F�VNڪB��S6�2�g��Jh.~��E�lk����{���i�ţoG�n&��~���n�;*l�\�9�M�bH�ю���U�����B�~z����=�NE�ǰ�/���jO�����?#NY�.]��ܘm�Հ�y��!�NX��8��$�1h~o��m��	߮�;�����u���X�����/�?^�v��L���e�Vf�H-]V��.���3su�Vtj�����2���{~������?~{�����_|�KzV��V�>s�m�ee>	^v���c��n.��ߏ��T=�v�knk�P�(��� ~��^��fS��Uq立�w|��ӑ]���ں���͏�]>খD䄗mC|�28��a��CZ�������/�������U�Y�Ϫ,�֞(��fVk;�|j�mc!і����^)(�i*�9����t=�Ws��!Gio��LII�(��d_�������rp��Gh�ϙ>�~�d4���zUdQ�����נ���]wtOjߟ�������0�TƥDGK��e�e0(/U�v�c�F\IttMϴc2�@]əE�.uq���F{�V���[g0���k9�@�M���{B�쬛~��L�řk]������F7�ÄB5�#�i�E���g�J�n?6S]�Mx�
C�E�Л���י=���f�X�D&*Й���Ꚛ��U�o�b��0yu�ʲ�\��UTT�f��t�f�����<{����1�m�D����0p���=N����@j��n �m����7�Um],�����w�.u�Q+�tX6o9nta"�d��rI�Z4�����\���,����2"}|���2=B������q���awV�=>�	n����r���˓��O@�-��gV*�:�������c%�o߾O�@W��MN1/��R݄�M�ԉ���������1����ze �g�����N���R ����0�"���<b:���������w_������cD�g�����}���$h��ߙv�/%>ř�%�%0h͂�a9F[f��Q+���5(�rZZZ��X�ƒP����C�
ʥ���wy�:��/e�,3��Fe���~��̣å��C7�S��V�Z~�d��vZ[x��(uM"Z�j������ $��9E�8W��qa�8�j�K]�݈}����������#��,�R�i��Fmt�HϨ7r;*@��4��-�k�]�,�Μ�7*�s�2u�S���r�ϛ����|��k/bE���s{U��+@���02$۶o�o�0{����L�2�=�ퟔg���X�u;��1��s����H�AT@a#@%���n���}��w��\V�M7��tC��2qɖa��ŉ����wE�2VH��i�'���ݘ��Բ��V�dե�,j��ӎ
��eb��ᗕZq�z�O 
L��0/�n�����'խ�hZ}�D��5��Q(�dPn�|i�TR�Ǌ؇����/���з�?��{�`�S�� :wxl�֓����87�D��T�_"����f�};�x�\�F)�hխcN�QeZ�ʼ��� U+����4�8T.C����;`��&������:t�`���!��[i����8O�R	>L�4���ΝC?���
�q�$��Nh $q2��tl<�ZDC�%��^��Npsr��HVK0n�1_W�_�	��4B��p�f��U�3]�=~��핽w"lg3��=��t�G4�J�`�?�c#��#�Ba7�Aҋ��u����n�r/�����`�6n�Xr	�
����g�W!#�.�.S��:s�<ح� s�3\v�d4{pՔϣ�NNN5��6��M�͏�Q�'������X��p�����S���+vM����3�%��(�^�m"'���*uC[~��y�9����E�dj�q�4�ٍ���r֜�0+�N.�h��兗��g��R2�����x�B�����W�O�N@���6��
Nt�����95��c��-��JF���9ȃ�K���P�y���:�>ʑ&z[P皟��߹��.ch5��R��酯l�v@��˟\g�<!t� o�`�G�.�%oRg�u�ԾlVK#Dw�W�ð������@�˺���K���#����s�D���U31SLe<4�TExE�u�ԫ��Zt�<<z�V���q$�<�R9bQ��@�@���Fm��BZ��n@iAJ��jp�Wto���6���VE�I�,�؈�cޓX�OW=D�����+���$x)���fy�y�b�a�
�;���IU�Cϣ�d�Ӻ8QPȍ1=�y�pa������zGN
�3�a���}~�L�ޘ�8�6)�u�N����R�\�v�֟y'P�e)��!ޟp &c]����� ���Zv@|���z�J����V��,Ѱ�z;([��:�4�7�~�ŉ���#@<v���	D�ƣ����|��Am��cr�A&~�ώg���yV���ͤ�P��d�P�oV(�Qv�7~�	p`�j����~�nH�����#>y�|�	��F�K]�;ɭ���"U&��h+�(������N�&��O�c.x&3��������7�t�BV�Z^���K�*X��'_)M���5��S����\ �b��+�l��&����E��[2�	�D����	��{č����������F|��0�?R9��~�`g���2�����x��) ��2P�h��$���1r�PX�f����?__�u��`��>�Њ�Oޛ�K���ֶ���Yih�9�}�o�хGG4[�P��2��~�/'�\|����Ka�R�������]��UUU��~���3�X�8;�1�^�(f�q���K����ւ��fc�}����t�A%�����p>����i�S�Oz�MR-~�٘ġ;B�h�������P��K4竇n��ރ9[�3>�t�X���vk���. ���� /}��
PoB�D�0�9���^=�e�`��9X�,�;6��mx��v�����%3׼�Z^��� �ܢ�u?|�|?�i��RSS�/�i��Q'e\ڿk�����)�{4!#�]�i_���.��:���a���{?���=�"�#KN� ,K�0�^�'w���P��;�-�[���)�C8����yv����vu�����n9��-�v6O	� 7�M�*O:��*7f�Ƃ��#�z�G��?㧏�p+'$����L�_�9n4 �h<�?��xAg�0�<ί�0g
�����5�r]V�� ī����� b'�L�
u�>��B���G��Ї\t�z�|����y,���UgMf#Ĭ�-�𽑁��t�릂�J�'������YL{��0|��s���9���'+��v�CQ}�Y����|�rPr��\�7��R�k@%Ow`��^h�� ���]��{�M�$�"��&_���'W>T]]���$
#5J������.u�$�vD�|d��
�qƑ�揭'�}gY��2�ָ��Y�;(�|��0��ɬ�*#ѱ�I�b��ə�����K��u��o�M��u{�ۨ+�@��-I@�ː0vFQQH��-zO���Z��0��Щ{S�)4�_��Ϳ�<���i�/����PK   ���X����<  �  /   images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.png�YeP^�'X��YX�C�$�������;X�ӥCJ�E�nI%�P����o��wg�93�g���͍��Q#1����H4ԕ���v����NI%��g=�M����z��~'C�Nzcw{��K,~'7o[��K~w/���2���4�
	��bz.k��wx;xq������[�����H�S�^��jz,��D���K��
9��+O��,T�"K��B��l�&�|?�u���YTT��1�2������3�a�!t��ư:��4��ޖ�[�\È��9�s(&�k��������]7]�ǃ�A�})$�%y�4�?u^d+�O�����k�Q�b��쫛�'�k0��b?�����ckJ�,�}��+�Kd5��Ҁ`͜�FJ h֊�d�OU�Yz$��D.��Ff�I�g+��\
1��{F�rV�7b��R����	��b~���&()�Rz�(����,��0��K�JQLD�9�R*H2��D��x�щR��㷸6ΞF>��U��a�q�Z�$Y~2�By�'6��ZQ2��`k$�bI�������p{]����1 v��X��f��2��7m�AKQt���L�;�{�Ե��h����czBSiH�D��!Ź��[La�����;˅x~\�%�f��T�ϖt��ߞ��ǩ��o���m��2l�f�:������>bE3^
�{�V��(a�r��^�.�L��)C�5{ǌ��!�?�W���ѝ>cl�4'�p���؊�g3+��G+`t��n����^V�L��4�}�DV����f�Pj ��޲dq�"m��BP^���[7�B7�\����7�:C6�=���\IIvZ�\����]�������
v��vG�,l���=?L
�0R=ƣ�S��8U���
�d� �?��>�[Nƻ�1���sLP@k����<�oD��ZY�U�\Q��q�\h�]� ���jnB�uk�I�ōre���<�ǀՉ(��^��/���3HԞ�b�M�-I��%+o�.���׍"K����hFt����}�a�����iiC�����7}O�6}�`���^st���Ƚ\�aB���TC 5a8Ԉ�,J�s#
������#�H�cS5G�|}�2����6�B9Z�I�&*֖_:��-i`�U=�1L����ӎW�o���p��<D0Va��qC���"X�_�/���7��dB�.���U"ST��u�(�;RQm�<4�E��c]��?Xfa 2��>�זY!����]��\d��d���9!ɐ�*�ѯ��o�9)�b��w�iF?a�
� ?������wY[X�߶:^OL8�-"+k�Fp?�f��M��]���v.Lع�O ����pL��g�,��&�L�릆�Qk#�C�]�g���*�_������N�F�G���i!U.�JlT��r��MDX	��J�L��p%����ƻa��k�>_� @��$��i�G-���_e|!o�Ш.�x�I{�XS�[5V�<0��`�X
�	,��RԝD`��6r"��Ya�[Ǌ&�+�����g��������^k��qBT~GG���Cޫ	�7T.�%=�Q�k�~z���_ǣ�u�*2�z��p(z������L�zkļ�Ŝ�#�����
e.6�$��O����ެ��	ZQ|��"Yz�	Qj�h�S������.�}3�����E�i�-��䲵��0MR;���<]Rd�d>Ɩ�c
�P�w�����ЂD}���{���zΒ��2�R7����;3��������w����9s���1����g���glS�87�*]�y�C�|6�Gg�4Ϊ�i�j?�3��i�9JuxT��f��� w7k)��YLY)�l�#1Y�D��u�-���*��>��!�@C��)�h��#��V"��?��Σ�d�?�r~R�S:��%�{m�F	};��Ě�c�c3z�}7ܽSa}��g5C���f�\Fr5�
�B?���(\v�7�/vI�⧥	3bb�^���������"&��,u���(�~���QD ���PJ�L�^� |䵖>L*� �'��Ԟ�URң�Gїv�Z����C�|2&.���ܮ:ۋ@�UX+�fG��Dn�m;,�oC�ݗ�{��/�p"��I��b��`�Ӯ�[�nXK�7a���!�WIې��j�*����eЦ����V�7��|i�ܴ�����фRO��/ţL��B� M(S���~��GVa>#u�����ӕ:DD��=�r�y� ���zi�D�� �Ò<� �J��it�e��т���+-L�:(�I"bZ8/�{�F`�i����1�j+�+!��qJO�B�ZM��ww/��-5¸��D�Ulv��z�2��!��P��G8��ZT���G��4����x2�#=�k4֍����O���V� ���pбe�ˎb�ǧW\�0s��<���{���Xa���:T�i����_�N5N�(��w�?=fd�w�Ƒ�ֿ]�|8�j�4F\'G߮�xً����a]0j�*�By�����@��1�L�����
?C~r�?���n����j�{�?��5�P�.G(]�8I�i�*2F5{�#��]�����l�X"ȓ�>So�&U��Jg7�^��GMd�`�@hhw�6�;[��1��YZ1)͍y���ǫ�q�l���S��-tMM����Ry�_�hf��Lf2�����4L����I2]�2�c6%�٤լ��s�ha�Iq�y�)%qP������ڿ)x��%�Զ11�x^��Da�t���`���x��H���;��c��20q?hv�4R��|�A��TK��4�"�����[������h|��hyg�߮P �J�ߞ�=,
낊$�\x����k�����W+Ԇ����(]�b@ER�J����������/�X,ү��b�	x���Mp�E��L��q �)TTlٿ�+�RC���a����"�v����.��66��϶b#���X��yNı��U�j4���ԥ�9���{I/S��Ola�A���}��Hԣ��Yg��5��p=8�)w�%�c�B�xyRLu��\5S�I=���BU��wْ�d���>�JC��_[s1�p�ˮ�(�Mkd�*k(x`0y���ϼce��"�JrU�_�6����X<��?"����ۄUD�Y��k� 	|a�A/�zЛ"����&��45p{�wo�7���˗�-�Y�63�n&�\�G)Ekq�#��b��S}i(`�\椨k�o��:/�'xL��.{���ǂ?���(i��p���R�$*�S�e��ͬ<���Е&9����d�*+Z�\���5�6)+��@�O�>���#�a�5(�}��?&���F����t�C4��p��Y�ݽ�0Dwdz۹��)KNؿ�&D����Y.����ʊⱢ���=J/�
��S����U[7���-p�AR��@�r,���t$MS�����XrZO�?(`)�֭R�H�i����]y20�EU"����=�Y�Xܭa�q&i",N�ɵ���j����]���������`YG��3��ڲ��*�ػ�y��~{M��@� ��:j?Ď,�3��7�頤~��1L��"���M��!�|'2�2����ʩT�۞meIR�xH����J�۶�E�Ĥe�Sj|j�݅������ �M�frP������n�U����<�C����]��@3z��Z=8Olֹn(�Z��Z����/i��C� �dݍ�N�>$��4�yp��o�rO^Yۈ�ԻB��Е�ސ�jFɉ��Ö�VYw�K���6����wYg<6���ɹ�d;~d���j�e�a��Ld`y8w�/��W/��Bl(h����ū�&�ATA(}�W܈��MIpT�>���m�uq� �l�^����R(]|��ݮ���i��Z��x�j6�j�L*�~��
�d�ꀯ�H��nq�G_2=_�螄�� ѕ7x.C��nyq$�R� �Uv�=eHF��cE�9)Q���m�M��&^^G���"�W#-5��x}=c��5X:7v$ԥ�>�,~Q4-#n�i۞�l��+X:TV<�ѣ8�xI��ε� ��Hr�3F�S��5���B������uQU6��Q����9"H�Zzk���l] ����4�K*n$��fg]:�%��ɹ�]X�Y�e�l^7}������hU�f�{�=�
M�r��^k,�^��5yn징k�Y������^���9�v�x7�~T�g����ʫ��n���p_�ʐyZ�� =��P{uz�6L�)�E8�����+� �^�h������j�UOs�R��t	�Y�\�J
����a� Gˊy��Q�xqq`I�~ 4&´���#�k>�M#6�Wb"w�����ڟ�VP�f+��h�1ֆ��������'Wy�6P�ei��Y0���w��L��@��ѱ0O��(z�p@U���`
��G~�Ӧ����pI�R
�f��F-��T�<�a:2%�^����4��
j�BP<�����=�&�W�������tn���y���1Ƌ�QF��_��.�8�s*_�՛�r��w�JG��Պ|g���+9ho�����9�ۙ��V@�fz��ȯ��u�}����Xq/k-���:q6M�H�欨�0R�T��q	�M�xf"���t��
.�B������/�*Q3����cẋ�dN���K�ǽS�bkFT^���"˼�����!kY]sQ�O����?s�r�U�G�a��2�^��ߥٹ���D�����f�p�ƌ7z^��$s$U���s�sfW�Y�+�X٫����?�SxN�;�� �%�L���yrny�e����`YNZ"�Ҁ�>�TEp��,��f�1N���DR�sD_~b�]�Q�|�`�6�+��bF���+kk���o�FV.��%9��7��}�G��n9q��@4.�}i�ܾ����z+l6E}��`_�,���V�q�o�up�e�� `�U<A��!?�P��tUe��u3?�q�"ʭJ®���@�TP2�s-p���,�O�VV�}�k�d��I;r�u���eOCơ���]�1��3rZ�l����q^$��Ǖ�r��D9�׭<EH��c�����'Mm�5^w��2�����}P#=l�1��I}�����꧵S����-M�d��͡�2�� øL:!�H!P���@ټ��ru}���:��S�s?��t�X��둧�bC=D|�5U��~��b����IH/��Ϋ>ݷ����Kc �J� �<�j⾔"�f~̑Iuҗ����C���"թL�C�_�LZ@�����זxf���(�В.�y;g&Д����P�2��H;�N��wQ].���t����J��XE܇���SRT�Z�j���ˮ�M!o!� cLS
U"~u�P�N�˻q��%o�~�"�a�����[�:�o��=�i=u��2�lHH'*�����͙��ï�w��H�3��c'Q7݉��������m��6���K��G{aK�(d��R�w�=��?�_�G���X��� ��Ǐ�&�' �5)����ߠ�œ�	�Q1u-\�5���x������������F���/hʤö��~ʉY��k��D�~� ��,F#N���Eĵ�����|X�=ԁ��'%ѝA�A��m�Ч��[�l^� ⷱ�����/��/K[��_I(��/���U)�Q���2w�y��mr�z�Jc��i�W�o����o��Z��fO�oi�6* ̳3Z�|��Ɩ��I�/���������4gt�S���~�aɒxn�6A����V��5S�5�=ZeC�1�W�S��ly�(���Z��K�r�N�C��2$��"}�g�F���N�u�hI��UZT�Ǘ���QJdgl�3���Z�l̐���&��U��?x��|���@��L+�U[�	P�i�U���Y�ݧKG��̡c��K���"��
�q�m'�T+���}����{��TY�3���/�z�Ș�>�E�"i.�z��w�����cW�1�o���ݴ�r�9�6�.?8���Me��*���?{A�E��c�bL
n��y��w�Jp���Խ�O��̷���X�����������#�T�5FP��b�����N�gO=3��+.�5��;�>��rɿ����=���'����H@��}N��U��3vտ�,�M�oTK�cX��VU�i����X�?0z@U!S+X���Зm���i k���O�Əzy6�x�",�XJWuU(�/S�����fM��F�������܌6�m�/(�n�Ѽ�ĉׂ�	�1��cf4D�#�6�lͫ���L���l�|E�
\R|�=珿_�Æ?1X�V(V�%7n�zح�*F�6@-�'�o��������*�����R�bϸ�j�Y/!ojݵgl�[�*E�
 ��Х0/��A���'Kd�+���^�,�_��0v����w�_�˝���~!�`�u~餍�s��x[�v{�Y�۟�8� �z�����MY�k��#Z�Wr�������N�vS�4���drI������Wh�,��ԋ�X�E�U3�8@������%2+�j���%������n��[)���+�Kǁ��3q �?��^֟u��N�S�N�Y�Ð�\�"��RQ׋�['��#�1��^�r���(�z�I�]i���4;2��ʙB��1p��[�Qno
 Q�+��u7Q|}g��lG� l�=������Ce?��޳@"_�L��X�l~~���Y5����?h�D���bD���U�a	��3��-��ۥld�gH��r�ޤč}�F���.�Q��E�i+$?��'r>��i�}�_׹b��Y�V�v�s����_�nk�J"#�N{h�{7}u!�����n��R3�s=|����/��s�˩@^7M����=��=x�級̢��a�{�.R'ٝ[ً!�!�L1�(�z��$z�����]����*�&��ŉ�T���1��N�3n���c����$�@��;�-��=�q�x�#�:^1�� �T�_�%`o}��?�����&2�}��:�5=����:4?�&���Z�&����:S�,2-d ��퓼Ɋ��р�JU���[!���{�'�gM��2��Z�}Kr���9��]�P�9��Ac���P�S��#�u�n^��sN*���à^���7�	ߕ�p>�l}�ӂ���Z'R�y��E�e�/'b�%@��3��Z���
��.����V�A�H�K-O����Õ�n]�it����6 ʆ�7Bo�'� �5H�vl�K�F��=Ԍn �F�c�i���̎~\���3�/"Z-���8��3p�z�}(�L�"|tYz~����?Kj`g�ע�		�
�x{��;s�$u9�+�Ĝ��|���}�]�
���׵X14�9�KO�E��=��?w���p�9�{i�ks���oip���Ww\�\��{�"XA=-c�b>����ǈi�����f�ǜ0:���sh�;����QC|+�U ���B��	��O���H\a'�N9%�[��c`n�c�N�rn�����۞��:�f�h�n�[vZ�_�)r�ۚ/1����S�í*	���W���hp͕�?�z­�����8ڸlx��d�i�:��/���zE���PK   ���X���7z  �  /   images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pnge�uP����iv	Y:X%D$���e���T�[@���f)Ii�R)ARZ:�����>����s�g�{��3��+Z]U���PA���֨=�A��U83�t�7�@C���o�����B=������r����p�A����|���ae�j���n�u(J��FK� ����>�&j� ��"�>ݽ���vЦ;������p%̑���a�Է���Z��R�P�Źy����S�3�g��'iĞ�j�8�Z�%�Ww�G~ڝ�ջ��\1��pY�ӭ�Ǜ����L�>�����֣�I�'99y���������_�_�"�m�g[#�w�G��,���o\��%�*��&����o�i�7L/�f��;��`�Ҳ���>r�92��{�H$�s�٣���<??����QИ���?��)�G��5���>����7��II8 �_��ia���0-��;���>������r9�ﵗ� v��eE�|R���k?�-?=�l�o<�Cj�A��Ӳ	~�e�t��w�´������K(�
�\���.?a�D	�:����'@7ݬ���� ߽�����}aG��o�d5�J0�#�I�� GD��i��p!�X�x�l��G��@j>lF{�����O���`�'1�		��`kQ��k�n�+�߲֕VR���@H&����ѩ�_Ĵ��� w����[Tx���F�s*�m�E����N�*�]cX|�<���"�P\��҂G����ؕO�i
�=I�Ҩ�8��#J�h�6:N/-��ڇ�-N� 	o��Y� �����O�E��{�
�/���L�kp@�wy	d�Dލ�V�����M�O�ru�Ñ���7�M*�P&�i�$g�P����ơMؒ�?J�x�]�'6J-M��%	т���bq��6K*e'竏*��ӰM�%����[��w2��S��፮E�@y7�J`:��;��Є�>�L�Jq��1x��J�
�O��[y�mN�P���].�H�ԋ���k7�ܢF�G�u��`�e�Q����<$��v��a]A>4�6t��J�`���&���7k���sJ�=%Nm��	�烥��+g����\e�tC}ە�nsߗ�բxy9�WW+�IfQ����ȳ�ID����)t-�=	�(Ke�z��+O/L8��0LDQ6�P6�(�T8��C`�)��ڔ|Ox���˧!Y��u��`���8���[�}��f�/�\��S���8�\�����^���B���İ���B7[�2k�L�t/Ũg_1��ǃ����p�ҌI[�A\����&I��ϸ�G�������4�ihI�	CX8`�<!�����3���xnՎ}m�}��Hui�!�6��ޟ�^��D)��_�]��� ɴJ�+Ţ�ۅiiC��
_�$���b���BF�GHā3�%���㘂>�{:���,?�f=�i���$Ga��m�Lx B��Ha���8���݇�ǣ�4_�(U�&���fY-2F�'"�A�^Ui鱋�lB�!具�"ZX)��חI���r�6�9y�@�nj��Y�L��KvQ���� 0c�'�[����ǘ��1�ߔXb� �ٙ'�x�˓�q�
�b�������Hά0�A�8�.���nc,��|qrZ�ޖ�����+Gٽ$]�6&]��L�u/,d7P�����O��4��rtQ(�U7���[PX���Қ����t�����cp3�
͵\Q���l�;�n"�;����p��y��!�;����Zt�f��>jg��ƾ=��O/�^���TY�� `#o���t�L���QD�����-��}��B�M��es���wh�Ϻʩh3im_�6Yb���lc�y����]�0�Cw���0"�M�2n;��85{���Mݱ7��uҵ`|%A�z!}���
i�VT"�X��e>'�}�	ռӲ�H±���l���b}�?W��qɄ�������E�W�M |��L"�!�2WW������tcPh���wDpo�F�P6nh�����[���a}��I#{^��X�p��ŌN[��j��*Q�==�%<2���;,r��$���7��_�k��ƚР��
ݪ�Fs�S�}[�|W�eG��������~�n�"Do6�K��u%����a�E8��F�D|��2��C���5�^��q������<O���ƹA��s��(��4��(gp���9U�0���޳���TTFHQZj���z�`�k����	Y^�-e%�ˠ���܀Û�����Dq{y#�r��G9�2I��"�Ke@;WҪB�y���hF�z��TL7�&�ȨD5�2K�> �Z
8�OfQyw�'�!�2�q��-o=lq�E�O+�˭�X��'n{�^YOI���v����y_�V��o��)�\q3?Kf���^��T��l��]�Tӯ5�Z˗~q4��#���W�`�����Z�������ed8>%�Y)-�	� ���'�;���$g���)0�Fǔ;`K���l (���y���S��O��߼�>��r�sQ��l6<njڛt�!
��<[mg���s Bude��g����1�\��"�}�&��2?���'K'"��/$b��o�2v��j��{���y�0j��C��3ngZ�;�6�`�ݜ$;��TJ1>�jll���8�6a,|��F�]�ٹ���۟�;��V�Vqנ/���õynG�jo�M�+�ݧ§��~��'��I�4�^O�����H��/Qδ�!����jz3�����͙�b=6$���nE�{��k'v��s���)���`�E���i�g2#�C�=Jj�MO2�����z�֡�?h��F��8��y�&l~�R\-h3U/�q�������������K�h��|�����X�I��r2F�54H'��O#(�Tf��*?�و�����}��"%�����ۯr]�C{����T3����0��6��{�Z�h=��~cdr�go��Įj����g���3���f�z�g�[&�GՉQ[. �WNn�wU�o.�#P����$t���!� {z�ѐ��s��L&�_pgk��d3��[��]p��d�*q'����wUN#(U������~o�0�����g���J8�rC�@g��%֤K}a�( �؍�Vy��%V���(d�ru޻�����q;��]�J�W�a�~�&��L3r�a׫n(*��l"9����t'0�@�fE������t>���Uen7���i�3-�7Hw�Ol��;�����L&L*�qLoFJ��?dǰ����H[5^(����+1$=�\���e�9�L�^�^b.s"vY2�j�|�Z��6y�n�J�E��j�i"�����kd�|��"�a� ���J�����B�F���4d뢦@;�7T�K���a��x�Ǆl��!y
6���	�,QjK�f�3�	~�X�)X����K�[�h掲�4O Ϸ���V]KV2���<�/�pn� ^N���. )��r�׀AᏉ�<�C\Á�}���Z���G��ˀ޺����v�N�"�W�ȅ�؊���ʎp�&{������*p��BZ�!(���������(�[�S�13�i��"P�%$w�Dd2c��[�k�Dώ�ǚ���ux������`�����͇����Q��
�4�T�f�k-���;��)����^��Mc�*���ggҊ�գ�n� SE6N��n~�iP�/�[q���ʮ-v܅y�R�ˮ���뷖�����efx��C�N���ɽM�O�gq.?���ֱ`�ь�ăz��'bSrԍ����to�7#���F�a/�C`�e��V����^ZF
]~p���6q��$r�`��$`�@��N���y��%5���#�P����ڬ^�C�q� 0��)S��2p5=�����d2���g�Wb�>C�&���]�Fހ~�Hl�G�����!~�UU�F4��魕��]��#�rNWN��r�~E�Ԁ���x����ݛ�:SUB�+�*Al:��}���P\����1���C�uRO\�K��X�}����6�be�~�ܶ�_�x��8y�iL�L�\�^�܎B1s�,<o'��=��$<����(�a�8[�B�Qe��c�3��4Y�Ҧ/�u��	T<?�N��F���r��|~��6X5A�H�;��5mЄ�Y�޴�m�A�eU�9���VtU���G��{ؼmX��6���tT��J�m����e�x�4�Mۇ},�n2�H�.E�����ʥ��Ftv?���f�[��H��.Z�;9j�Z�����t��~����e��V�K�*ߎAq�D��,�1TP�Fm��c�
��z-��]����6�eX�������l{�U�=N�u\:�M���]M]�T6�c���(��:<&���!�w<�q�� �F�s
�6� �`��|ѐ�
�����L�����qbЏ��1w��;�i ��7:Ќ�_�?����B�{���F-�`d1AcQ�o,�b��Y 5�d�{��A�l�������;��_�U		'��=;f��?�U�	��5�|��������oWtp�F����t' Yi���g��4�L\C�[�r$�	n��4�F��μ4�;h��ޫS��W[4�[��u�jX�>uW����G��ٯ&���ۚҗ�X9�?�Ur�<�6�O��'�[�F��_^Vj�)7c�1�z�s��0�����oRrNq��t���f�8_Q��2H��q$?��AY�j9��p�_�{�U�6����-��DMn�u�z&?�ϸӮ�dk`��Ķ9��_Ā��iA�5��yv����ꋶ���M娖~,.��^�gį?����J�a���%Yz��v��#K˸�������*C���}�Hx�ټr:/����\��,^�A�y��n��k����>^7�t�L��'�
D':�ϒ����/oٺN7�]����}�j,)Ѿ�R��ɲ�<�2"���	Ym=�pXG��-IgN����KT�lukL�>����L=�Z�zAC�D�F��VZ�q*��'��������Zd���6��7��g�M:�7^X��Z���h�!��Ŭ메"X������x�9A�6�	��O��4
e3���h��zDxg?)��Y_�(D���,49�jN$��˚ůE�C�	g�Qe��f�{z�0j�Nr�̡�9�s?j@Ǳ��Ml�����C\�n��{��9�ۡBھ� 
��t}����|��Bl�t$�#7��57���~����Q� Ll�d��ͽ8#� �1S�_?�1p���������-�JZ���]N1�Wߗ��9�pP���@�?Z����3�U������H]�'��(5�F�kx�<�@���qbM�qZ���(�����|������i�A�n�<&D�V��̒���x%0��=���u���y���h�����kӶ���K��v����yMc�t��8ZvR���֪z�~ń'��rb^����w��{�$� }�i�R��*|eciN��<`��Z-����0�U_��e�3���K�s�֠W�]�M�%�hh��)����fO�3M1��b)��?�]��l''�M����sTBKӨ�4�׵�j��
�����9y��ऻ�����j~�iF�T�M���k��>�����3Wo�`A:�FH����X��p�>��
�/�ii̮����g�DU<�&&͚��L������,(=��+F�:�E�,�0]޾8֗+�_<b�|}���u����X�^j���cL��5�Qb������Yytl��k�ǨLM=��?�/wĉIX=#t��qxG"t#��*ΟY�]�t��7�1��_#җl�U�S��q����d��g&t�znn\��{,!�)B��q�P�P��p��K��M�	��޶��C��μ{B�ZHR���x�X�OS^T������9�x�sS��$����R��ǹB̬��F�1>z|65l����M��h7,��>�ٱ��2�۴QBb�(9Rz����ϲ��>���e�������%�z�8(s�IS&�/hDu5��o��r�%(Z�
���;�ρ@�S]��,R������ڬJ��@!�_��4ƒch���%ѓ^R�6ihJV��٨��{��`��t�\FΥ�E_��+�le��_�o�E'��V�MmE���B��������5FClwh���&�3�;J�K��X���HM|ląv��K��D4y��-��������[�V�~���<Ź�@����7�:I�j����H*N�W%J9�P��O}Q�Kj?�Ո6l���>݉�g�����r	^�S;�~;"���Տ��z�n�f�2�����XBDF�ڦ&Fީ�����>{��58�QkH�';�:�1-Clx��t��i��)W�X
( i�ޙ��2�Ow��9?�׏��0�-G6bdN(�����7�Y�~�{l�vz�������mg5\�#{�����0�N���3������\F��7�H��rTD3S�~s2������:`�8�ER�,�;��[���mtܻ�ݫY�!��w2CS�ܻ!�>vK`���Uf,�&��xH��,9]��c�b�h��R{���8o��K��z���
�y+I�Z.t�Ӽ��:q~W�Pzh�Ֆa�Bɻ���
����+k�]�|Ȫ��H�U���5{O��ǔ|�I�͡��^	��Y+N2W���"�S���V-$�{)O~�����g�;5��d/"@���J��W��txnh�EU���Z��.YL��<G�3�
'��!::�'�J��؉/�Z��F��-1�͸��>�������M0BV��ہ#ׂו!����|���D�Ko�<�EY�4J��mZ�5ԓ�n*��R_�|LMܫ�\�Xr���(�bx� �(��SK��t�2�|�x��]5�Ey�KI�i��c�A���K������������=�	����h�U͡����*�f��� PK   ���Xp>r�  �  /   images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.png��PNG

   IHDR   d   1   ,�   	pHYs  .#  .#x�?v  �IDATx��|{�dWy��޾�~NO�L�L���<w�v���$#a�mDJC�P1��!N��ʉ���RvL���*Ɗ�`L��Y���Xi%����~?�{���}���힝׮fK�5)��ݾs�=���}�;�������O\��ͦ�o��&X�z]�д,��ʊ\|�WW�ihȍ���f?�y�Ѵ�a�t�6wձ��Ӥ7���}��5F��֩�ٕ�e�k5���0�4�U��|��;���|��ݨ5Lk�g�����\7�k�wBZ�K^����60eT�@���àۅ���fs{�R����é9�o���-�	o0�b>_ �j�, աNT�E�X�����V�����b�PD����h4갚M�<^�s[h^���c�~�jQ��՛�6���C�4Jyд�HLr��N�vw �÷���Z<_~���YM�K�	���)�v;͡��GWu��A�,��'hhfGnkT݁�_{���{�é�/D_�$6�f�r�X��O.\����+��!Ē��AAHoȏr�!T)��r:F�"�ȗ�Dm%Oɵ��W�3Ff����H�͢G~+�$n7<��=r��Yt%�omA����AdWV::������(
0�Qd����P�5��9?���1LNNbhh�TJ)caac��p�d�\>/�m����33�������A�]�ő��ҙg0v�8�����٩֞�d0 k`_c��X\ZB(�a�����ѣ8/s���*Bd��[����~�a�5�r��w-Lk�jqY���y8�=������}�r�C&�����I��N��jRM^״�M>�ԍg����(?X�	��X��	�¢�auy�,�а$u�#'�D�Úb���&t,כ�K]�\�f]�o���!%�7�-ܲd���O`�T=d*1�t8��A�yz�aS7Zo�{xO`I�wI����J���M �ǲ�w�u�	�(Ε�+�G0q��:a\�b��=�����cM~u�.�Wם�����(=-�(=,ck���H(�Ǣ�!����%Otw�+�S�)WED�X���E��R��S_�oL��	�h�Q#W����Hw�쒱���_"@�Zǲ�@Ƕ����Ւ�D:G��p,����#A@�4
Eda!��"��k��qJ̮򙴙�6��g!�+�:|��e�_�Z�)�隅��7��H�\�HG���.����~/���MIT�5�㽘ns�dG�"���
Uge�>�`9�����;�_NB("�]��$�/ͣ�;�� ��ea�Ӊn:`t��?�+�a#� �y��:���T������.�`w}8���� L]*��BT��^GY�n�(�J"�I&̺L�lH�ti�/�Pgy\�w�B�A/2�\���܆R��+��h*u�CC!>]*#�b]�u� �&J1�>+�?&<���%�9�]$�.D�C�n*=��Um¥GEĮ)��ǿ4Bd�Sɬ�X���"���ґRr� �VQ5Bm^4u�b�Ʌ<La�卢m�5�\zt%�A�[K)+����ҥ�B�k�糪, ݬ�QS�g䠔P5������S�H��Z�"�oʪ�69��]�r
�F`r�T�"\��#��(
���� 6"�ź��Y!�\���cT���-"*�O�HwXʐ�!T�9��B,�H6�b<7/�r���]��˹$���ɪ'�ůu�����k��R��w!�K�VW@b�ȑ7� 7ʈvxQ�6�zj�+��b�}[ܽ������BiM�%Y<�m	�P��v�ŏ{�eۨ�~�]�������7�C^�#�Mnl)b��.�����<r�q^>��f�,ȭ+1U��wMY#/�N�|.C"�%��-���K����1d������0ot��#9���=E4�\���LY��7�Z5[�SS�Bqz��l9P�Gm���s��(����^Dؔ.��P��G��"�2�gfWq~=�L���;-6�u�5ҏ�>��Q�k"��D�h"�SĒ��K��|#����dr��b�H4�%ѭ�K���(b"�'��-!N/�����|�{�_,X��"�\.;D��h��p�T�A���qE��tZ &|{�Ĵ�3�6����H�IM��fڢÒ�'E�5ſ��_��\��	c0��B��>(��/��U+-?����D��Y*"Iٖ�E��pA�����*Wip��Ҏ�2Y()C�����R9�m�p���"�0��*"+�J�J=����l�Cd����]���b�|QL@q�j&����+�p��f:���,E�,�b��17��/އ����΢�t(1�]�ؽK��hÃ��N�ΐP�[�5Zh$���j'կ�J�>���t�R�`�7�i�?ԫ�֒��h�i�z���l)u:}��ᑖ�k5��ۧ���C�ug��KMkY���Y�W�R�"?���U<1�Al�L�80s�
�h�Z"uGD��NQȤn�{�/��b�~"�H��|��e[�+���
�!ѣA�\���D��.ie]�¥P��8���Q�RH2���;i��)�V�{{n�������"\�.��B�N���C��bn-�����('b��|�4�+\�oD�}�!�~���2��v�R��!T�y��N_X���FS�Qr��2DDquC*�$����p�ًaKqP�P��2��UAC�ԪR��Q��]>����Fw+e���0�CN�3���];�p�Dφ\���؀\�����0K���$�?��$R�m���Y��h����ex�������w�Ƹ�>���Fb��E&�.0`}�Q���{����������|E(�D�X�Xҡ��Ԅr���sgyI�w�E��gr���ƺnᶁN���1�:�8���Ȥ���8���yg5W@SD�߸Z�փ�P&�Y����$��iM��'�)�ծ�!C������m��CMGQ����:)�˵ֺ{�%�-��s���xj&g;}�(D-���'���.�wee�1��ư�ɪP��Ӌ�5	�Y�B'�P�ni�T���4�e���q̊����&>���_�G��uEB��o�#:V���cZ�coC9�#�!�,��3�Ю�ZADR4��ٲ=W��i���7{GGF�$�/-��4�J��L�yPG�笋�,�v!��!��V j\�p�GS�9:tY�+*��̨�-�t|��wQ�����ĕ"1�:��)
�n/����0��_����=Jw��k�wcp�%
ZEz9W"�q�h0���~�ד8���tFE�a��b����8[�G^(9��{h���ͤe��H��Nn�"f��fE������;fz��=A��r����ZΥ��ٻ]d\W�o!��@"1��X{��Xz���_?�B�TU���ۏ���B�CH	
c���jc�����s&�EMĘ������;;x���um���\Q&j�x�j]��5Ok��ɺ�P������T���&y���{@D�p�6�vw�60��Gw�妎'��P�+xO����ps�I�D�q!���@�܏�?}�P����ٛ�c�&U�ײ-0!�r͂��|fWLr��"i�Kٱ�.J�p����c�i-5���%�uu$�5T�oˠ��H����Z���y�a����
��K���r"��f/��	ȶ"����_�"����R��-T�4������J����/a��3�'��s�����sO鲥�����Ṅ��=�n^e����B"H�D�AK�&z���^UO����"?=�Ӊ��2J�+h��=�D$��H�����u��{�@7ַ�j��g!%o�3�j�f+(�"0];2-�.����8�_��_�ן@����)��!���٭�%�^�ήؖ��3�!�b
c	?�s艉�0��3��(�D=N:j8�яb����cڏ�~*��'��t ��`��h�o�nLtca3�D��,B����I6`uD�ٰPsy�����Eyg�TCI��)qdoL����&F�!��+�w��l��ld���GQU��~�u�\8�l�w�s�i�t�|f5�G^\���k�����3p�8�?�t�h���V��� ���T9
�$d�+G=dk;y���k��فB��V�3j���johT�-k�R�P۸V˄"u��K���?8��ׯ��V�t�զ=�J�ڈ�\N1{˰�G{�Ss+����x%@�{ؘ��RP5���QR��f�f�g5�E�x�62�\ �r��������N!�3R*�j{�~%V�U�zl���w�������%��'��3��Af�t6�̨|�JD�K�q�C���yԅ�F�r=�v��2_�b��k�xS�0HX��Ⰵ����c����RNcL���x�ٗ񫷾�x��s�G����-�".�9��A����<4ػ�*����"\���Ԣ�lq׸l7�ہ�߇�D{=���C��^�TɁ�BH]fq{��w��W�XJ:���k%����5뚋-4�8L!�:�~�����x�,��I�����p|H���_�����b���݉}�[
O�.�t�T�,��WIps�J�!��x=�B�ob[��j���1����&��f/�-�Ft3&�!�nx�`�fY&4��u���ģ,�9~J=�v�f��'^��>p7�ϹY|�k����|����8��;nƽ_~�r�8�K����p�/�ŲP/s�j"��N��%#\��D����xV�8n10�]�!�{�px�������e�n��-��>��m;D�̕-��ב�_{��B�ܩ��_��������o��ď��z�Gg��g2C�p#�]z�B��i�NzA�S��R��D���r��$U�v@���]Iؼ]�W/V��;�콰��b�rx!�_͛��fْ	'���,�������?����?~��ދ�gV�Ȣ���K_���v<��ϫ���~�x�sxaa����#	�[M�	̹�Wn4�)����Na9�)�[-�R�PW��S�s����ѦL�V)R�Y���Ĳ�ƀ��;l��j>4s�̟na���ȓ/�)A���.��K�
1g���R��G;����_S��4-.&Q��>h�������ž��>��*�O")������Q4}����%WV+��6BFGG���>���U�R�v�p�L�z���Tc� �ɪ�+��`23�#`|���M�w�x<�+�P�=�kT�T��)S=��F�SO�,H8=��R|�@���Q���9(�n�޹E��xw�2}��B��c���B��$�����zJ�8Pdu���`%w�Z�1����@�eǌ��ۨ4�D�k�����wu�pa
���na��
�=:N����yL�����{'�VR!)��N`�[@��%=�ɍ���=�Y��'�vּ$�䍩�dm{ϝ
����P����f�w��XIe��q1�W:y��G�����6��M��tv]v��Xˉ�<��J,ߘ���>��8.>
�|��_=�WX�D��~'�ٯ~�H�|���xdjf��>Ni��:LQ^w[�Xv۽�gD�������'�l �^�}��JK��6s�9ж׏�8���,E{�5r'���~���uյ&�guwv�:�p\\<��c�j`u�E<�O��N���6�ʶL�����-<����S}�puA�?�'����W�X�=DH۟Tl�j�۩ ��]��@�L�ǽ�\�������m��I}�q�cv�U��C�N2{P��$N�N����;�<U��4p����[7���(�Q]C����alb�Z}�}l�F���au@��	�D���S�[h�Evg��X�k;^�^h���V���g�-��l�5���<o��3�e�>b�,vZE������C��+����7���9s�i봕�%
��B8UG".��P���JU��fg͖x!P��*Ң���ZU��#��"��Ib�����e�E�im ���X�u�p9�9z��c"��
��ф�:cC�D�`GH�!x��f$��iJ�ch��b��m)hM��Ʒ~�[>4+>�3s+eC���}j�-��$��u����Xm���1������ut��^�BY����7~7�����{���+����9@��9Ãe#�O��?��֖pPC(Ɖ�x^Cѷ�7�;�%\��i�l��:�H�sH���::@��0�G���Pg1��b���BŚB<�M ���c����`��˧_PQ\"�ͥ�9����_�
8�o�)�k��?�Q?��3�U�\2�4�,�x�u�����s�>t�B�erPv"���:yD��{Q��DlY.��ݨ4�0B�B��ya��0�=xy�������BIwb��B.G��h�x�R���G�\Q�W���nLt�{���Xr���S���ʨ��J�0��y�I)~��� 
b��Eɦq�/���g�j��2���Y�C����s�!ļ��,ƺT�J8�}.r�UǓR.r.$"k��;X�xW3�
w?�<��������8�=��Zωǿ!��K���Mv����� kn�d���g��Z&L�����$4� �?�a�6�ؠ��,S#/�V��z����Xb���i��>��#X�[E�j���E���\�����1��Ry��|��re|~�k���L=�`�k� �{Q�)v�2�a�X8�tY�/���@P�s��5�)8�K.>��yq���fϟ���)�(�|���3�#��x��C~+� *�]9{�,z{{7�B�V0,z��#��5ܘD����׿��:1�(�n�XvY�-eZ65���7E��=�Μ�	⚁�|C>~���~Y���$�g�U�~lȽ?:�B0o9׫g�&�v�n� �����
�צ4$H��v_�i��H0�؄Lq}�!Y{�F����9�N7e:V�ί;�wM��*�y}2Nv����d�E�땺��R�����`#z?����
�-?=��d�x�r�umy�_]} ��'7;�����o�F�[��Kr������l#�`0�B����pH9K5��z��133���qL�o\X��)�1��߯"	bũo����9gRI�~��ȅ{୉�|����p��������a�$򻾾����H���e�����o���j��K����4"wߏtt .���a��2����oJ�7�g~[���)�_G�Mw!;J�~E���Z��wO��$a�O�8�t�9r2�jY���K�o�5"ױ7~�N(��1w��v��0��h\��@�1��C �DL�����[�E��:�N�(u=�a1��� ���f�e����(�&n��*��qՎ���G�J����N4�.�W&2���8Rސꓙ�������/q����R/sxk'J�n�$�1Gd������/ɵ.�{��F1���*�\��%�����u�\"����lQG��	�:�0�ힵ���j����rw����i���s��#�8��wn�~�Ĵv��m�s�:M��םb���M�o�8J����n�p�Q���:j�i�*�    IEND�B`�PK   ���X�GDU7� �� /   images/d628d844-ce42-4e82-be63-f5fdfa438334.png�wTTٷ.Z6ݢ�@w+���6�d$g[D$�䌒s��
[��,Qr�PD%I���"�Ud(
��Cy��w����1�p��[ٵ֚�ߜ+P��T�~��+�����1q����u�,��oT���g�����{��%���Ώ�����3-6������k8Y�#��Z �H$������gn'W�D��5�O����5���?�9t	��T�;N���h?ڏ���h?ڏ���h?ڏ���h?���-`�9����t졚֏���h?ڏ���h?ڏ���h?ڏ���h�W�����w�>�d��c̯��nq�������\<W�^�)�����WvK��[���<���N��s����vK`_���jv�z�n�����[�o��p3�=E;G�oZU�y#3�{��4�.�����o$��0�5"���x���ȏ���h?ڏ���h?���Vh^���a=)n�$�pX޿���g�\�+S�(�6��](Ӏ	�N㱒�w�'ӪJ�����K!�:Z#�|��fXN�Ĳ�_���F�cv�n�|�؝v��T��m�"���2��/�r�f
y���f��XH����S�V����z��y!�R/󘭮3���g��o �3����Z]fk�>�)IN���;���n>����9�}M_iX�X
$��D���������+��\����4�ͩ<Ƨ4Ƨ���)?�Բ��W�`T�SY�V��o�j���$������eObՕ\���Ն'�k���_��_*K���5�\��ubK$��G�0 ƓT�g �\���	��i5O<�yfMQ
%��ޛȻ�T�����ښDq���F�{L�ڈVav��>Z�f���Ԑ���dC��^��?���~����~Z=Ͽ��%.�
�d��m�%����_�)��$��e�9��LM��#����s>s����4Ҩ�S�n{��)���i)���;�z�ֈv(�]sh!:�v��|7����e?�o��O{�'�T$!Ћ3b�V@^n;^Z��K^~_jҤO{j�/kM���u�<+F�K��)��{yY�T�������^0��,Sy�/x1j�N`!�X��6'C�c!sB�]����E=	��CMf��]:퍹����jؤ�gq��c<�����Q��.V�Ϣ�e�C�J�TʌquoA���Gs�������3�9-C�퍽.��>�ٞc�}���E�'���q���~gJ��^,�)G�M�O=&KyA,�$k5�呕�������.���5�9�Ӹ�?��6 �jf�����5��� ���˔��l�2[���	x���r����!-y�79'�f(K��Ȉ�cl�� ������]�R�?�g��EW�󝲯�l�]��B���(�	Q[�%h�yM^X����/{�kF���Xy�ZӤ|*p�W=~�
k����N��s�?*�K�.?.�KGi���>4��w��r
�C�'�8ܖb��W���Ȝ"iIS������)�3���/�c�^ֿ�����?�;�,XF
��ߋ�T�:e�b2`ȴÏE�n�m����.	��Y�Cj-S}�22���k��ͬp��@8A�(^Z߼-�H����$u�l�rg�a��,�:2#�'6���ϭ|��j��^�>��=�G�O)�*Yf��mڎ���FT���)CM��4Ly�'���>G�=:Iqc�0N����M��9{��I~Sf'�߅�=�WV=�,�9��Bed�H��Hbל���KN�%{_/����bo<��K�X��0n��U�����}��8f��
h{�춡+1#�f����Q��!Y� �!�~9/{
V2�����qK
n���X8<�#(c�!(O��m�G
� x<׎���������W���Q��T;4�����3���~6HB���ۄo�.��BF8�l�0��ܹ��G�d]y,��Q�Gx��8�oVSR(>'��q}�%�"�L	�5�#8���R��z�����`K���t��AygP�����A��yB�#'M�S�=q<�5�t�N#=�� ��|t�t����tS��r�w,�h"��J��\��.��mW48,:r����[C�":�ڠw��ˤ����Z?�������DIx�j�s�Fk)ec)��!#�矂f�e����ؐ :�7�&��l3� ����	D՜����~��x��`������BM��	�A��]���&�R��l�Q�ZD��G̅�,V�
�5Ͷ�"�&�����F�-�4���Țm�&����6�\z�Y��8������WF�y�×�����٤3J@��g5��ne��ʧZ@B'=֙��(��QÆ=���u"��ƫe��0����t�pt�����(�wL2Z�B@#��}�ݯ���HЫQ���Y�k�g%��Ǹ_l,�p<~�q���s�U��	�����<��k��9�J�7a��%�ԉo���y,��v�*&�?d���\͗�o�~�b?g�}d�џ�S���X����M��p"���������4�d��<k�z*q�A[���R1]��h��Ē��F.afG�ec/@Q=�mt�|&�caK��q;������_;�?#m�u��I���*_�U�+�ىPo�<�?��9�
�:Z%Y�G���6��^Kt�) +���/Ol��S"N[ɤ�~h�d=�n���;#ЮB��C���I�����	�|�`/Na�z=�w�s}�#q:F�����d-�F�\�b�����r;�kM���d�� b�B�q�
�hd���ȡ��k��5��]�Z|�F(>� x��+獩���"��꽡ͲZ�Y��:�m �w���-��|J���:xH����rC�p�b�@#���+�2sy����Ȧ2�וAu�"[�y�Hm'��};���� 7����z6-�L�ג�E�V�5Z��,S�-���9���JEF/,�hx�4��6�T�cޜ���z~��j���I�oGNoS���{h�͛q�v�~BW�O���	N5��≡p���Qdw@�?��	��¡�9Ц�PL�u���9{�F�v��k�z����iw8��_�P���5�@Pkհ�����_���(j�����Ԙ��5e�5�np�`�':2{���`�/���fج�NwbĂ�Ưz�����drQzDʆ�����u�B�N�z�d�{�T��9݄jy/��v��F�	��G	`cS�����-Czk�<38jOM!n����RKg8�wZH�J8{>�a�r=��^���ί�i��g�}���k1��Ff(�D�=�kQ����>�;�m�x��k����|\q_���
�*fy��ZDK����R���*i睬��I-n{+�y*� �X5�Z�Ū�����|��Q��34ఠ��0���T��[��P���Y(��Rr&�6�!��m�J��kV�])�f��t���?��n?/���`��I �f�����X.U��_�蹤�O/���ʻ�����X��¢ʚ܊��E���*�ApZ���<&�
��9����ƻ_:��6��P=�"���OD|�}�8&3���VT�x}�>a�}�ԑW_�7� }��]�kP��T�,�_�$��J��)���>��Ĕ�����f �r�:N�������gf�m,�&�h$�y���AM�% [!t��b�hz���$�9U\S�Hַ��7�©�����!���m��fs�%���}�n��:�ǖ𲃃߾���Yd�X��݃�A����I5�c��Қ� ���`�y-�vG_�F�^m����q`���U#&#�>0�λkK�����tGP��_�@�'"`�w�	2�d`�NBv���e�����,%�q��+A]��X8��tҗ�a0�r�	FU'����� ���K��%N�A���B;��w8Y\��u���ZB	CBl�Bi�T}��4����!n��!GF> $J�v9�v
����?Ɨ��qF��j���_��CwW�zl6���ԛr�@ 'L'gY���?3��O ��`��*��r�� ��W6%;�VzO��~�+/oP���1z$�}B��'ȵ��%Xc���@τZ��;Y�Di���ݮ[^�cQ�SYv�/ݰu��.�V"P�V�!�Vˆ��h����]�MM?�%uN(e�.�,��l���[�4q�+�oON/�] 0�޹�f�
�x�V������i�ow�Tp�Y�#@N��Ax)���.6�!Њ�;X󶁷�}i6��XeH��#�D)�}��V��k�Sⅅ�D���v�U)��$�����P�c��_A��d�,FQ��E�5����&�K:��s�g�&Q�}�da�aay& a/� YO���F@�$�I�&�#c�Cy��&�Z�u�x�Ƹh��~����/�1+2���%�Gx�%_z
ՉJ���`*
}���G��n3�,��$}�~�n�n�Y��ӵƷ�G<&M[XU�S`�:)c��H��#�_����fd��|ڝڷ�'2�;�\,�jP��� ����0����:�
/�dGGZ�!�q!׋�&)G[q�9)R;<��SNb�ኇ�1����o��>E�&!�֡��ޱTc��F�I������s6�s��R�<9Ҽ�Gc���	����bU4�/F���1��V�.��~m]p?��������� ��"�,sٗ��F;�QBF�=a^Z ����P!S�T-'�f�8����A1݇�$*�Vf06C��M�ƒ�do�A��R��W���fc�3�> �m�wq&�\��e�N<p |n Ӏ ��3�:�f����r�"ڽH�0n�;�$
@�
v;�Ku�H���j=���-��_�ç���F%˞�7\�PQ5-���!�n�"��?�?*�ҷ�-������P����_����Tu�,��?E*}�5��V�.�p�#v9"���3�%��	�R
���'@�Dޙ�����M7�T�o�X)�Z`�����ܞ) ��HX���)�/� ���i��jʨTt����f��e�?@���~�هIo'�)l�(��..y�1�yǔb���_�]w��{{�[]�t��4����N���K&bȓ���� ��]_!n�u@7��s��eW
 �V�E�ǆ��_�;�ӏ�����HR�H�c��/u%���!�b�)����=������:�F���YO��9~:��� !{L�$��O����Wڨ�F��v5��'p�a��;�m�!�
z^�"PH�G}������k5�U�FU��[�%�8�H����o�2��8�uиa-��f�.*	u����X��j�]q��7С�!�,���η�!�=}�����2����qK5���6���;�;���d�: ǝ����:��/s�en��u]���S1�F�Ě�b0p�Y�R�e
�/H)! 6�L�%L#�ч[d81p�[��~i��@��h��)�x�M�~��}t��V/J��eS���lޔ�p�����DT��"�Y��$��2dٗ�l��׎��LT�e�g�H�_�����a큏��I��$�?Y�� �Q"����HȍJ�F���QɅ������,$��򇕑��Ɇ�Z��kl�>��HUyW�Ң/�:4��&L<�������6&:���<&�<B�;����P���Ϩ�B_li��E�K:*t6��e��n����8�f8�b��Í=��j���4�^$]�����	;�=oL� rp?��L]q��L�<
��;k�j�=�p6dk��{�2�gS1�����>Nr��7�#��ןBR&��Rm��tc`<���Ȕ/4C�U��"���X&J�O������o�U��;���]��%�;�r�!�YC�/�U�H#n�'�+W�k�j	�'lO���1)(㽸���<cFZ#�!���lϔ:�F���cJ�PqE�:✯@B�man��R�+�"�E���9�/�0؆��� [��l��w��R×����:������ ف�s���m� ؑ�����0�H Y�h�!k	���*w|Qу���K҉��f�t�﮿�@)8��q��+�r��j	���Ie��)�ۡ�LX>up�ك�xC���q����k:��bZ'��p�Ƌ�A �D_������y��k;�|�f�h.�9��6.�s���zl�p{�1�GR-���v��h�H4����ґ&��o� �����2��0u��6�rHI�Q[og�*6,N�Q 4�$K�x�&���;(_@-T��ӎ�Oy�{9��h
� �)s'�NR}M�jiCxC���G�R$�pe7�G�e`ŉ��B	{z:�q@T?,�58�;�U K�R�$fd��Ԯ&4�ǉ����p��#�f���(ӷthA���[���-W��p����j�� ���0b���+��B<9�D e�;MMdL|Z�໽(��-h�x�H��^�j��2���>#4/��u>�����R�/����=N''%D<A��pM^���z �`n����o���ete��4����DRX_�v6�é�IJ�����ƳnC�_�#Ƞ��M�7
Oړ�Z�f%�3����5��nӰ��rk����,Ɩ<+4�? s_�C����%����+�y��P� �޿~�V��S�N}�̩
Y��S�RQBNÅQ�>�����h���g�d���D�Z�� ��X��U�D9 E�j���r���	��!fA	)�������Zqwh�n3�ސe�jû����G�ztp�CLA���r;�ѳ���6��<P$�9h�L��[��/��o���fj�� ��ɻ��#q$j���2Dv�Ԕ�
�O��<]��}�s����օ��T�����mD+�lha
���n�S-iUuzOjK:$��B�B����>��8��%���PZUI��绛i7����i��\+|����1���^����q�<����������x�͛J��
�������+u���p�� �V�T�SBCu�x4U�/U���|��5aF�xw_��;��=Q���f!T<����%o@fU�+��~ ,�2������w�L|����{��0����/Y͚pjܫ6�+��c�&���=2<&Z� ��� >8Х�sa��3~��7}�pV��&��m�g�^�-KG鐱������,(W�d�f����n�������$!�SF!��hNڽb��t�72М��p<��[L�����ca;O'�S]�Z��$Zi���:ӇϽmv�M�}�,/`�|̠.�@�n�U~�����h���[.�}���>��M;!��ܪ�sQ�i�����P�?u���Ӿ�̴��������:vE���z���͌UU5���GN���l���;`"���Hٟ6���űY8:�wA���]'�Z�����o*S�i@�vv�ȎԬ�_��G����D-��)���R.�3���e�����X���l�Ӗ4�\QWʁKK�Gv��)sR����Г�)�{Y�K�~ӊaշ��=�n�σajJ]���k-��&Q��H6ĩ�ݴ���5<N�lA��OH�6��kJ�]c�W�@��x����H�f�'R�ǖ�9�!:�0�o�MN���$���``�@�D�ξ
���T�y�ogϝ,x�q�d�$Md��w[M� cL�NO�g�(:�唛���L��13��,_	���Z�-l�����@2\��p�&�+�&�2u�J_��u6��9\۽�u�|]Ľ'6�H-�E��&�mf��y�:� ���z�,g�se� {��
�.f\؎MD&{��߇٬	�M�X�Q=U�Ho���.Ąͻ�
	���s;�nB�?a�L��5�����4����/>�K�7��}�������a]T�_�+���5�)qB#�w=��?�-~3�k������5iz�*Бj��fVc~�bI�X\����2��&a_�Eq�er�d�Gͮ����=j��r{+�'��<��{�n�з:��7�6T��i�9��L��Y(GTw��8���E�i�q��i�'2kKLV����������+sP=5�M����.�M�Oږ�yKQxJ�P*b��(��qR�׈�2�Oe��pe�CM�r��fx�֨��N���@������2�7u�%o������=`���$6���"��}� JHFҲ0}j��6L��(�n��S�`u���8���
�M���@�(�4.G u�
��)�+b���b��j^���I��)�X���.��i�FD7]Fڝ�X'n�2�!�d��/���	�N��d��XD�3��l!׾�ۻ�m��Ś � "^�9�5N«���C�xVט�y� ��o¤##�b��Ò��8|�À�!��m��rq�vW��g�{�
j��=Ӱ��uk�@o����[k v�r����5���9h��>�4�����z�#>�S�8�3|��G2Q���A)y
&�!Α���T~���o�aC�\MH,�]��Oߡ88y�������`uL��bAw���sY�����9���ԝ�2���od��^~�"j˖��9`m�(7c���t�/��:��tbl�/eU\,��N��Z}��y�R$z���ג��Pi^��U�禤I)w#�˽�!�[�Vh	�Z%=^i;�D6�d����e�Wr��VQ�R=?���]�M^kr�='�	�<븡�Jcm�r;P?ry@�	/bB�vo)����"!�0�t8�=l��gaS���Y`���NLT6�n9�j��Cb5��@VU���zA�� �){�J��u� �Մ�'�
�%��p��@I���1{�*x�J��6�Jɟ��>�c�o*w���S 	Ӥ���B�K�Y<�|�fN�D�����0��Ǉ����۫w`sXFy�tӈ��)��5ښ�
XJ��*zۖ�%}%���{��UB#��m�[�s�O����)��keDڴ���B����ה{E%g`h�oڀ?x� Q�^C��ȿ4&���0�k3�ةxB��&+mN���DCs�+!��G�մT|X����.�ڞL>8*F��|�?#���q��G!2m�����,_T���b��SjtaP`������^�ʛ��R
7����h�
�%~��0:�g�Z���ӷ�l� �/�W���&�i�d�;��Z�֣��V'�G�7��_Ϟy	�L����\��w�ӱK}#�)��5@C�#�3;ycT�o�����_�:ё71��#F���+
���B>�tON�������M-m8�Jk�=7f�g�`?���TX�Og�d:O�ߥ
\3��\�6V�+�z��{irn��"��ʞc��R��v�y����`r����K�4p��yQ��Z���Qȳ�C����HXL���t­�~��T��J�~�i�l�t�h�N�r�jo�����`z���
�k�Ȧ�B�QN���-5��*N���7��Ve���*&k�	iᰲ�2�Rg�`�M�U5yr&�����j��a<\վ��o���p��z_�������s䶻�@Q�]��x��c2r�~+Z*��k�Hl�2�]0ji�4S���{v4+b��Ն�W_QF*v�Eބ�� �����Ya�O�%���w�7���u�cW����:�������j��]J>�,?�D�j�2]�5��l�J��qx�qz�@���C��=���H�>��x�~��Po �:��Vf�4Y���gz�ܦ^�kK�Jy�!l�d:� ���A �x`gUMRYPhp������t���A�nTN�~1�lb���n����I��� ���h"�â1�n-� ƽ��d�-ݡg{�N/+�JV��)���U�kgz��a	k=ˣ���gV��!�M��	G��݃�D���� '�/��$Jx�b�T!�gL��mz�qÑ;�u{���h�����  ��	CgH��_�5V�O��-H�U���0ғ��TDU��8� m;�L�U)#�|��rimRî�S��)gn~��81�t
'm�XV(6VV�OF9H�n��=�M���v�����;'�i�oV�Y{�2�rx������`c�pG�����^��K��+�e:[;n�T@����n�T��	���I�&3��9�QeGQ�j+7�Y��<�u�fR�Ǧ����d�	�J+�W��j��S��	���z4T:�3����ۇ3 19t=�쫩X��Q�@�f,���2�f�7�KB�"|7
�H0���@��w%z�w+ZԷ'��]=Aw��Y�0+�m}n������JK&Hi3(hEd�Hp�>��#���Ѧ��"-�F��5��!��
g�y&��A�:;���|��������UE��g~�g^l{����9�����Y�b6��f-��c-K��=?:��Z(ͦ`�kLs��/���1�q�/p�6�;��8��=��ڃ�!4����Y�_,2ȵ�a��`��]�A��>e���lj{S��a��CG�����@uv�������@ɷ�D�e".�Hp!���K����NI�;~�pg�A�jA8�a�28Y@�ޅ[�"����rF/C�:��nPg�)*'���ΛVY�+ʄ2L9M�����<�9a�3���Ϊ�uʧ�
Jѧ>}�g)�:i���v9j�F�'�w�^��;��q�(N3��Uk���
����-Җv^�f�0`Mw�
W�#�jBY8}U0.�΅�p�9�#�xJG2R{gx�i^o�Mp�s�Ag�Уw�cq0h�{�f��5Nn��A�,�:2�C�&v��n*H�I�o�����qU�,O Sc�d��6��&O�#@�.��䨝�~�������Jܛ
��k31f�!��%B�y�����TVQ�8Dǝ����y'3ݪ�OP���1��ĬQ�ݼ8&��Ғo�蠂����}-.�_}����yk�؍b�bI5l�bG�̙p����t��?��%,a��6Jo���yN�8��t����� E��1:�Y1�'��������L*�J����δ͝��>&y�.��mF��o%�����O��)�]�I��G��?�3��iuI�Rk�(���+ez�W�AN��\U9e���0]V��e�ɚhS��W ��̊�S�|����3�{�\�����L�r�Ɍ��i��>l�qwY��Z��u��S�A�%i� 4r�9h��|Qnn�I!��v4�2��q�����Jp}-�0��K����%�}�y�Y6�+�p�6��@�3�3�K�n([V�`��)�
�t$L�U�+��#��sܧ\���fm���7�e+?{O��&~�Rö?�E��?��8��3�?���5���|4Um���/�6��o����fR}e�[_lc+��f�C|�����Q�>���]��+�'��Χ��DH��� i�h�@�����#$�I��o �j�����Fm�4�)��x��f$���h��=�;e��z��Y�U������ �v�B�-Y"/���b�a`�{=��8���"���_K�=�,W�`�AKq�Zez���\�t��r�>2w&����XT�S�~��^%\��CWC:�u�Pj��3؎*�O�c҉Li�"����PY�h�hق��zF)x?s덷,qʳc���A^p���2P/e��{�C{���"!{@�a��H	���6�-8b�Hx���u�#��yՍ>K��՚%�?�_y�;Ej���W��7�������e�]�8S�0���
&{�Q���[�4͚��L�*N鎘��]?/�\�)��|(�%��$H[�U�ꀷ��~�u�NE����X7 �h�w�+>1*����DE�	�#*��p�WU��U�*i�#g}�"Ȃ��ދ&+���l��\چ�g�~��'Xg���7�{��j��K<;I >|�KR�n��K�6�M���t;㙘������>�1�@{�-a��r����Zc3����!�+lT{�N�$RǤmѢ�ddD��y�'�'������Dl?2�e�H�s��'0{< W���8��d���[��.˪���;t�zˤ8�s����t*K��]v�d���&dbd*��4��坠?^%�U��Ԉ��M�'j�Aoܫ���
R�Do�sA�!�&*�?Q�ؙ	ތb���b�t!c.��jx{:w�<)�k�uj�k�&�����R2S���7�i*�N6K�ٙ�Mn�����X��s� $��%z��}�D�S�Y0j3�%.��8o������Y�
��R�zn�@��:�J�"��'˴�!����"���D��
��ӽјyv�G�z���i7J��	�A��)(|���X�Avw������b� ��n������+h�P����J�L�J�N:Y�c$*�)W����0Y��I.;]�&��k_��p��5:=�>��1�tv!�:���T���C�s�����=��@��"y�����x}�
r�� 0@�[�_�1����$x���b
��SKF��*!-�G'�: B ���9|m�L�f��'��6���S@e��Хjƾv��|��A�/�L�n@�M������
�#IYC����11Xs�ob�=#�}̫��PJb#|��m0�g8�m�����&�¥�:�T��`���T����̀AiGB�?φ�O��D� ���۸�7cS���F�\J�}��*�"`ę�;��K����������x��������� ?5��-��$�;�O�Ƴ9y`��'��cv�17�)�Z�ջ��8'���F��2Ż\�\�q����:"�z_�������&��/������J�M�'�o�ċ �ԡi������(��������L<NFa���{M�j��X1��<�1;�Y%.9���=U���j��`ڮ���} !�j��v$��p���:h�%l�nY�]@���C������cx^ӏ܂��W%U��)�6��䭦���e��2�$[�K�s�Q�����c����A3�{��l�C��%=9ЬV�@�>YW���a<�-!��� 
�He1��犹��&j=M�:�=�P����Yo^� #{"��q����~�o���Ō�~V_����X�j���tl�/�&)Î��&{q��Ϋ�fo�E�a���t�t,tJ�ae���v`��\"�X4�N�w1��C���cR1-�.24�^��ȕ�kr�������˂փ�Z���?�d����
�����-��}����L��.�i��5n�X����`�{��CU\vW0f%)E͛�e �z�=�̙���=M�[;OF*>q�<���a�2��3
�g{^8Ѱ�v�6�� �d+�~��a�	�����8�!J�����W ���v�Z����NJ��-�h���o��z0[�n�A����Y�hYYh�. ϵ�>����2N�̯�1���zoj!B��3�2^\?2�%��ש����.�r���6f]>�~[�+�XBh`��t*��X�W���O�J�A��-���\!1Y�!aM/�'��ύ���V6�����H��`CO�v�)N��]�9úڙF������<�� pz��p�&����Ƃ����%�/Z�:B�5�W�Ғ,Y2�cg&1��9f���=�O�`��5�I��W˒Wy�_`���s��w�(�F[�~)��8(��;:a��������G�Q*R�t@IlY�8�n(���Ơ����6E����ʑ��]����n�����W0�
h�H�P던ٮ/�+t����]D��;%�.�Z��D�������jt�6^��;T�[���2�׶[����5k�kUŨ>*�b'�)t���چ����ai��n��(�k	��q 	�X��!����W7_�ܜa��<6"3"���3��F7��T�Tn�Ak��;�	�'Vv��/pXs�w�ȫr��p�:m��k�A	+��9���.,L�ݲ������\�[��v2Lq�ם2�>cG[z��)�mo�p�2�Oz�������k��exr�aW���)�*`�/�<�{��HLL��i�V� x75���3u������0P�4+U�L�-��<��o�?3�L`��������S����%`��	����.����	�ap���r:�u��8n22��LĢ����� �3���
6�"z����7������:'=ԟ,�ήDȽ=�N�@5=��s�>�Y��'�I{�,�f6+t�+[o�<�)��Ѣ��ݥj��@v��d��W�~O!�ݧʖvb��V_�Zo�<D��� ��V	��z�\���
J�lS
=�?Q3��Ь!�B&G���)oGv#M��ahhz�]5b��l�֋Y�2W\r���|�����"�/c0㣟��I-�����5���O�݆��?#�!�I4Cqdx�}f�j�z�O%L�j]���"	Sǝ���!��'��U�&�J���4���pqU<w��2�{�2
k 6\	��[��̪��BKॹ�;��,�s��r�]n���T�����`{����j����b�*�ʡ=�l��&I��5�%���Á����-i��|��^H�`(�=:v���]�`'Tw�$?�@�oL?[3��49����D�C�dU��yō?�Xn����l�9I�u�6�Җ.O8�$���e)	�\�@�o� \w{���f�I
>�����X��OA��gm�X�͍9Ζ�3��:\f�.fgҿ�����`B=C1\�&��ݏV�$���"E��"�o� 8�"�����tA��#if�>[# ���׆��}_�:��NM��8c�'��L��I���u�:��?�cu��)��T?�� ����Nd{��t��;e�������	1�t�s��+�-��������������78�,⼕�Jzb"���6ۏ�۪�
������k���=-\۴]����B䏷ѭ����l#+��@�P`&�䴇X�z�?x�4�_���V��h�&�s���}�X@ʚ/SKTw�{���Z��D�L�Jh���է-ȃ[&��:L�Nˑ�O|���-���4
4�&#��n��Z\}N�Z@�y�u�3S�����'�;=CQ�(˻��ҥZ�/���m�[�b��k��������8b�G����;r�Wj�x�ᗝ�͡_̢pxR8����̤2j[9�dC1�vۡ�mt��sj�4����O��3��&ӱbko��y<�H0x7x�K6=首B�\{˶��d�q+����V
�`(�o��~�
l�U3���l`[�O�;�������>L�,�7n����{���%�{6�C���VJHD��?��W�v��R���3�N�:ĭ1W��y脏'\9��t��y]�ZR��h6T���]�z��dqg{`0CX�_��X�eĤ�Fh|yU�T,{+��`��ٿ���F�^��f�����{��A��C�q��;P@{	��SMF6��m�jD.�r,Q��O��}��4S�b	bXHhx�?�aB��9�N�:C�/|��/��4��d0�{_�'��K���fO�r�V����gF�s0{�'��Yl.^��ؚ�,; q�~%74Y��F�*�����:5.-Ѥ�s����s|��?ް��
0�z��\�~��bJ��G��ՠ{���*��v�j�/����o�~'-��]�1�/�����1���N����5�9`ִ�Q���~R�ڃbؖ�%/�o��� ���h�0B#ɇ֞F�ݎe�ޒ˿8�<�*u�8(�/;!li(@�����4�s��w�R�1�*AϰgNE�}��	<��
es�y��=�q�_�8�ݗ901�.$i�7"}V��0��2�x��BKY��g�_������Ƃ�n�{7v<���?!Ď�f��D�B��7ό�S�@2�/�Y=��m�C�G�7_��3f�|�şu|��~�s��<sW\v�&��(�$�����7�ߥm��)���%%F��)�쵌{)�-�~'�{���=��r{�=]��"�G�D�c=������3!�cv���ps�*���93?-�'o��a)��r����{����p�86[˵��[b�6�q����#��t���Ӽ����2�Y��'�i����Ҿ1�t6
HM]����5O��en�Sld��b+k18B5YA7�k!���,:*��W�ĥ��ڽ垈D���!6��>�)�|��}U�B7�k�=v�.A�A��lC��p��� ��&���N͘��%�^������-�A����[�3�_��+�h��D}�ʽ
����w�ఊ��]�F�Q��"��Ho�j�8M���wv9۰�ٝ" �ꂢq�aҡ�~�RN�ߥ��*F���O��P���`|�y4
�����E9)��[i��A2$���ۗ[�Uyp���Qb�̬[`c�/�d��YOƑts{�l�7��y���nH4>�Ҽs��%�+.F�R��x���nJ!���܆���&XSB����Z���vO�M5@�rkȦc�f)��ft+D���������aŮ��x��C�Ql��ˬ���l��M���,��"z�~*r�@
S-�(�Xt$.O�������_T
v�
�E]0ʪ��b�sN��ދ�p��`4)�r������Rv�y'N������HVzV�؆�C�o�C���9�{��=?$����` �����ۅiξ���F��l��J�jn3@��o��4���G]Ɨ��D�:J���J��9�Wߒ�?�p�&Ӭ���w��HT�Qi%W]��8���$ߦxY��S`��$��k@�8:����ހZm�i�t�+F0�eD�!���+�ަbBXj?n��.vrՎtF/��u<t�6��0�Ap�%����sզ�����]G�oU[���������%h]F�]1���~��I7鲺eOR1d�ψqP*�٥�4���w"����aV�Y���n6�~�{ĥ��_$oQ$�o��,f
g�jX��3#+м���p���>P��#Dv�[ᕈ�7/�$dً�OR(�/T�	���=�:h��Y�\�d�\�1"G����G�������.�#$5G���e��ܕ��A38�䵙����Z�5��xQ�k��1S�
�I��xf{0m��M�bW���
�����5�̽�w�����BUn��%��ԭ�����uߠ�;��	���U�o1�^��+O,"���QW���6���~5��}Y�������2������D�{L㾃IS�����?O?�9>.����_}������OJ�=��u?^��i�3��Hl�q���ɻ�L�
��qו�O��FR_q���Xt{�Z�\�?���<DL5�u�3�YP���s�x�o��L}���ʽ�<D@���S�r����ؿ�f`�;J�e�i�
�?e/n�.$t�Vbq5Y^�g�C�շ��O:X&���з��}����"6I�=��T6�w�C�KD@�ҷ�RYN�(%&[.�>L�����uB4KD#1H��?�*x2h�5��7�5KH"�g�ʅ���*l�|�\�
��)L}�"����%[Z��I��`���ց�����o�;Ța�_d��h�x�6��N�o��1g��:;���of��'�`! l/R�ĒA���9y�ĒK������Bĉ�s���hd��Ա��B@(R�s���T�N	�
.t �c@'2���;�fd�oE ��Dc���'L�D)p�X��]�����O�N��Ab Ckyo<h�,C�ݦ#�
ñ$���
'�T��X�&}aCOQQ�I����6��~~{8�T�[i��D>'9Y�J��[���wgμ�j�����v�,V�t�f��5O��]�L�hA�������tZ��j%�����-�U�Ċ�O?�X���q�/�����{�]j9X�p!+zg�Ej&��2���d���u����-[��m��z<%,�6݋[ԬY�W�*F��I�z������Csu,J�ɑ��yW���^�gBz�n�� �D���{��!������ATT	�R:��Hw7H7C�
R�Jw]J���!9t�{����>�~Թ��}�^{�}�=7~�	�j�oC3f�i81 �H���W�#��cV���7��?�!v�ŧ�=J4N�VOh{���	��DjT�N���Rd���b$���J�J=�XC��I��=�G�X�d�r�:EL�& ��$)����,�*A�k��6�����/M��]4� �yuǀ��#�5Rt�CiE�Ѓ�U�6��i>-?o�m:�!tU_���A�=N�5��(�ME��!Uh�A6�]�[���J���ƹC�X����^5��Ĳ��-� z�3�z?��T��8�c-w��E�����ط*�&S��R�������S:��_ ���ƴ��+���؂'pU�`D��p@��hקּ[!{�p��"tu��f�MT�-��D�9������t顸�o�����Nge�飯�e���zrݡq��A4/�1ʣ0���p5��t���G�8��Dȶ���L��u���X�8�ẽ���%j{q� :���l&�.l,�<5ta{���$˟�{����5@l�ʪ����{��hX���Jo#"XA}kh6l�L��q5�tn���s����*%���{0�u �����k^+2����M�R"w�*/M�$��:����ޓ������[���*���=��!��� �"�Nʴ;AJ�2cǋ�LG���웗�xth�AOmΙ�o�K@�e�k��IZ9�-	��|�)t���H�I���.�����θ�\�{I�8�J_��5J�����ا�g��G�w���I|�5:M���)��Aj�ġX�z�3�c�[��+nƲ�ܩ�k��R�N��a�r�HrS ś-%t����.c�
w]�`�G���Ӡ�b�i����&��0��a��\�U��� �V��K5�3 Oj<���=���Ņ��tm�g�܀�ȣz�����s�_�,����*"����d�/X3!#�<-׼&���m��� 88����VMJ5,վ�`�����em�����;���z�~;�z�$k݉��;/!�����]T��TI��%����&�\�ڢ�����SCbp�(v@�l����:o�͟�V�I�u����]л�����!����?�a�<�'��p����ޱv{g�⵵2dM!f��� ks��6�t^��^U�)�����4bg���>���&���w�ݣ-(�q�m�:`C'�<�t1t�9�-O���M�I�AX!VS-,��r^q��RzwO��x����1
Թ
�ߕ��%�T���/�<R�?|�H����o�q!2������9P��T:YQ^;s���/�Ї^���Hrx�ݿ��.� 9$P�
gp���T�]�P��H
�,6f�����i�UH��he:͂tBhe�3NCZ�I3(-�:24���!:�QD��M"�xԥ�^/.�6�LT�&8)Q�+6y����J��o/ �'��>g�jd*d;���y��*[�h�(�z`n6�{[�P�J�'�ښ�V�|��!��������(e��eҶ(���r����o�Az��q�+�]w�Gu/��x@���T��B��5(�g4����ᦦt�׼������s�4( ��U�W�P���(���F��f(���?Z����b�"y�\ƨ��E���Q���Jd�V����k��]��� �?��>bX����le;fM���̥�G:�O��.��rH`b�s���%t����5W���r#�_N6?2U�`G=*�8���,����B�H}�Lb�.�Π��~i�O,7h�`)��o�o���^��8$H{�q��a�4.���;,QҾY�vl��ŻJj��J>M���^��2+R��c�>�B�E�0SA�2V�~�΄q[�@�l�TJ�k�����*o΂w��4i��
w��9�.�!Ζ���ܵ�	?Giv��o�&��F��Z@7�	��&8�l�c\T�+�?��������L�"�X������23:����m3J^���6��\�s�%X�Q��޸/v����ib�;n� RHu'uµ�r~�r���Ͼ�-�}�L⌲K�{Wm��0�/�ڃ�V�j�(�o��w�=}��=�o���e�Vn){�Jx� H�=�8"J]��՚'�v-�����l��r7%ݎ��5���P���W�����6�����2Z<��	��w���L�?�+�	��_=r��L=���@[-m�Ŗ���Mo���_�S��Oᕭ�A�Qu�t����K���z�>�ѵ��y_o�bR62�������%�xj.��Q���a���eB�민�]�����^�kMoן�/���-�9��:�侮=7<�J&��OY�0��-���/���-�@(��m�B�ᣝj1�fk�=������s^LT�o�`�H�A!���)��	����Wo�+����)����jI_���tR�7�Y:=h �`���U�=���'�6/]�-�Sd_���r�#���H��<5b��W��R����C�^&�~-�p1f�o��������?�`0g��?�<�����$�Q���6��؞X9I�������2_��	��0�dD֘�]���7�D�%X�/5�5ܧ
��ރ�;��D,�K�w]d��c�-0��9Gm��H���݋�ͭ3D�-z��f�����xy���_�*��E��80Z�V�e�ܑ��1�-�6C��'�����J��?��\3�f/:���%D�^\>ޏ��#���)�����?��`�e�Ѹge~�ypt�3�6G�1k��

ñ}9�o��4ǰ�hP����`��p�$	K�S���*���ڛ����b�~>��(\u�!²�QMB%��<L���:H�>��h�~�(:��N��-���M�x� I��|�g����.�j�,,�w��;��ɾ@��]�=�#ԥ\�y�v4+�b7ER�˲jaڲ�Z>�y[�Y�n������]Mu�U;H��$��P�#T+�O�˱Y��}ek�(��%R�O~��k6vڛ\�z���Q� ��>�f0�Mݟֿ��ٔ���M+��d��W�~>�����~s��'q�'��V� ]��;�9y6��7Θ��6�9�.	~Lr���Atu�_����P_����� v�.<�E�Ǵ��������ƕ5��4�]4�y�����+�ɖv�QUɣb�g����H�qh�!mãp�;8�|捔W�RK�#�^����; ,��<����n1���-�����6&�z���۬X!�Ş6�>��A�r,���x��7h߾�{��{;QKA~��}R�Ӣ�}}�7d�~B��� }���ϣg��:A7�{p�������������w�y����M��
�ʎG�꺣��!�Ş6$��6�5:�DV�	���5����^��O��R4�_r���m �x���]� �����y�������:n��	U��j͒ʖn�'�͖�)0}Fq�U�I��\jBf���#]B�G?�t�63���{ϼMg$Ĳ?"�ر�&V�# S">-`GX9�\���f+M��9�+�_� ��4p�PňPw�@�K��b�|�Z)�ƅ����a:��	rbӯY��ո����4(K��:�z&��u���ݟ�Y�J�iy�ۯ�Qc��;��#�XaH3��ł%��zu�(�{f�l���ˑ`�׍֚�`tٍ2 ��>Xߵ�_��@��׺�j����肥�<@� �t�&ߙ֒I���Uͤ@�]�μ�p����L�yy�D��f���I�e���c��R:e���4j�Wia��S��ԵV^o:�۳u5H�|�[�,��,���-s���Ȭ~���~�E	���
Td�MLcj����S�|���i�o�C��7����V���}���}��p�X����E"f��O��~��������e6xA(}�¶@Y������XI�/-?Շ�.?�f"~)(׿�V���8}\��PU�(E��eǠ5>�38<��I����
���[�5m�Oט�g]n�<6o8�oq����]t����%y��D�(J8�%�{],�X�u-%s�I��A�����2Y'�/74���C���(?��t��I&>���2-�ĩj��{E�{L���<o��菙WMx��{��e��S������=9ՂX̏X!K���Z�1��Fqa��ه%}�h�� )�=�7��d疏�*)�T�]\�GQ+j��cQ2l�>x9d��T/%܁��lձ�����o䷘�E������s���Y�(�ò��l��X|ak/^�)��B͍����an����!�Z�>h@��dw��F^#�+�~�����\�n����o��g�Gٺ�$'9��K0A��t�� ��ujVhPns��py[ӌv�9�p�<�W�:�3~�����C=^�ogk�"�� ��I�C�H��U�n�QA��j!t�H�Ǣ0=G��x�O��'<`����d��'"5(T�6���Kn�5�J4��t��^�7[������.���
P0�E�ﯤY�?.^����7O1��t�*���a/�1@�j�f�hԚx'�Fg����a �A�&�,�7�r��"9����?����I�tH���H�TX��d�w�M���G+���҇^n�ALbȶl�V=m!�;�AƢ������>{k�H��<(�e�߳��G���f�j���k�\�aU�xaؑ�j�$!��n�a�oĩ�|ޙ��7(/1P`�#�	^p䏄<��'�͉���ﴔ:�Y�>(Λ}�VXUc�JȎ���g5��m���>	u�;3�/������I�jf�xؐ�l�L�)��F+��O�x���y�|J+��%)�(���G��7��)�K4G�*��lͳ�p��g߆�ɛ	��w�x-76轷BTr4n[#��M����PF=�b�������@_����@}������iH�M6�d��U�P5cɓ1+# �J�:T��o����v�k�����oWwj��!TǊ%R�1K�m�{�񝻒~3e�]���Gc�~�k^)]70�~�d�Ԝ"\Q��u�3 P�+��k�o�/|p}�:ݝ�l8����ک7��a4�Ԑ#��_����`rOfN�;p;�A�R�觔	w�qt��ʽw���� ���ͣ�/M����	K�����V?{D���&	Pa�����W�஀l��`^��E��G՛]�Mp�!_v_E�Z�����_$Y�e�L,X���D�RT������Ь���2���O?��Q���^�:hɣ�RAGq�gq���[ET��Z*�a���O�g���� ��Ǫe�~��Meu#8�~�����f+Y\iH��m�,��d8H��:�D>b���X���UHQ���޻vX��QV� C���w}�xD�b�%�n<��DJ�PYd��0<�g�J��K�C�oA�����D�3n�C8�����x �|f�qE��SUr�% �N�{�1`V�W�]~�%@^�F7l8�IR;bV���l�v��~����wv�����6'�Jߎ��>�{��^܅�$E�7H��ͣ4L�C����1�&&/Z�������/�`^֭mC��;�t<~kH=B�۝���;�{k{ё��@{��*L0��'�uw�k��{����º}*<���4���p@ZhR[M�U	���L��	
e��j�����$����4ɜ���;��������*5f�煫b��ªx�G/MƊ?ho���0� w�;�_�&��Y��7�jP��Zm��e�D��,��G�Ga]���в��b,��y	�U���ü����%}l�I}MA���~0�=�	S[)L(�z9�wjc�6 ��}��'�*f��P5�.Rظ�dvM<~V�PiP~%!M_m�w�X1���|���W_��	��D�<{~hG\�#��m%�Pnm�!rl6���dƊ�ؓ�֞ow�zVYa�A���ث���D�V"���d�H�OGq�G�a-����F�Lڠǫ����r���]�����7H�*��f�w�F���+���"������n�W)Qm?�a�{Ǽ�B�֜�[w���),\��+��"vO��c#�Q�{�b��"����jl����;����������iI�9_G�X��K�Bgtt�ݡ�yYUGe,��|.,n��֢��
g����r�ܜr��r�^+eԓ���;�c��T=�.�dR.����zK箕���v���竄U	S�N��4������2m��S��N��׃��-x�=X���_ ��h��s��� Ds=�7E\k�d�9߭\���# u�le>�͕�ſv�*w̋Ö"V2�$l5��^�^�Sgl�[�s��N�h�R��tn3��h&?�����>��o=a�.�^��\�f��ż��ݨ���q����D�9��;c�F'�t��Fv�qa?.�+����j�D=���is�����UZw��n~�i�PxE��gz`��;nU3|y��$�����E����=����jʄ��t�k�|$X�e8�c%#�X�����Ht�G�ol�@դL�Q�
%*)C������Q����+�`�pKT/r�b�������bP����3�-���/ZO	�@-P�->i�Ns�Z(}
�?���zb��Ј����0rP�.V�ro���*��z(������+I�xJ^������>���0�[Y�^��=�����_3x�Di����������T��q!�|�J;�]dY~eg����)�i��QO������r%��?�N}��5�GJ!k�FƂ?�Mf8n�`H�j.>XB�����f;Q�� (K}s�YP���]�M�	`/����������w�>��O��'�����mz$�J6�G���k�C�Ϙ��cP����g ���N�^$W��QA�,u�f�����O(}G��&}����v���=?�|��Z�N�W�%�����{��2b O���bc���'Р74DN\4gk0��>����O�Z̭C �� �sd�jP�[�q�CAM�2-�S�9�k��������)�ּ	Z��Y��_�bg؆l������Щ��Ic�%����"�@I,�  ���.m�Ͻ�q�rlAG:M�N`�?#�R4G���CY7�৘���l����:n�0K� BW�^}��'�D���t��spR�0|l=tDXz��Ǳ.��c�>��.�Nl����=f;��v.|0����O��?,�=GM��z�x ����������[^�^f��Bd�)��巉�ER���#�w�.�m_�#sj�a�x����Ve�U��x�x]Ȟ�7�^eװoH��KC{�^�q��v�~��Br���5/���R��%��� �ǹ����W��������cn��}&F�2К�-lʴ�
LN�H,���g>�q��_�
.��oS��
�Ᾱ�ϙ�p��&d��I�^�Soh��Ɵh^LU%��by�:������*��`���j*IS��#-ٴ ��P�h�ʂ7�u�����ok r�i��σG�n?ol��nj���l�γ�/��H;?�U�G���?V.��g��|�j�_:��CҠ aњ#�#��9�
k\�eC_D{��d����,��ok�-��GG�zG^f�����w�1mPe,1L�tK��u��|764�MF���@��OGIe�Wj���3!�0�;�g���}å(m��A�7%���s-*���6~7���%~R�< =T�s�`F�sEgo��_�n����'�ִ�o>%�0�Y��tj,��A�~`зn�TFY\קQW1l�pz�l�4r�"]�/��a�\P�'c�A�fr�OPڂu�'H��.�5{oH�B7���������>���4���C%ƪ�a��@��=�����s�"!J��i*�D����3/�("��)��o`9EF%�m.�m!]`��H��웲[��VO�/P�,���~s��Q[��\��ocߴ������eHO��.|8dA��M���Mu5TG-�]�bmf��>8_Tr�C4c�
Y6.�4yz\�I�Z>~�g&��&�0�k�	�x��M������&'��ٙ(���_���� ;���L�;C�$��������aj荪K�	��m� �N{���O����7�ǣ����/�=���L�FP�J�����.A����R���]�B��j�g�+�#N�����O�fOp���xO�Y������OU�E3Y�!^^���k@���٬�5��}�Rme�\��{z�k�j�$7\��;D���Y~<Ll��{}k�X�p�U�DB�Pwh�ta�u���O�����²�����B3k�$���kȂ[3��`�m�� \`�-Q7HgA�diw{:�GMf`�W��GF�.���
�u%.�R�m	&��T�͠�������� <���[W]l��=8�s	�5<8qt@4U��Y���D���J�����������(��'�&�!BҍM��{��v���f�tb����e
� $}�NL���� �\�����Ypۜ�7�N��r��W@D�+�t$\�OI��;���E���
���	M���lA]�]�\�W����J��}B�p�L�П�>12�c�A���E�8�MT�2$�7(��o
��E��U=���J�$��Z����Q��t��}@���4�ɻ�+�_���6��I�����I��ųDa֒����<q���'�����{c�K��}2���ᡡx�t�M7d?��Y>��%��F�%G	h��kh�(�����T~�4�z��b��)h�_�ߒ�h�Я�q%�=���{���i{�FA�7�"������V�X�s�r/����$;�]��L���}��9�K����Sߋ�qr<�6�mB���ښ,����	��B��NA�������ѣ�|j�s12�]����v��Q�v�{��p�����A��O����������<��,
|720���X*Г�W����ݭ�%�)�����p���f�q/��}��~����9��I�2�е;�)n0)F0U�a�6�)�Ǿ��&�M�.z�lP��Ļ���e�gS O�!`���N\%c�i�+�������;խ_��b;�Z� �L.��\:�����:����ܰx�ӻ�����,#�V�gZ���l���6����c#)��	���`i>;�-\��Y]:%�Z���W9;�ڲAK`��먳Q�#t��9�&<����-�|G8���r��F��o�3bf-��Da�5B�E�K/<>��!���.�������
YG;��F�9Lo���U��X#\n7:"d�����N ���vOs;ȳn�)�w ��]�p��HԢ�p7H.YK���i�83�������H��[��a���5,G [�G�b���y�6[�3y�2�D9��\mU���3i�߮�&����(��w:����,}Vȇ��R��$�O���=̐&��8�NF�����em�-aչ�؅�
�(�*��������P)�+J<�;c#gb��3ЀZ\�G����:�4i���3)�vd��$ �]��'t9pC�X��8{f����~�hR��o~�zǪ'Dѥx��C򌧾�<�I	�0av9eӏ�M)�|ڦ	���޿Ia�����2B�Ρ�C�w�XW�b�����/���=8a�Z�zd�k]�|�_�^��>�|��/
;���F���"c{���^/0@��o����Y�1�1,
M��]�؁Ң�*��+/Ei��8e֬�%�P����ۓ�+���W��GQ���
�{,1���la�k�1K�,LrU�t0�8�����f�~\�Xb9��0���!��$��tM������3�T�Kj���f�o�,&Nm�=�Y;���5I�we~`��1�X�=�ڣ��B�MVK[Y��f�&��U�K��<�<[�ǜ���zK�"1u�s|�͏��,)��o�mt�/����C5��zU6��D]����Ok&��N�_�Ҟ�&�n�i6�71^y�σu{�X�Qh�_�	(6����l����=a�I�Ez=:�����%l�Iͨb)���,v)Ġ?�.ye��,�d�Ɠ��
��-��QoC6cr���(�,)2~t�7s�m�@��0�TڗO��$�z�0�Ӹ=a�˛ȧC0v�^C��	{�2�+.��*?`��+�m��.�E��歚C�����ֲrA\{#��7t�fLct�2�b�җa6d��{_	��ڛT��K3��?S7{�u7o�e�J�~��-��ß����B�\A^��;�E���R����m?�K:�Z�]YT�C�Q�vz��R�x�XjGœM ���n�O�$��u�oW����ĭrl.���/#�����Vo
��x�)�b�V���^���Д5�gN՗�p{pΈ^�F�%����s��Y���|]�建�0�k�+U��eEn�	&��˻.�HjfH]5U��~����^��+���8#�qq`�1v�Ҏ���C[�h�k��q��<q�����Z��,/�K���g~����5ɢ�c���-���bh��3�ԭ��XгK�=�G֞
�1��Z���h��yyy�L��O9����?�פ'$4�5���q|�i<J�亽+pL�9WCm�F)v-^)���`�`��?�^�ag�n���j&E���vvFEQ����M" ���=u,���x�4�ſ:W�ẘV
S�+����U>Z�-���cy<x0λv�y���9�k����xz�V�j'�VV���R�]��}X�à\
��n�a<�=_j��ܞNU��kˣ��Z6�*b����\�{D�p�\'��!��V���*�ESZG1�LP�c�y,��fh�R�AtB�j�t�ʃ.mo�{��Pc.���J��۞>'ӈ(�QV7���;��F�QU��y��-j���m�~PG�|�>n�kn*�e�#fz�4��LE-�(� ���V�/~��?R�(�Ms�K%����e�L��d`w��Z����/���ݗC���G�O�G��d	���j9դ*"�"~S�.���gv�p>��P%��r{Z=��"���l1��e��ֽ�;+�[��}u�ׇ�x̥�*�0lN}<Y�,�t��Lw�[Uəu�K�>�si۷Ծ�^�̻��#�UC
��9y>V�v���)W���B���e
A�q��H�6����?�Lds��"ڐ�v;Y?*��й�=�|y��U��(��Q����o󋨶�a���\6�IP&`R���5/���_�d���oyA�:^ʆn��Y������^�P����|Qji*+�ɟ���L ��L�Hy/K{?@�{��b��s�~E��f��lJ#�7��\��\
�t24�./����qR������m�E�F���-ѫ^��SOMwI�X�-�`щ��<�pW����LA����?��6 05;�1GU��P����
-L�ܾ����14{N��Sk]7,��s�=�;�1S�Of��WW12�˩�P��o���ƆEmJ�G�|�Aڃ�4T�X05���5�C	4k[p����C5�Ч�r��$8J8�~���H�����L����^���j�YܒO���(�]P6�H��=ef~�������"� ���/�^�����pU�'S��|�C��_X��ܷ�_�æά�$9x]�%���vv~.�y;f�f+<�zy�]xP��)�A��l�R�39�%�	:R��<��&-��alGQ���	��ߞ�W">Աh;L��`S�>Ĉ�w$0���j�#�Bѽo 7���Rr�q#�u�V4���ON��[#�PowS��5�������!}c���ӎ�C���iU��Y��HĆ�C}R��P�	7���7�ӕfɈ�l'P�L4��G�l�o���f��J����Q����K�����U��]g~������ψ���y^K���B�w�w)�s��q�k��M�ĩ�L|���{����κ{S?����ԥb�`����|�و	��Z��|t���;0�X󽱝5�?��P��m������4"�^M^�cc`.���=KN��r��W����O��3$e�i���L{��S�}�;����"���ꃮT~m��	uy%@�b�@��KG�'��#���N��m�'�/�b�$���E��5���y��^��i1\�8�)�$y���� ��IZ��/�Co�Y<���`�����6h���������;��q`����'�|����WH���itF�A}�2���F�M�}�Zhz�@H���v�Q#�\��T����ud��\�k&���*V+���.�<�G�n�x�Cb�;��t�6�P�kXW x=�e?V�@ނ�ꍪ���/H>m	���A�#�ݎذ'_����#��~@v�,0r)�}`w�ķ���S���ݼ�P`��f["��d@e>1R�P��h`��emeM�����,�}om�����T��%mE1�Gߔ�9Ʊ�v��ؚܑ�#pߔ '��V��m�l9?�Pk?Z�.D�R�_]���;�$o���h�4��-p��ޒ�V�m��΋�>�۾n�dgU����x��Sh�$�_��șZf3�R�:��C�5�x�	�k:���L1��kv�4���&���ֹ~k��HVz��\S�(���d���idY�e3e�1x�o�iʒ��վ�_H卌�͸�W�1�y�M��9k�$>m����i� �\��5Y��w�]d�e�I6���;0P�?c(�����zR�kӇ����"�r��FҶ��ʿ��a7�9V'�L�;a���?t���(������j����gPVف�W��q�$92�A�	� ��^8]Y=8&E�k�E0��I�p�}��!����RU`����7�����;G�5�L�U�P�k�.g��K�wK�o��8�, ͑�m������ ��Յ��J�#�X:��p� qVS�����s���2����h�H�O�N��ȯ��U�X�*�������>?��D�(҇����ǅ�1��D���pr�>��ŗ��*���mOA2��.Z�К�Cy�ޟEcB49X��(�Z�HZ�fZ�Ju��f���_6�6H�8��dǠ��ɮ�*�x��8�Ã�eo5Y��M�հ T����r,���8��J��AV���ʜ�H�.#m?$�%�~�4��)'�;H]�t'qCMF��a��*�L?�@���o���T�dʅX��a��S�Ĩ�8�}�����!���5��}�!%B��[D1Ι71���N^My�<��U�V����\�qTL�Ov��Z2��7�g��ݍ-��B~���%���R3���+Y�9??��fe<Es3mZ��'
�������6���C��������V�&��gf����Gm�Zd���4!�b�B�]i_�N8���\��$6���� �1�j&���v���Rr+ܠt%�X�W���ͥ�x�zꕱ�,���T[,����d��9�����¸��w���ކ?�y@1N�7��B��J?$L�Nu��F�H*���LA0��a�j(Q+Q��o��� �}���0ƹ�����)���1����Q���k�2l��	KҮ�̄�Ȼ������u�n�����H��z�0�'�f}@�
rA&��"��*�.b=��./�Ŷ*�V��k˵WPa�l�C
�]�KU')U*A��x�+�6�Y�mI���w�]�L�2B�Deި\#�3ɔn��j��~��ӕ����{v~��҆&}`��ּQ)O�������#T1��C
arn���E���}CP�m=�3)>�h��+��{2bZ�R��C����a��Ո:o�m1[�f����M&*%JT�TRn�~t�쾢��be�Wjf�0��.��y;�'n�w��O�E�F|��ld&�Zʘ��m��R6Z	Ǯv0_���Ft׆g	�u�O�%��3*�|�u�B��<P3F/`��;�'��ƾc����e��8e�F�Íd��~e��T���r�Ԙ����{MN%�T��Q�O���F��v��U�D�>��76�8�����$俯Ҁ����Ŀߣu*�I�R���2V�����aa$�l�_W�?Y~�kޤ<�tW�6K&��yHo��;uv�SQ,Ϫ�Ang�X��3�RC��R�G˰�� �ogK,fm���^L��3�J�E�\��0,�w�'
[(�?؛�*3�Zd~ �l\��r�Rvŋ�Rb��×w�w2��P� ,�!�
c�X��/���D�zc��b���ؙ/��YH�47�
Oɘƨt��^�W!\`����hG��x�Y@"w�M6W��k����e_G8��)-��1L/��c���@Pf�<��V�.E���>�p1?��u��gzr�c"HR3ܬ���`\G�IcX`�X�I�Ӱ Tef���<<́%����cc��I���07�p�>�W=d���\����o;
MO��	��^�m+����Ll�������A1 ��B'�9��.K��6����3[�*�%��`��~,L�������K�vVh�IO����hF���W��0BX�f�f��gM�p�R!�e|������`"�n�Fж�wZB5»o}�u{]v��I�Q�7�����2���S���D�s��Gv����ɠB��
��f��H���1Q����WܩN;ʁ�(�\���t]��#�Up0��դ�dp��R��5h_\/S1L#H�{�e�)`�ݣ����#Vu��%R:��F5�>!۾��˩��A]@���Ͱٝ]f��tFｈ�5 �ZI�S�`��>�`�E��U���$�jbK��[����Z;�Dd궷��� 1�P�A��pW6�~o�>�W����XzNd�O���H�r'4���������e��+�FH��@���RDNC����Y�Y�i;���5�*�O�d���9ޕ�g
�Y���e<11&4.��7v�7�j�7��*=�5TAkR�[�8E5���'Lob�����n��v�!��� ��c�lyE�@�l���K	��@���G])7E��>|�e9��4t�n�b�=�=a���U�d=R����Q��qR�U�n'jo�R��C��V��^��*�X3��u�Fu��Ah����#t���T�J>�Q,5{�!�½�*8�%?t��)jlG�J�#K{Gь�]f'�{�����x�I����ޤN.˟��UJ�BĢ��h�~v�Э�a��d3&"
�tP���h�L�u&@xn_tW�>���ȅ�d�;�����K�\�f���Je��ߟ.��)FP�X����'L��4_��Dy@�q�C-��w@]�r�r��2�A��Y" k�;�Xز5���;�⤟�5v�?bQֺN�V���Fz5;/�~���γ0�Y$$����s����׷=����o	$���KZA��5+��p�0MZ��N�;_M�\~w����V㋨K���3��,�vț���9�X �V+yOҬE:�e&?���Σ3ϡ⭹+9U2�U����"| �~t���y(Vl9}��W��b�W�;�\�c�ò��U,�ml�B��"ݺ�AD�j+��1�9������g��+��3�c���l����w�2�/%g��^nG"��!N|{[1om�������A9w+ʒ�T��]���ȯr�9I��~��Xh�{$rtjE5�	�? ��J�H���ņz�$w�g���v�*���L"D�V��;����L��(�M�8�l%�&��W]�A�W�Ki��wK�4e��L�ȿok�V���o�Û�eǙq�q�ȝ�ޕE���N}2�` 5Y�M������}kw��gj�a/��,n"����{����2Kl�͝9��fړ�e�$ᆽ�`;.���iIe)�Y��8��գ ��8X�SK���d�!�@���������~�m�0�@��/���d��y?�8iFF��S\/��}�I��^�ު�"&�OA�&�7�O�*	ZdV��eA��p�6l�^��B��I]��O���O�.}�\O)ܭ�t:��Ô<�-or��K�t�A�Ǌ!��Sj�,�G蔓�����KF=f�顈�oy|?��qx�*[�i&+��(*z�T�u�u�T��O��9hF,�T��g>�۟���]:���V�b�h����_����&��떁3�zPᏍG�	��r�wV�1��Օw�4�:Zs�s�v��H�F�B���?{I�,�����m��]:�O=�����l�����r �񘓧#��'ϝ�cz^��f8�P8^]%*\�~U�Z��]	/���ʯ�cPΆB�U~<���"��\�2���<���+��+�K�bm���=��\x,�3���3-�V�V0��6��A�����n�D����j~;x`%gс�?�HA�d�M�/�o��$��*rEW������c��:C]�5=T����3���3��C�Å#�!��f��]�ۆ��rgu8��}ߌ���~NJp�P�����^��Ma�]�W`M�?���Ҟ~�Rb�^�z��X���/�w����T����l�{X|:�<�����(�Ry�;M����h7�.9+F����>�]�歱|��'*�v��I�����I}����94�3��i�d.v�2
��q���	T4�XUĚ�`�f�����2NL���t>�Qk�t0�B�c[���+-I��W�aP�#K󸕭\_��z�@��-7��D�Ǚ��ȞXv����B���y�[\�eZM՛��H�Y�;㫁k����X��t5�:���i�%�]Tӫ̈́<��rߴ�{�~�
7��Q�7�r�т�w��_�B�JĐ�8w���u��x˩J�s���j�q����+�BM���C�?��*�G����oʛ:"se���\��@��r	�f=���e�ۻ����v�V`DeH�ExK��2@[���K���d���Y.��ڥt��ԲVʝ&�ј���������ڜ�/OƠ c`]nd�x��fޑ�����y�q���]�o���b'"����B��ގ��ld�$�f�$xS��V�zh1W����(aߵ���Rh�F�Z��ZrGWG���)���#�K0��8
�$�6��wEy)��o�k�(y&x�EU����9���uʻv҃�;���տa؇m��n>�T��a D�i�\��(� ��@iW�u����WD�oƼ?;�+6�N��S�F]�nUW����@s�����O]��'� L2ً���ߦ]�g,�8�o5A���$P�T��Ȑ)z9I�8�l����	���|W�Z
쓧=V�1N�bdF�~��	�����79]Y��T���� $6Ɖ>�LE���g�դ/(W���?Vz�,��P~�=�M~�_�;�9*D n��U��#M���PR:u�≥IO]rV���o�<�z[-�\��&Y/45�,��7�/�(�m�k[{y������Y^�SI�׳��	�]"=�C%�M���s�'ٚ�v R�M�Gu�Vrvƃ���2N,h�E��P|F�\A�t�A��E�}���7j_*P�j��z���9lÛ�Q[Y�Q)�މ�����3�Nj�h*_�/�<�K=�l5l�Z$��z��HL����?�ӂ��S���3^
�*w���7Ģ��z���^����.9,�_�j�C����� ��P;�٨�)���Fׄ�r��Lz���O��2�ݗ�I߹3��fU���r�$陫���z�(��{xXVp�`3*QA@W����3��$IR�HN�$I����4��<���a��}���s]��s�=�������nK����f��'a��pF�{ּ�&f���03rx<�u ��`�oԳ�p���O��z�+)*Δ�>x���Ѵ��W�I �X�g1R}=��9zF=Oi��۷|0�f���|@�iD}�u8� g^0�^OS��`8�HJ�	�������pe�?e�P=��ĺ�����o�h%e�2V��7�$�=꬧�ؙ�>�Y�)��y��H|�*ς�Q����#n�s�hjOE�8�s>[���7�8-_VSX�_�u����65U�16��M�6��f�k݋�j�����"Y�ћ2��_r���Z��5��6�h������,��T~���%�n��(a]U�Tja��f�.�η}f�����T?3æ}�'J�t�� �=<ò*O�Ct�u�Ps:���?8Ѿ��^�ޛv��c�c�	���3e/�>�M/̅����ŉ{�rZ�Z=�Q6sm$vc�5�(`m�2P����1�ٱ� �T{+?�rPm�6}i���)�ĥ_�'\�&�rB��#���o�T9����Ci�����ZފcE�dg�W��sU]qL����a�Ms��@�p* ����k�MWUD�$u���<;7;�ժe�;;�g�vДq�)S������1���E�y�|ѥW�,?��x(�Y���[����|�9��d뛞L�u,�4����tʬ[��ð<N�p�(.��
���I��J�Ȩh��_vM{����3=I��sX��T`P	7��Iˎ�͇<�I�E�����}�S�� X�m���ӉN��]ݿ&����_�5ӡ{4:k�����z�x�5�|8M���:�7v�@�d0��V�ڞ6ۭi%b��G$.�-�Y�Э	�v.9����u�vO���*I�\���,mǪ�1�����(��2���&��G���j�~�	�F��|J�M�9�����l��A	��9�'�����w��,RY4��n�{߶-<���G��z���1���nc$r�Tt�	�9��F�V�5㢰5���_����4m���'H�qŠX�^�.�1�z���gK�I�ǡf 8���׮#����<��ư���P���uQ�Ӳ���'sOm�æ��18�e;	����1(����;k쭛1P�m�دmoi�6�E������8�8�(@��6�V*.q��T#�J����Ǹ�6�_����(7�W����))��q/�%��l��B�������|�s�#�ؚj��蟸ab�$�"�)�������t�*�ܣ���6[[^����o*'%o�k/oׯx������#ʞ�$0ks�Ӡ�IB��66�i̥5���?k��T�����sG�vO����N�����(z}A�R��v{C��O�뱾NУ��^V� ����ņ�t�C�(1�(�4WY�<��cW*
�����6�rQ��qZiz��c;�4��
�מ��� ���ԃ�J�ě�K�@�l|��G0
_�,E�������W��0��
���pm�����`܏C�%�u�镠X����Rps�����t��hVn}l�@��Dg��Ci2[�ffP�~���fl�W��ofҴ�]wRP�r=���|��M�b`���2:��X����_�jr5<���閼���;ZcƊN,|�*L��@~�X�0u2>-��$���ϮF%�i�+�T fm��P�Y�=c��]E�ȷuN0��1|I���f��g�����8�"���μ��</)��ួ�>�[�*�A�Ot<����8���MnFj*D���P3�Bo�������s�X��� r�0��}5�ߢ�xՈW�w��#��j����^�(�]a 6��������e�L��]�FB���E�|��oŜ��	����A�Lo���~��o#3|�QN�i���t�)�+�)�3o��xM\�9��[H�ǉ雂h�E�H��+�=��f�8r�N7$�D�E�(�U��S#�Ds��S�Ⱥ�Քva:��d�S^3���we�V��jC�y�T�n�KWPES�H[*Hې�����68Խ*m�un,�\�SZ� �J��}��pIn�P$⪂rN����C�'Q�Ɏj"�s��Ď,���J�<�b�Z?Vn��5qnU�L�Ꮮ}B�l�]Ĵ������q^pĞ�z>Ɂ�3+2N=�D`.\`$���H��Pp6�9�����Rمe�Q�� �v������?L07��J?�o�Z�������:]�-le�~�Ĕ������yw�R��O�X�{V̯��zy�P�!h�Ʌ�K�� o 7�eڳ�Q��Ƭ��>J�O�4�A�����)��S��9X�f�/ F�H�m�
B��c�l�k�[j�j,�?����oZ�}`����,�H�H�T�u�.J=�J����z���8ORc/s-IN�uUKPCG��ȣ,K����l���4sg�,�TÔH6|���a�|�$��?&A�����O0���t���ӯ�d�K�ڠ��B�*%�8Rp8��IW��+���'��c�e��>�����83eB�G��t�'jϫ�C�L�fZA��;�
�f 
m��}�4|��Q�Lz���;Ysց��Nf�y�sTU�b�w�����㒢B�����#���ܭ��;]f~��6a�:�'���F��TT+%�ޭ.�?EGH�{�K"&>��ªs�k�cRk{�ua��i}/ gk?(Q�e�՗��
x"�_(=̟��~3�41;A���@4&��sz!�+��Y�4Ղ9 ]�5�J��<�R0h5��vJݚ�_ϥO��B�b5<�i��sC�ߛ�r���b�=�a��&_�)8�����+���^ �;�Sb�7~(�_ �\
>Q���i� D��Ȓ<�i���X��r`��&P��TR��.�kɛF�^�2'�w�I��	���~�� ��5 KyM>���V=^�j��!��o�.��#��>"w�f����S'ݝ��J��q�ف�^�/�F�n*k����#|��ə�^{���+���~���!�O�˴������fÌ���iBX�vW�
k�W���;d͸���dV�����:ɕ2*;T,�͟Ng��t��G�B.�w	_�:�13-Z�4~�J۷�1��`&w�����(�A\jXsH��!{�(���}�j�A=���0����O{=�~(�{ZN9��{qn��B;�Ij�
K����	Lp� �o!��D��>��� ��N!M���C��ߨ�+�Q��]�p<��yB"�>��ϊ�(����5��Q�aNET�
p�Ǩ�(��>F�ܼ=7��3V&)���.$c�����R�.<CB��@e�Fkܼ���-`k C��1�T�e�q�M ��Ǿ��`��@���bTqތK���&b�>�:���nz�0�
���cx�����̌�(%M0�M*���\��7�~YWB�F[(Gu�K>v|>�S��T�񣅫�	�e�> uG5{�3zޤ�����䤅�H���b���+���g'��7���^>�'��Kb�k�OP��p�1bpb�l�h�ut�A� ���W���&l��=u-�ٙT.+����3���H�6��A�?����7j��a��O��)wH�����v���wH_�s�e�OP�!�=!1�|�T�+��R횒�y.o0�u�#<��9:
H�7�jހ+Z���e/���ũ]bd�����y��t�3�ވqR�y�5�/�)��gD���o �o��o;hy �K�=� /\��4*��<ؚ��=L�Y��=(7� O;@�\[;���@�����Y罭�r$����J�`@�0̺�K� ��9���>(�U?�!1kd8�[AJ�7WL*%X�X��hFp�~~08��}�oY��]y�u,�w�,�P�%��>��ޱW �ǸҬNI�ŠQZY@Smem6�aͦ��>��AӾB�N�8<	��ʂ�V��3��)6��׶�?#R�u�h5-h}O h�_���<^��/�����Nѓ �����=9����_*����i�Ǡ[�����k���^�q�B�z��IH�N�һ.����<��b.{0��Ye����%6;����i��6��'0m{P��L~��V��-'���߂�������I�J--|��9!qb�|`�� 7��6ٵIܽ��Ӥ_3�PB�E��cr};���B��{�w$}�M���rY�o�a#3�UE[)���䀗�t�΄R�ϱ�8'o'iě;��*v�_����+MwR��E��_(��+g�����-X�0� yr���\����{.��x*wt�����}�Ɠ��p~((�xi���ko���[�����S��4)��!�R���|������A���v���c��d�WXb#	P1�� �ԯ��vE���{fv����|K��DQgOh����y�_؁�y�R�E�VK�(�ԧ�J�1���9�w<��CEw�����D
܀V�߹���G�	��7�R�T�W��1����`"%;��2������8f����)�Wl�,V�,Z�ՇOS\���\����;1�
�����z�H֒�al� 򭐲_���H$%�ڮ�T�\���;����bK��`�� B暈��}��`�i�'e֩9#�f�с'���P�q�is�w�y{T�q��TDy�U�|MmajJ��Ѷg?�l�,��}{�w����B�}�:�j�Ԍ��!ץ6T*tʷ�Q������͝�Z�xM�.ׅ�y�~��zsHAU?�o����.g\�Z�V!�֨�p��i� v�'ײ��)���SoCu���9:��Lm=~A�uw�u�d��{��-Z�~���A�y8��¨�O��6Ew��z|у��Xll���g��F~P�oz�۲����b-�x1B��
(eޥ�;oM$�uvv��N_�/��u�	�����.uG�@n=k�ށ�����#��Ϸ���|8Y���Lv@����bgx�ǈ��.�G�.J��gEG�,��#eLz֣��k��!�K�vne��M���z�=�+�G�
hϯ�w��*�Y��9�
q���M����CM����g�W�w����2Þ���)�
Z�@�>nWo=�&����W����	, �'6�γ�f����W�9u�k?��v*�����������/k:��G��K4�JRv	k��W�oAd޾�i1惰�T��:�W��pݔ���F�����;�k<�C=�����-�N��w�Ue����c^sj&+���'i�xQ[j�l� GWZ�A�!�t�`y��K�5�-\�o O���`���@����5��t S3��/�G�In�-��.4>����[tJc������`ס
>]����/����� ߩ���o���k��ϩD�����K�OQ���K��9h8G�|!
�ݹE!���A�ݼ�/�p_㫸��|���*��-ᕺ�/�?���l���<���7@4ε���ޮ������$8	�矙��?O�����y���$��.��9����mJ�jRF�X�<K��ug��V)�[�9@��mFBM�f1���T�Yҝ�s]�^�m�:��6��6�W�#�|��&?�m��d��T��N���fU��rIu�\'dW뾆�WGvZ�g[S+� �)�I�O7^W�};��\���ڭ"K�Y����=�9�I:`��mEv�3��VͻI=I{���6�+��=J�덫�EԎ�,{��'���� m�����?���0�2��{�sA�&��{��oB�P�(ݙ�"��Vŏ=�/�D�U��������� � �b�����cf��d�fc#'��i��F[Bq/�8�-��3��w�QØ�&CǱqF��c�fOO�K}�Ț��V��<����i/o����:���#�>��+���1�xHf� fWܦ^���B�(h�;I[= ��Ag:�*�v�`^j�٪I!f�o���C-s	���[k��|j�,nP8���u}���ǋ)݂Aݗ�m�|����rv�6�G]�(�*Stv�nl_R,/%o@#L�i����A~l6w��V�����}�w�Lx]�&�;�s�A#�MWz"節?W4|��<v}q�կ=��sР���<AY�Jx1g���	h��12��pP�n�u�>$��4��pjG0���K��{�,�w�����R`f�W��A����mom�"D�'0�h>B��A�H/����^�ꀗ���
��**^�5�⼘���DwC���_�ˈ�!��7h�<�(���їV��ѽ���8\�f��JK�޷����g!���y$�-0�O��w�zǇ}@�
b׌/%Ń��8G��x`�W)Il��ՄLG�/�[`��pŁk2t]0�U�*��v�!	�U�U�@8'M=^�(�}~t�]7��_w���`a��b�@�Wz�͞áu{ �Z���h.�� �?��]���oq}f�K&��I]�m�/[ �S;ሧ+WmU�.|���������7g�b͵zR/�MVs ~3:S2���{u�u�$�o�q�t~p� �ӷ"��D�˙/�I-mqʹr���%�Kr`VՔƕ��=��j�xϋ�!;K�;,��������z���F� g�|���T��>	7�ؚA�A�������|�o�'9P���͑��������h^{��D�<mna	R�8�I�I��v��.|4[Y�ѿ�W����Rq
�Ĉ�����{���=�V/��]Y&WAuK�O����k�H���5<�v��{^���@"Ѻ�i�)�(�<���WKC_W�!߻�|��Ǆ�!?�+�hp(��N��1L��b���'/w6F��.��z�nN>�c�DߐR�sn%�`f;��8s�w�c�A\e>�wE�T���J��jSa���͘�:
c�#i�=���݅ �JV�S�l�糘���ͅ7$�_(����Xj�Z�i����@�+
���%f��	�]LJ�X��B��8s��wH�ǝ�;E
�e����թ	f��Y��"��mN��*�,1�[�ت�5`u;�!���R���oqIe+F��ry�Y˞� Hq���������֤�݃hAu�����ހu�&]�Ke�*t�9vs����ā�ͦ���1\SD67�K��;��ѕJ0�53,�5��Z6���7MV2|��&��k�q.�7�f�DAٯ5 ������E�w�[qQ��^$�k�Pׄ�l��W�.m/
�����[M�z`a�������f��Øk��wLf��1��粐&��T���ou��_��7����z�� |�""�O� 
ڰS����v63�[�!�L���-���VQ�%p}H�_��B��i�ƘA?�:����&�?�;+E%e!c0�@2J��NÝ���Wa ��������|�L.���q�%����ދ!����s������ĖnZ���F妘[�͆���tg��V�z��Ns���0���n��n��[F5��?�k{��w`�c0VyP��.ֺ���fpՊ?%}`�Br0�L1|����ݟ���[�^�Nuk���.�Ʀ0@��
zh���m}'9r��c����@��!����ͼ�>MN�X.�������e�8�n8ǭ>Z����%�f��a)�Su��H���S�:-pr�*A�'&�6�r,ÞՖ36��@��%�:K��������I$�;��ZX狂��ފ���a�!�,���k��EH7���������k�W+b���BMf��Ϭ�Xdp��~t��f�`�X�]����4=M��ᗹ�ޏ<<Tv�����z�{�x�{x3 ڗ�8�P��O�~���z����E�\nn	%�YR"��5��"�.���e��F�ma�+�����������k[e��+�2��J�ꦘ���B��4D�(��m�xЇȄ�>c�V�)���ˤJ/Y��`_�e~���t����6��ÃC��.�8�($⩙��Ӟ-�E��;m{�MW�: Mx����a�A�����a��6=��RB�'��z�ft11�_�]Eb���
����Z3!��B�B�K�ކ$(n\"5���:��x�G.Ɵ�`9+�Yi���&fh�*U"�����VF��z� M:j'���%�`���3�B��i���w䶶&P
I�J���[w�Qt���T ��^%K�T?�)��_�%�Zu��Z��X��6�h���k�&�{��Ȥ���ėX�mO��Z s�Lx���Q��ݞ|I���|�����H:���\ϟ����PhO���v�C�\6l��ᶼ�����˶�����1-��: 8�!���th�{�p�������<;�0�:E@���gǩO�-(��("%�S�q�����425~�9Qr��O� `� �֓�k�գ�y��+������g/s�{�!�ۭ\K���G�i��C���U�X�5&���������Te��|6CC�ݵuO�}�׿�|#�we+@���	�e?� ��5ݖqD�%;Xڛow���2!G�(b��)����<d��t��퓐��`�8���Q���0X~Y�� ,�Z���%��T`�e�:�������B�#�z�����>���:
�H�y���+w�)�So��E)����
sTL��͒X���}K�T7�9����_Ր��V�����X��%�8i��/�E��ں=�!q2K���b=D�۴.��a�A"CI���h3���E`�s��%��ۄ�ض�m��>)�LO�H}E?g��1x�@�	G�X�� ?�iҡ�����g���_ ��v�0���&4�Q _�+�/=�2���aR���Ue�`.Bj0��_��`W1 �5��<Q�F���O��ټ�US�/�C�n� �w@�8���ڳX#���h���PT�PRԂ�E��z#���v�gu��;�`�x��L"3 ��,xw؀:MJ��-������G送�'�욹=������u/�9]�P� 
�6�}Fz�����4Bf+���a��Ǚ�~��㞟4��4b���(+@������K0̕x�c ��ծ9���Z��1is�[ܪFi$�I=y�hEv���^��1�+�B�K6�1�v�{��>��K������C4HIӱ�ZkBjd��B�	��<.J*z�֮ϗ��@!t��^�wB� !���Ӥ�����&����p���c.�3�g ��&G�JcNb� ���񌍺ѨT^ҧ�;%J%�-y����3���v�i68�öo܃IY+��8�W9	��Ic:�K�B+�R�{����þ���Cxz��a��I�m�#�#�U��0x��n��(J��QO�u'*��!PK�a,����rm�?7�|t*-'��!h���[RZ���M�%䚸�&������p���8mW��g��e���Ez@n.<�(��2�f�]�G��t�����퍐��9�"�?�?����`
==�A�T������6��3�tq���^a2 w^�`K��h�����[�����ִo�",Y���wj0�ʤ�1�S7k�@N�PB2����w��7��!.�
K���;셉H꣼�"H��K�;�st�Ğ]��K�g�GǾ�E�D����	�� 8P"W��ٙ����	�Ϫ��_���B�a^�nl1j��-beY��t���H�	D�|`�5�.h�b��@�����}�j�x����<��"-=���(�nL!��>�V�m����i�5�tN46*~�2��.;�x�l\�l`�k�+6�X�Du��"(Xbc91gJL�?MR�V{�
pK��O��ޢ|>�ó�5��'p�C����
�xt|�����J`�T
b&��(�?U�B���f@��;�h�#���$!٫�Tٹ��3���b� \}���ʞ�ZB���'opn!��SPt]�SڬH2Y`2?i��g����/��,_�M�ֽ�������*�������$�Z��!�LQ%��'���>/��D�T��|�����q��KݤoDߋSgv�xO��u�n-<�K/4�ѱ����䃟�����s{s��!e����`a��3�W�^{3to5g 
�W�4��g���-m��"}�Z�/�x�/�S>��UC�3*0��aV��5\ɞxS�IzZX����@�1a�z}���qU�Ge��"��U]��z�n��c�B4f��n�֥��,�DNt���]U��P��]u��y�P�t�L�aq�}���a�7�|���'4�g�j�\�d[I�uY����w�!Q-�z����6L��� �+�~B�����7�Vh�M�|��&�|TJ+�٣�e��O��6���Gy��h��[JZ銂t|��j��]&�#��*MSOᤢ:��F�͏?�V7�:Y�(Ѵp ���k�g����^�������\m��×8�l��������n׵M�
�|mM���n}�����ᚧ ꘴a?)��ў+�K�5Z�K�UA���u��W;]�i��e�2�L��m�Lrp�N�ܮ5�;F��D�
r_��6���m��L���ӛt�߅�_��1���K�a�-��`�	 �q��/35zk�%�S�IଧR+^l4 ��N�9 "|�/=��� �ܬY+�/�Y+u���'��D:�o �um=:��@|}��#ff�¡8�����Dq��d�{6{��
��U���gO�"��O���Q��/�N->�^�\��͆N٢�Y�i [��%�#�={'z���V-��K� 4>پ�)���g�PѥV���ͷ���;��i��Tu��O�QO�L�]��.$�;$=��i��xӶ�u^]:�U{7P�%���8�&���L�MM����f�e�$���܎�-Ӗ����І�^�;�2X_���_ȝ�����r�h����R��x�B0�4����:�ہ���7����J����ȱ��K�0/�]�{Ig�	~#��U[���O;j����!d�I�>,ޘX��$��ל�~��B&������U����w�.�;P�ﻺu�̒_9�`q^�!q��+�W�sxB�R��h�-�F��o�6)���Y~D�� �[-Q|%�z�Ԕ7uf��0��W��U���Gw���va^�'��byeC�����s��@����V�� �=Ȩ�C����_�Ƕ>xL7��2 ��o��k#w�|�(�t�5qD�旉�0�/LSf	e���;�l��jHC���v�5T�y��@�Z����X�V�=^��~?�����x�C���g�v�F>�d�����;r���œ�T_:]v��7ӑi�7'�&��*����K��*��D3��_S@��З��͸� wiGO�yϿ���1���/J<�b��/�Y'���<�t��K-t���Ao��?��&5�Sl��qhV�,k9����������+�F�Q/�� �+;P��!X��:�k��?�_��������N�K�+R���v�
[]4k5�]��G��_C������M
�$��Z����^%Y�1�\h$�D&v�"��u�8U�����_�o8�N��,�0--��F��ϋ���*'�ޏ�Y�Y���u ��Qgf���2.��N+������fP7��yYՎ�D1�#4T񱗠��뽯�%��:4A���[�;IE��L�olQ06ya�����*_1��h�q�[oWW�O5�U�X�7��X�_�M�W��Ҁ�*�BQo2Z��ī|�TS(o2<���t�~p ��\��V�l�X&��xPk{8�E9"�؈E�#3����;Q>�k����,֙�,f�W٣� ����i�3�������Lø\���R����w�ĭ�U��[������m�ѧ"OSJ��h21M��kUop�����'C-�=#��޲�����0sv�K��+�Ĭ��A��l�6ЛԜ��B(aJ�9էg�O*J��(�N<� �Ur B?O ȁ�����-]�9`�-�%���m�lwR��^Q��e0�]�SQ�P@Wg����Z����������x�8���a�_Ո=����o��>�_ā\�^rx�J~ruQ��ƕ�ja��9F`��b��崪�C�9����_
GIT�F�ʱL�E(^e%S�$꩝ͭ�@]���Z=�Ew�c�BBɓ��,��G��i̐���T��Fl��'=?G���ۙ�5{<C�n�oM| �S7Y�x����<�;z�C�Ŭ��$5-�4��*&���P܇|r�!�ԗ� �׈����]�^f���澇�p\T���=ضK^TR�Yk�XW	��̷Y6�j�S4hr�O B>�h K3?z���7\����7��/&�By����i�b@�K���=��WXA�|k=�'՗DzeFF���L��Yy��~R�|��_ -!{9�]��K���_�8*2��]�y��_���h	����9l� ��o�Ț��ݗ������L���~+);7Ru����4}���6tZ��sԙ���|��S;�K(�9o�'���4[7A�J�����S�O��+���j24���^V�hY��|�I���*��x�:���C���m]�֍9h������t��-T�}�3�ʃ���� ��:�m���G��m_�6�o���y�����Z�2��}9�i�I��x�)�1��'���/G7���Xl0��ǯ7��_��L'W�?d��ܒ�)3L���������ӭ�DT�#�|��Cs�4�[,q�4��ȳ#@k\n2愊��, ���D�h.�rK�:�B�T�^��㐿���ً��]@6�s�#d�zǨ�l2H�Ro�Cq�)����n�D0�Z�P�f�����U�����c@�X�9��@�*���'u���R
�3��-����M��:[R���4�!fN�+��M����_��H?���rݒ�U�ɢw^�`�A`HB,g���� �*Iᢔ-o�(w�/Z	�1�'�x�:�3��v��!��5o mI����i����4�^�/W7eE�4A:x��{_���+�n)��f�3��.uViR�r,�ꁤ�Y)������V���#f`��݋<Ĭ�Fr(;:h+ ejTB¤��u�d"�p�c:�w;���Ar��hF�� ���RY�<�V��l������tx� A�Q��#�T�y�/J�;zI7e�j�V�kC�/�OE� �oq��Aq���^N�,J��Q�,'y���4z ��"�;���ֱԉ/� ����o��%ɒ���0�}>���(����{�#z��h�h��]x���!U�{�]�	�T:S������Y�̻f�Z3X�;D�<(e}�r�����_��s��E� ��,��̃^����Ǘ	���xOB��-��!�9�B���ԑ�ר����iW� 4�Xªߪ��h~,i`h�;3M>8m�2d[Q�l��BO��w�&�.�N�N�Dm)ˤR��b��>o�=�[�����b@(:!��M]$�;xx�mv���z�Mw0�������:��I˶����}���JI�
��1��{��Q8����r?���J��HU�j����A:_�'���4w��ُX�uLBIB�T�\�Ş��ϡNz������#&�
�Hԡ�̲�)�s�v[+[++QZC �����B��"�:��[�N� ��ˑrR�cyk%�D����̝����"���X�׆�ɑ2S����8��������'0U~6l�[zgȄ��X���(�����(*[�i��*��M�1�>.2�g{[�~iі�� �53`��nU�^���6F��VJ�q:�7apOKUx��,e6d���PXL*��b�z+OX�%(�x:��"��[�	����M)����/�� �V�g�8�����q�p/�c �o8�J%h�j �����o9��j��e7�Z��w��l��4��-�ݧ���;9��a;(�@)�����yMCxC����'.H�Ev��Q�J�±鄸�R����@�CjLpő��c��[�~�(K���)�4�K�1E	K{wr}-��J���S��!���E���䱍^����������3��H0���VJ���_`c�a)d�T�R��콽��x�����&e���`"/�c��:|��, 8���b��w�;$A�������*Dд�g�ኀ�G),���0�t4Z,b�*��.I[� ���mFg(��j!c55�6}� 0w�exp���cp{��;�Ձ�S-y��������|��O�|��[v��ݗ�����ٽ�\����Խp�p��Ra�m�4��x�����uc�sX���o�Iģ[=S��n-��ʊ�h�8����.�|���0��[{$�`9|_���=���ׇ��,�b�a�
��'N��\��ֻ\��VX�U;����pi�5L̴���j�3����=5� s	��e/'Ε�%X��y��m� ��l�l鬨Hu�U�{W6���8�l��۟�w����q�D��mۡ�g�_{��}��l�c�c��`������*=ʝP���ъe����Oڰמ�z��V�r�?ͯEk�>j%���ܨo6?ܚ(O�"���b�!�_;�qP�=�K��.�{lMIS����B������`�hy���j�a
85�T���v�Ϊ�rt���簐����BCk�2wG�����e���{	�-�a�1�����e����G�?���;&� k��š���]�jڍ�3L%-.W�(<ǒ�|r��ܨW����;��d@�rѫ~�M���W3B��-�կo��=��	C��F��J�kk	tȚYW|�G!%�������]�ɟ�C�\9aʠ�l�s����JTm��G�[���"
d�[:?��C��B[XyOșjDJ�M��ؖU�2�*�!����ϙ�m�|�d"1����!Q�!k2�$$Y�owL'[ ����ŧ`XP������Q�?�d���_�g@B���=�X�lF��f׵w�q�W�(=G�� !�d�J2��
}��s��!��������rM�`[�_���r�έ�L��"���n�n� ,�z�X�%�$�F�58��N1+ ���o�Evq��Ӱ�X�@�U�w5��UǍ�z*�W�C'5�[�D����}S������]�=���XWN�I��2�>'fv�̇����W�כH��A�ߕw�9��⏞�Y�����/v�%��EnT������!���(�BP��S���HҍAZ-�����d�����J��u �w=���P�[���Xu��5e��&,/�[�O>�,�SO�! ��4�]�p`x��rp#F�}�y���L��4r�Ktj����)��U�I�y��$�d��w��E�+����e���~>@��x ������a��uǱԔ��~�l��w�0����F אI�����$&+�vN����w#p���{�v;���۹����}V�L�;~��-$]���BǮ�5%|v���Ξ���]_=��?dֿD�����0tʹ/.l�/&+���}[�q�`.�J0L�G�4_��k�l��k>����;���o�$���
:�$�ǧ���k'!sa�Q�V�>$zp���d����DeomA�8�'������F���N3����̐3R�c���7|���Ɯ��wv��#���9s���A����`��Gމ���&�+`)�27ko݉h���%=�Qp][}�<�z˼���濡D�y�qy�3 W��~w7��~q0m�Z�&��L宆vqtF_<q�M)�˴ܾ{VypOx�ҭe_*���Y�Pk*d�Ȼ�C�{�����"�4ծ�b��6��s� �gΏLf�Ē��������Y?��`��馿[������1>����C�%�C�x�ӽ.�a�t*"���t�����y�A���d��Q4r���l�)X'F^q�)�\�Ǭs�LTT���ԩ�Em�ڐ���z1�o	��f;Lqm�E�.���<1`֥76= �!8��s =�bY�ڴ����g�D�,;""�6��4�����C��z�F���k�9���\�`ܛY*y�,aw�[�K%��y���u���q|�m~L$Av��*�ܧ}G�ύ"�X�>!�����W4[��xL��ub�B-����%6᮷@�����Q��G��OO���!�ę�X�l�S��.(z�9�����q��Lp�%�V=J������B��-M2y�|�k�(�1�O�e�m�2��$���A�҉X�+���b}@�f>� EKz#7�v��| rh��M��"��0�g�'{���X����l�庫t���P�㟾�4Y�����|����@��w�)�ח��vݱĠ{��4�4�lNS.���Ԧ�a�;NCs/|9���������1�Y��|z��`/��2}�����	�m��H�$�!|{���	 �lÂ˺Yt�"�&��M��qP?�gr2C&jիA)L����2$�rn�A���j�3F�G��9U�� ?Wx��P)�F�+'�p5�����?�m��h�$�K����XS��shqXe�[5�6vcҬ�r����ږM��k��~�*�@���YYq�닾 �Q��G0�&�'9��m��J���)�k�l�m��g{;���@".��5N6-�}�Oi�@v�iE�-��!�<O�4������1ˡ�-*��c���|��c,��^��!�X{S��ior�6����e��l"5��w�� �b5���p�L�f��`�O^Y_x�g�jЙ������ۋ���"��wfn����HFV}��AapeJ�a:΁��6������A�ܴ���c':�a�#��������PakȤS)j4�Ю������҆3|� K�fju��T�\��2��N�����������f�����"�OW�G�W����a���zѨ��Q�4�^�3�	��a�n��A�mm�iD�u E�!��z�|ri�r`v
�?{Xy;^����/��b�eb�O��ȹ'�w�ז��$���_9}�U�#|:>���!��� w��|n�2\�E����1��7�n��#m@"<@"ȉ8�'�/'����U ��+��������;�P��#�R�}��-(��+�����*�H����I���ݞ
5 
n�e�붯}IL&XV,3�y2�㼫�4�Z��#���#_�f>��;6�z�.�,�^+m��z��7ٌ&���0��yk�=���(�����؁gC��d���U�_�E�O @q�DӲ]��X_�� ؠ-2����#��4Ķ�"?���\bl��/��"���s����Mg�'�|��{�����:� �7l?_%�O�!}d�n�!�!!�	��4߾�,�6�E�M\g	�D5�I�1�������-�e71*%�������8R�� ?%�3T��|�Y{f�bhG"��Iۤu&������o���s����1�Yl�4^."E��WQ 	]�@UI(��Zq��K��t(�]�?��[ ������8r�+��g/�9%"Z'�϶O�~��:dZ�!�Ds=��靆��\����y��<��(�(�����fd}�b�����d�sQ/�2�j֔w���=���kn�1yt�p��)��N�\u�ABU�c�0]�CVi��U	�����ݩE����B���!MS�^ [�$�u(]_n8�����x��+��1Y�?�m�ҕ����k�z�p�5�L�c���w�����uJS1T�����D ��q��L{������ТQt]��Q�2�ɗ����4��F����料3�:�%��Rg�n%}�(�#	�u#ߍ�������j��O`�.�'� �	��RX�4��-��d��I�##�[���VSv��n�J������`�ik ��hL)kJ^�����d��=i�84��b�O��ǀv��б�P~bG����dǙ��Sg��fD��mZ�jXz��h�S�7�T��� ��ͼ�QY��WL<���V�&�²�a��t	.�e9�DѺ4�:07�j��w�q�o��l
ߐ��=����7���g��K���nW@R4ͨ��7R�ͻ�����:s�^-.K'n %�!�]3�ɣ�ߊ�q�4�3���|�~?�����R%��o�����R�����?.�(}�ڢ����m�4w����zۏH��B������5~�c�߻y d�cK6Ba_L�7^�n-l�����`{��}���1G����-r�~���Oܚ���S

��cF�X�H�E]�v�3و���#ː#y�A����@�s�ډ�JpJ��B��L5t�q��w�MK$*&��Ҋ�`�rփ��V�d����*z
���> M��&��߼�A=y�I�>�ewuL�I�Q�16��D8����Cd��r���b4�J�5�h�Ͽ�_��e��a���x� �Z�J��,�D��0��A����&z��=�պ=�kށ���:�Z�C��~!{��Ao�}���kz�q6�ٳ��88Y)I$t�I�?=7�X� �U�tz��p�
5�1�=�x|��k�k ��㓽s�L��{��E��뮸�]�iE�`@@� .""�  ŀ Y`$�₂��U�̐$QP� HΒs򯪻q��u=o��?�:5]U���>�9�ӥi�Gk�"�?�[��ց����)�]�����a�;� r�����i���"�����޴�Xl���`��m�@}�(x�%6�2�����c�����F�¤M���M?�M�Bp�	���r���� ������V���;G��-�5��l�u�J+kPڵ'X�uGFIjߎp�XZ�T�TAlf�[����1�j�&'*s #����܊d9���m82e����b�س��*� r�8�1�),��FӾ6�e,��w���1;?�-a�:{,���e�C_�[���C�/��Ye�����i�O�;�og����p�t��(,gV7�!ԭJ��s6���.�0������y�M�h�!�}��|MOt�LGbï��c���j~��1�ĳX�����z�}��Т���x�aB5��
F�;�~���S�����/�R�BL�+Ua��^W�NlѼ"B&��Z {*/�\��M�M·;�9� �v�V��q$R �K-J�o1�� ��v�۶K	���z�����Ά!�G�+ف��y�_���8�����o�����*X�|&þ��جΥ��}+�h�ZJ~!�xڄ)�-�/��:
���)�!`1{�u9�٧z!zCX[��c��V�R��x�ڰd���U�P����&���ry�᎝�@�A�"��hf���9��.���Y/���`����$�Juگ�/a�d ٻ�w^t�	�|��&vH�S��A�޻AldE��_���q�0|��|߻n@���M�ⵯ�xJ��⁂���r�o�X�)H���F>���8hMt&�ӿ���ۡC�V*��m_�[�d�K�R���6�;/���Z���י�Cl�����FS)�ZB#'�\�ָ�f׏��1� �w<k�=��q�(�"e��|�X>�	����O���D�T���툴�.���D�������2�j#�@��o��!B��z��N�ހ�˥�,A�)@4����s�/�X��*ܹ£K�p�b�R�,����TJV0'�x�Hk�ol�w�qY��
`%�)�";��e��\�ǌaK�
�׼G��/Q{��L)g�.�u��~.��o���#������&�iTZ'=�=�x$��$�v�m�(ǰ� FM��s`|��q2�A��m�M����HM���bam�dk��|��[�%v[ß���Q����o%�컗�,M��c�;(�l�M�MG�d̪O�;�ZQ�G7m-�l���K�c��)�>k�Z�����)w@>�����=�	��{`ѭ�&è�Kzo]�k��|-�e%\g}��}̡Je�^R,�M��,R_�=&�r���ĝ�����/�"��Q�U�6c�4x�©�팿A�����C���A��M����+�x%��6ੲ�hn�F\��y�O��b?g��N�a>ݲ�{E���~|�������CL�&�4(-H�l��_�M[Y86p�����:�Jb�5�a�p�-}m�nL�{0�v9���_�jf���6���-R>9b���>w��O3�O���@#��,��3e#L����l���ZP 8ht��QȈ�I�7@����ҕ�A~�A��J����,���Kej���PJhilk�����Wt]~L�l@�1��e/����b@j�J�L�N��8���S�)�Xk ~�� 
�W����cX�tyG�������dR����)x�œ���V�<��&�E+�M�@������S��Д�m�ࠆ#f����\���C��7U ��2XJX2�1�]�섽�<�X��XJ�������H�ϥ�pཱྀ�O��уR^Kԁ*?�<������ �xi��!�q����������&���/5).�x�O9c��~�]&0]��J�o�#�����{Fd��J��Oc'�@D�j� �F��{<�.ƙ�X���E8QE��T^j����m[��,�ZQ L+�UK��A�X�>˒E�Ya�Z�ne��
aw��%��YI��2�CT���\�Or!s�����ۍ�@�{l+'��\����,zC:��z&q��?R�қ������(/���XTfZ�N|����%�xU	(u��-h?/;��� ��c2�!rM��~����Lx����3�=��������6���ͦP�� ��(�]��jbܙ�݆0̧(�E�&��[�*���y�����aK#'(h'z\�73�0cs��G`0t��Y:��S��~CL$,��RȔ�^����G&��z�Ԕ'nVZ2��niT��U�v��&��*� �#O=!�o����c������׎
� M�e/T�tI�n�N=��:�~�Y'�����}��c'���(O5Y�;��D"kk�����S9[q�
?3Z�H����7j�b��}�e�7��#S�R���K�7����և�g�C��r��
 ���������`W��9��Pҁ���bsk¹��-�lRx�cv��#��L�����OY��æ/����l:Qmz뚓��B�o]j��U�6+zq��|��W�<0<��m��$�3R����	��쐢��?���ڷB��j��9 ?� �!"]Ʌ�Cn��p��%��e�KBAs��cD����nc���� ̐�	;��ݝ�j�H�Ch��@%���J�l� &�H�ܴ����i�gj!r���J�
Z��2s�[�N-B)����|�e�N.�w_	�%�+Ͽ`q�I�Z�e��_`�J���D�^}���ȯ��nkPY�nV��m�d>V��n�n36�����N.�=@M�����ޘFl:�&�BX
p^�>"ŠN����	���L�^�R�Y��<@^��H���oT����6K|�=�xʹ��l	F:�1~���",�G�g+��ȝ�0��=�����k#�U�T'��^��s:Ժ���U�� �N�T#ʚ{9��&RC�������Î�Y ���[#z�Zb6���[�5�����co���w�6<�`���uE�i���`RL��	���}�%�ݺ���� ����ODB�;��[��ͪ�����Kh�h�ws!�t�ZK�_�p��4GՓ�b&�&$�L1�rB]��T��f�{a}R	Y��6�n��1��A��gw�y�A��?!Ƽ~Z?�c�Ύ$�Uկ�����(@E��YAE��,�j>�[���g��KQ�%#�Q��_�a�I|~R4�0#�M�~?�F�.w�.�?�F9yU�A�y�%Vxze�+oY8/�y* ��n��G��;v�܍A����X���L�漜:T(4"�k��o�\���$w�~��2�}��|�M=���| �u��Μ�Y&y��VD�&��W�����O*c=y����{��Q���$��:ӐM,��8��k�m��h/e|���n�K�*b8e����-:L_qAE�5�4,��j��K�7�N�Q���m���H{��P�M���?�v"}��f*�Hl�Mϥ)����P�P��3�7�pB��:�,�#�E^g+6[jϸ�}���]�|v������/؟�<�T�����uK�x:&>�٣��YLP��R���eS�Y�`���A�X��L�jn����4�r�!\B����A�Z�m��,G}�k#�4c�f�i>�E#��W,3O	�Su����I��o��@�i���z.�uO�r�C�QG���0c��9🭒.\�����5�UG���ɨ1Gޗ<u�g4�@K]��<Z,-�eW��/�-���ǫI$��c��J�<�6�O0�nzq��_����T�U��ѓ9�Մ�n�O{�e���}�A�����Zb����ǡ����H�n�p�v7�=�~�ȧ�ϴp�%ԭd�z8x�E<w���_CJ��Õ�W]|͞�}�l��������>!�n�Jw�L3��n�]C�gʍe�W�,$��C8q��x�`=��ĔB~��(lX�2�����}������>�߇�������}������߇w��&Rnh͔n�_��IV�{��Kg��b���O��U�wM�7fM��ow\�tڞN�(1��V�r��Jz<Z�����k��+��k0��a,�A4k]��&G�� Nk�>{t�C�V:�gyA3�#}ETv����f����ؽV�}o���^J�RS=4����[̽�7�3>veJp�S�TM�t�.8[����f�A�2I�q�н�IU�2�+7W��%�ɌoVʳ,��//t^I��6�6?�>#������4���6�ʧ���?�V����L���cr�-�}iO/]�L��ط�����<|=j���S��RB�=V�`�����9wbO)���a����o��������$��G�0�J��O���g�v��y������ �, ��\;$�C\"U���rj�	�,N�?`'�5f3,��.şX������R�7���^�;�Bh[�{�S�ŏ�p����y�^���zU���_��8[��~�m�m���Z.b��cǿjpGr'Iڼ��h���0X.7�Z}��fn����ޝ4�J\|j�"�#*az�+9�\Ò�y��vM�&�ZW�j�l_,p	�Noۦ��oyf;���t�Һ����N�^��0��_bʵ������il�>Z\t�'���h��ө.�tO�z%�H�
p�d.�B�z]K��#Yo�ɩr�h�ҎBKJd
�Q���e�,M��=�[�3,���F��ќ�g����"�x0��위_��^�O+�7oڌY;A�^��F%#wv��.�`�ǹ|�7��v� 1�Gu5͚�Ф�}��2K�J����"u�PO���#�Lv ;�"S0n<a�Ԗ���Xӹ{��P�d]���kp�MaW��,�Ľ�����u��[(��Mر�7D�I>K_�y&/���c�j�q+�OF���Iuqj^��A_��5�lXa�CZ�dh[݂n�	�`�5�$��L=���H��/-22�K����+Nݶx����8_�5�.r��=��nh�_1�6~�N���w�P3��*�?��p�2�8�a�#wMU���m�L��p*�mwﬠ0�0[��yib��a�j���4��8��L��v4�4�^���X��m5=�$t��13�^�~�o07��7�k�}���y��]���l�,Z�u&�o6�&ee����>ʒՊ��V����r.�Cm��_g�{%F�g���32l��u[���'������C���j\���%��X���3lZ/�n^�uIzhV#�\����*Bcm;�4ܸ��Z_|6���,�|�䎷�)��`"נoIQ�b��6ȿU�1�C�ں���~'��BЯ; ƙ���[��9�%�a���ř1�L���_���}i���18v�_�e�\-Y*_<�;���oj��a���r��ݕ^�e�M���I��n��q�:�#l�>,5�W Y8��挡Q�9�>��_����u�Ƹܻ����q���sM�$�2|�.����Q���w�bNR��7�Du�Ǽ��z?Z�l�(ꕵ2���lޔ!<���R�H@l�)WW{��	|m��y��FZA�dn�K��pi�<h
3>��v�������+ղ�}ߡ�T����c�ϑ�֐S(nmVHjN)ƫ����b��m��vJT2+� /��&�k�8��7)S��[�\�a���4�[�����lm]l��6�<�zr�X�x����x�m��Ya��Y���QMN7�V��s�t gmHM�@�xJz4��m��G#4�����HC��FG����ik_=z��������낦[<�uZ;WÉ�&�96��H�TZ�t2�j�m�)�� �����}�#�"�����^?�=�̍�ʍ��[�qi�8o�r�·�P��w9�	k���Ԍ �Ѹ4|]`k�lu��ۋ����%f��YSL�y��;ȑn�q9}=������1��}��� �Uk���q��-���)��<;�����/6�'�����h�gId�۝,�_����Tb}��&�]^uC&�4�����©Ǒ&7�c�����9��V1��חT�tN���c� >�й��&?ߨZ��)���G�nd�,�����'���/z��Rh~��R��M��������o���	�նj�qF�MRՑ���Z��vi2�Wejx�*������ :�{���=E��[�ήܚ��'}�D���Ԙ6;�L33̽��1Wh�څ�ݶ|���\�`^n����!e{h�Z@"�'!B��H�B�C�0����I�cT׌cъx�{l�k�
R�<��sP� pj�w|ݧo��$=�_TTy��c06�.k�%��G�Ͳ����\?�H��,:|���9[59��/�5�w7����)oSeL�פ޸fK�c�6wߟ l�a�j��V����?�a�p�9��Sd���R��׌R� �j3�0�ܙ�/i:�L�� /�l�X�:�h�ɇG��9������t�믿�Z�L��-��c�[U��}�<1�G�<����\-ێ= �-�s��QI�a2d](G����7����N���M�rJ�g��� J�ހ��4#n4d�H)�m�q�����A�D<�s! HB��L_�hӉ&!~z&�TԍE�lq^󣒓��΍74%;R�Ǡ�k6t��gMέ��k?��a�� �R��SMVX�ä�د��f�!��b��B�֑��Iʛ4�xf��)��������[᫦%��[���H�@5��S9x"���x�uk��7�D;ܼ�S�u�����$�&���������j!�.�@q�(�Mp	m1=� �A�m��W��^0�W�m��&�1m<�;�+��/��˄�] �;�������H��4ܑ���y`wN�/J��yyf~�[/(2U�Q���~��[j��ЉOx�l�ι�ݷgj���/�(�I~)tnq��w��y�Rf,���İ`���5���ݘ��uN�"�Ó�u�L��L��r�w;&G]��5}�Ѝ��Hl�0l�O���_,���H�T�r��S�7A���͏W��ރ�V˝�_fb�uhx�!���*,���D�Fɘ̤���X�9Ob�O�fY�y_��?/�h}3�*�r�=�8��J��^�_ev��͘���y�u��?���v�@O�|�p��Ə�\M������:�m�-�W7I�6��`l\T�n�:�4�rWx���P�Xl;*�Ĭ(�����=�����LlK+������� j��ݩ��7�-]}@��h����+gx�2JڍS�P��4��:o�ju�oB��d�aoF�N�n��V���ߦ�>�l�=�^�W���3'�>�40�����K�U<��m�ٱL�s� �wӲ�WI�r�/,��ıT�[TA��5g9!�)v˳i����R��N�6p_ �'N�դ��x����ϔ��M��
se�]�^d�y�	�	��e����m��c�yw�����A#k�7IJ`��/�����k��^U���9)սyST�Y7��.��J�s"�.N���� Z�ĭl��"��&�A�^��ç�9����盜wv���ݚt� P6-M�s9�������r3���_���������m&ҙV�w�.����B��m����٧WV+m���M��!ϭ2\q��@�v�1�Ⴎ
�43s�O=��|Y�[�������+�g{��\Y�����
�v�+� >�8r@V5'�a@*��.��s�ƚz�����dZ��j�Tz���/�4��L�����(6���x	��5���Y��2�=����r������±�'�w�W�� y�ܼϻP&{�Z���l�U����� ~�EB�˩����fh8�+a+(��Q.����VJ���C����_I#��4�}?	����,A��ͅ��,=��ձ�t��2��Ykt�zCɶ�P�:��6�Y�9��`�jz��/f��Y�nFX��J�	��Ǔy�λ@(��$ ��)�����m���"�?PrKٷ�;||��9��-.��^��&B��$����s%�����'��V�ra���� �R�$�q�M�:�,:��;�b9�\K��i1R�������Qg�	a�Rj�ə\�K8[��o���n �X��ej|NCQ^N]Oy�Rx�[����7%���P����+)!�?�0�{GWI���$������e�eZ#��#���9��^��ƴ.q�1'����^�h��m���]����z?n��ޝ��-Ե����>S���)�m{�ȝ1}����	�,b������-Ԗ���c��__�ʘg5���Lf8\a9��6N���k_q�CzI��8�I���""�`pj�\+D_o�����������E̸2?�[���D��fC
��b*��+�<X .�\�5P�:���O�S���oj�T�r=0U��>�+���0�nEi#݆��h�_й��=����;9�)�QS9gr-�|.���u�ѳ�j݋��tu5t�i|��ƮhI%�I*L�s�s��g�9yb)`ƣ�����GA���r�A�`Ͳ���{��Z't����p���/�	_�6֧Yav$1�@�:��-�V�8v�M�1Չ��(P qn�]�?݀^{����1K	*h��`�����$�
���yS{�^��u�T!�5�S��UK��:��[R���ή~ �dL_)j���{�Bi��[q���?�8����R���?ٕ�CKb斃?똈�,iđ����s�)������k�l�a��=��"nN,]�eZ~#��C�!��F��p�1@#�M�r�����I���������BRϮ�j{DBE����e_���e����h�u2�P���Q��
��=��G�d����{5��!ݲ#���YݒR�Қ_�/�b_���?��#��&���
��RSWcb���F�G�����L����.[e�n\�/Y7�Z�?���=w-�u��~��RB���R��G�5�z�HW׬�:�ʥ'1���Iᖫ ��Mɏ���g��=!�Bl���~��OӍ�H�Փ��>�=�q	��ܿޘl�'�C2�֢d?�N�p�Ǔ�����4m�οhu����~�
j0�,F�)����'gt]A�<�B6��\eU�6�1v @�~�����v�:	�ϝ{��!\";��'p�ΥQ:kA�[�{��ʈD��������x`Zݛ�Ni!�-��50�Gx���N�y���_+����%�o[$3���P�����0��h��8�c�����f� ݖ8�74���`{��g�Ǉ��Z����6��g��C��Ԕ�ICkPx)iȬ���y����axK�d�	��{�M}1 ��Ĕ�\M�#s�_?�~ez��s��C,q�j���K�2�prR\�k��̹"|9��NZ@�PO�����!�?��:��?���ӂ5
i�HZ�{���c<j�Fx�WA���1�]�9��D�ˠ��jo+�u�^�������O�v�aZ�����P&�zAZ��l%=	���x =�Q_m�ǔ]%��ߖߦ�c<��Ah)��-7��M�>^�#�?���+E�W+��Y.�R�5����s�T��UyDUI��T�t5n��0)T]��
E����Q
�o�p���/S����� 1:�Y�\_#A��2��[�%�;K��@�p�����r��#TV?��!��������@J�q���?2'�U��:�L�J
N���a}�b�Jcc"B^�Q�/ܐF���+cި����{x<�XL�V��#!�I\�������0s����=����a�٢P����Ǐ`[�CO���,���FY�(�y��ۛk	�1F�ɑO�N����#Jv����+�3��m%s��#R��<�⚋9K����������U��ofq���߉?LK*���K�ϑxQ���D�h��L���ui��]�#-"��d^�e�~�D��۾I��b%�G��.�+8�ߪ�Ƌ�3bq��<܁�\�0imw�!"I�ÄI�0�u��.A����u���C�� ��Q�?8Q����$Bw��:p=K?�iW]@��mq�B��A����F3s}et-G�ú`T�g�l5��j@�tw�M��
�J?�yh��Y�rGF�:�]@pGC��Zo�,��0�,��a@b|�p8RwR��aT�W~o�>>��@�ړ����uS��J~��M8&w��+~��?�p�;�t�h,lT���t Ը*BOR����;�C�AY�����ʘ�X�[�nX��p�@2Zm��W�S�3�ͷM�. �Ø���	�s.��)��CZ)i�9���5�f�D���F"��c����ŋ��~.�Hs��2b�b�!͑�����l8�`=��+����*`^�#��o�.tz�����m�Lm<{-a����J�iKL���%���'�/�g�=jP�"��1��(�Y�lm8�E�罀�ĳ `"��tR�٦�{�b�It�\B�]m��߿[�q?�ǲܲ��z�W.�� ��,�\ind�%"��W(zAC�B���܎m�����¢�;H����V�h�������Ѷ}��'���c���m�&Ps�����Z��Ыj$o��Jb.��N˖a��zp':������ˋٞD��7���3b斜�+1��Æ6�0q�V/Ag�L-]ꔇ��^Hc�}u��mi�v�u?� ɕ0�nȻ0�(
^��*�m4Y��BPY2��bDЎH,B���RJ�5&�X�Nb:!�{_�|@�'�@Q����B
��Lb���Y)=�;Ψ����@��y��b���Ao��f�{��ό��	�k� �k��g����)j�YCƇ�h�'t���ɫ��\P�䤅�Z�精	�'s��$�&TF�Y��R؅����`*=��Z7<	?�ڟX��N�����.����G��%�7"��ǐCV�X��M�ʠ��(o��F����[ �3�#��t�7%�b� ���zAm])�;�;p�"eK�9�E�| �� [������K��>����ɟj:��5�X< ���F��r���b�ϕ)�A��0�q��J�&�#��
?L��Ϯ�㳮gl�|[t��2�������ϦY�ƛ�L�Bn�dV8�0�X�'�	w���V��F��a?u����K��	&�?;���!T�� &�CD	�겆�Oi��0�۲�D�� +W!�ҋ��v�D^��}W9�FRl�!����W��[VLv`lII�2�,^�V=�yJ�k�g2V���L��woF� .��+�ͪ�a���}v>�H�^�����=��?ƛSeB��w���GMZx~| �{�����D/��{�h��v�\�_�2'�{Т��oXu��j0��a� �#k-x����7��Q*�����(o�C,&%���n^H���,˄���>7�=1�;��$�J� )!����O\�G�C�xo�ƱcJ$�<uC�����VB�k�����S;�@�@����In�v9訟�<)�9}�޲r�g)�kG$�şX�;�j\\�6K����d|��я�'�8�4�peO�S��ߢ&q���I��O�G\ѝ���}�l��_p/��H�O��/�Z4��(�x�tn��`�'{<�/7��W�e�t�*4t"�D�����<�01:!��G
R�z>��ȼ�\x�h!�a
��u�K}�d���ƚ.����ܡ�}aK$$��~���L!��L�?��=V��x`���D��:,�+1�+D�Ê����I�<;��caN������(��7�Ԛ*��F���.�R@����D��,J\��2N�^$b��e�s��ɚ��K�ͽ8�;�p>Կ�ၩ��( �f���sm�+2WB���WC��W�4��)J�&�� �ڋu��.�c7�����0R��:�|d�L2������ �wm��}��E
7ܙ�#������������!�O��e,��b����CK��yc�`*b2�!z{�����@�6���/��m0��A����՗�y��Z^��Ⲣ��ϝ�\n�<r�)2q��^��)�a�5�V T�ܜ6�)�C�(��Mb!lw!?U�r	8?k�#��	�=����>��r��kU����Q�Z�g{Բ��[�x�]v=:�bD��ҹU<�����7���c�rɕ`��{ȜY�B�ܰ`N�_pHCs��&a�X���ER�0��i�P��A�sH� :m砵M��$2��W{�1�j�nz�?������������P;��ϪJ$���;����W`��Ӣ���Q���0���RƩ�R�$�\k&�;dr� �%�=l\+����&X�.$�F"P�s�*D)��}1����&�r��˩�9������	�����b�D�b���4�c-5"H���_�M�q�&
��k��7	�����~��Ab ޏ|> �)j�0�����C@r|��D�^'�;P(b� ��?ݾpۂ.��t�zn�:�rd����R��dH��Ȯ8ul����������5�j��>�?m���N�_B�ٽ}���!ma��OE%
M7��j7!�]J�m�t0P�[�%��T� BG_��Z�M�+�I�D���F��&��ԼcZ䛸(�1J"_&F<��,��r�N�O�Kao��-Ý4���?��5|�<B���a��xS�g�����9��/M[���f��U�mڌXn��GY���׈���k����L�/�~k�(���w	r�Dδ�4P�U9���	����i��Uo��T�������#��b�����<��&�`�Fѯ�]����-|��q6��J�Ԍd*&Z���"�r
'����$���ɦ�σ0D���d�GM���"d�_�`�-��%�a�*7%�\n�iɔLW��� g��AL$a����294٫���%;?x�Ʉ^b��X�}��@��d;~WW#/	Ӱ�JV�;�r�3�J����Y�`n�
�$��
�DX�'~,��É��>�ҤK��%�e��A<_���.	X�@�q��
��#����k���`�qph^j1䦠������绸#5�x,a����)����{�[�qj��C�߫�d�����\ż0
���Ejv'���b�Ȍ�*�����x��L=|�[�8xD�=B���׍�c.sq��xG����e�]X˔��_�����2�@�sd��%���Ǽ� .�3O?�/��J�ﭪ�,�ݦ[�~��+5����8�b�U
�E=�$j'c�h@�B`-|+�r�kq�[l��#ۿ<�_������"���ͪ�ck�XӇ�6�G�^at�;���OT���,��KO�������Y�I{x�/B�R@~b�K82�W!gL�/I�ו:%�IO;�Ȯjg���/�70�^(�ͩ
{���z�7Ӽ/߫��m/�_�92�i���cý���m��V���q�k�&Վq��Z!�R�ڗ��[)o_g�����ez�ԛb�]��+��v�s)swv�5��q�d�ZY��P�ԭ��6,�
���z!;"��sl�⑌:������,V.h���s��->�V\�뭹�8͸	�����♅kӵ��)�Z{�##�&sii���p���X�n��X��5�pA��M��0>i��ʬ�d1�e�s,���\V��g��[��U�l-���/�4��FgLS4ѵ�QU���Kvd���EڬI��g(���.ɏ��J\���p��Y�tlؼ�џ���:������\]��CMuVj�[���g8D���bV�#0��o�#���v�Am߿��B��i�����J� ԬLp�%�!�955_� ��״��_���ްG��l�>�w���f?a�S�ݔ��䛌����ڂr����K6_�/�eC�������;\�'�FV4ί`X�.�&�H�	l|Р��}�R !rY��[������P�ȧPk���*�����S�Ғp7=�9�{���ˍ�yOf�zFSs�{�i�LFG�\眇���S�	[gQ���¤\w"����3�Tǎ�[�	/���H�G��|j��P�|��?KI'�z)f�5�(~4�����{f~[D+;�Q?���)���YD����&3e����y�C��%eU�9�q=2Y��O�iM�f�y�5���̠���nB��/0́�܋q�pR���t+7R�EAgO-v���}m�Bg�|7 �"���GRhe���C��lv]�90B#Pf�@��v�+3��`�ߐ��B���������!�C�\7Oa��Xz�{���O�+UУ9x�|N���	��V����l�os{�WŎ�}�
U�;R�lN�Tu6�ǛBw���$8�X�	�SL(�a��="}	ڽy�Be�E`G����4�ФɨT˥����-cm~���X~~qR�ͻmOqu�R�S�/�Ew2Tʉ����8{�Lt��i�w{X\֍�(�:Ư�/i�Մ�/�MlF�E.�5�F�0�h�/����;����*����MvRc�c�N�OU�� ����n���)�Z_j�q�2�jͪ��TKd]�e����tJs�i�_I9/:"a=]�M0�G`��{�'����^����O�>V���
��(c,1]-'b��s�W,�d���_���a2�q�>�^s������
7X+����&�5�:��eW�B��_�J{�˶9���4.8��-�g
G3��d�y��;�Uz�:~�n�]},�G?�<���H�f�����,M_s��U���>u[B&�������=���i;��k��6]u���)�ջ�l�X5�ݹ�pu誱�b�;l�y��gD��<t���?x<����꺧1���>A� �5�4#�V�ط,��.��xE��XFM[ް޽Ŧ��y��C�����k�u�eLs�һ��r
���x'���^��fq~p�f���Ma�X�:��:���KhNmb������=�}tsݡn�
����ߏK�7}���ԇ��?���A~��|e�����C7X�ikWl��������hW�������{�Aj�m��zx^7tnR,~��a����Z��N38j6)�;�56p�S�,+7��b�ji���wy8��9~9��n�w[��D��id����O�)�n��jޗh����4i\XO� �������&�
�Y�����x�Y��8Aw�u���a��NPW�L1�n���8�Vڧ����>�D
��3/�^0�
9q�x�\���]����9���`�)�29K\զ#q�>.ne٨Ñ�7���I�Vs!j��z�v]~����A�p�XU~��� b|�Aih�g�ӌ��{m64�s�5/���,�����]��b�{;�6��{5=q^rQ��K_�-�3#�^�/�Z��PM!�/U?�u��"Ͻ�'�n�2��r<�e�R?Ԝ9b'k
��ճ�м�m�Ӣ�G�[�H[��bw0z��n���)v�M֫EۧT�&�7\�ʞ:T0�v���rs��u�%��|�2=4��y���3[i���t��;ÉO�k^�N�9N��S��R�|��5&������͋4	��d�R!Sv���������g���mz�o�gʐ�MbӴdSD�?�_����A�:��ڝS��3�����8�<�A��Ow���D��*�����p����;�Yy��<U{�~�c�d�!��9��cҽ�d�)=F��!-c�{;/�ջ:���49��� T�[o���eSÅ�zǙ�a� �U�ѱF\��I �4ިZ(}�"Llz/�Ȓ"[��н��S�TvM�g���wS�:��B*�w�.=�d���$JK�~+!��� 0�+�m����7�/h�G��u�������e������N)΢��A5(�E��Ŋ�L^��h<��I;�x`םG��;��f�|R�	�pbo8ߝ}���l��m�URvq���gw��8zr���hR��}?q����{�e��p~��i��	p�eS*g��?o*�u(S�n*��Z�Ul�m��^Hi�񸑮Ա�[S����u�w�NW8�;��'��=r��W�a���;4�s-�t�ݸ磎�o�LÉ�� ��1ç�m�~��Ҹ���
Y*ˣ4�������_�����!���n�������ğ)߮>�+�5���OD����l���'��}p������N��I���)�����.��+�,�Ub�ZF��VW$��i.��X;�~�Szm�U����.�>]�i�o��ѡ�y����G��T���[+��i�'z��a�����<�!G(x��Ū�xG�k��*^X�&@_�$��Pt�0��8�{5�sR�ǟ$"ծC׸�(�53ڃ�B�^U�׸թ]~�r�G$i�)�'$A�z��e[��@��t�z��/Q�������v����h/�K�ߤm��ҀMX��瀾�?�N[9[K��/P�o�n�R�7��[��]� �-��K��cqzA�G}q"89�UG	�u�sTuu�wX�Ast'��h-0�o�Qs�5���4t/���-���r0zƖ/���ǲ��t׍��	c�FZ|�#;a+�Q���I�!p50��e���hX*ҡ�s�Xϛ�^��d����|=k��B̶I�;��ǥCِ�5C�����>ơ\�BԸˌY�:%�<_T�EF�h�x�&�94��J���Ɖw��u�<Z_�V�;��ķ�;�9�ʍ-Z���0�'���< 4�
��Ӝl~���_`�>M5�ۊΉD<�V}?��:~Ţ��i���J���(4F���a����5�VZ������V�i}h/���R(�yz������vd?��Y�����t��jRS�N��]DX��4��n�~����=O�*���C[��$�"����}R�d���) lK����(?waZ��4nͩ��K���������-���P2����:fC�(�\Q<d��~Ul�&܏x M��;o��A�AL��z�(ԱO;¨$�@d9��P>l�w��e�ａ:(���%v�'սD�OF���&���F�`�\:ۛZ������ۚAu٢W�����Z��b��n)�&�4q5:G>l�!1�e>>3�@L�M��q�@kq�@NU�9��q�
ݻ��T�΢�>Q� ,� D��	��k n�Ũ�àob# R?%-��[N�'��Ҥ���!�*�u��߃�Hz�1ʕ���r�2�{�|��l/���o,}�|�5ѪΙ�hz���g����ub1(��8v�#P�k�i�ʐ��{�xa� (�k���v�B��Jb.�����Ո*G�q幧C�x��n�&���=w:���kW�b��%�E��ɴ{Y�����K!�����cHg^�J<�yo�o���nY��+��
�$�'W�����£�� �?I�싶T�!AX=G�ۈ7mN������t�!9�6�"D6|�A˔��H "�(0܋�7~-Q�Vʿ&�����%�RV��J��5U���{�Q�m\��$�E�;��*����T�*��C�",����q����-w�Q�Q{2.[=��J�a�y$��v���)q�~�:S�T6u,�T���{�����+��2�W��D�`$�>ܹ��`�7?�����y�K.5��ࠔh���˵��,������_IW/Z���(��Me2��<�������Уڤ4E|A�eU*SQUi9�`��s��i�6qT����r}��̫�(�(B�~�܋�}��ԟxl$�8<o����}ښ��#7�73�n�/�ә%�H�}�МG��2T=� 26MQ63�[I8���ё4M�Q#-��D����L����*3��݄z�$m�v�W��v�mBS�FZ����>I����U\�j��Í�$}33CC\�1���H��������|��7���ER�m�y2�����Q2��� Eb�K(jE��hW�S�@�� >;~1����ĩJ��fd#��NG��� �x%��>D JF"�4���p��|��*�՟���A�p1m�I�J�r��pU��D�B�����?����m0ɹ���Ę!;��~G��k�v���8��1wFm :���f���!�����Q�T�I��U�H���{.��֦nk'��.0m��#�AO����y�0��С��}�gq�Y���vj�v����,��.!���+��E�r2�*�7y�F�ă�*{���G�����kZ��چ��7�9k��k`�>�]��K�
�s/���K��wA�/sX�6��>���(z�8�~]9g}�Q[#�$���oюNb���+�N9�0��Qf���������?�ӄtézu���-o3�Bn�3T�`̽�te�������=���\�&I�
G{����W�/��R״6�tV��O��O-�r#FU'4���*?O�5!�Ώ7�Y�(����pS��'z��̏�k1�p�ɑ�K�o���I3�������� 
gf��$<Wr��M�����49�$��	)�����~It�2��3�{�)�vB7@�7s��c��a}�j�}�ct}��4m�VgV4�C���_=M���qͿ0�L�=e�V�YN�ϫ¤%��`[F�A�0�g5}Vg�D�W�����,]���ųg�ߖ���}��gND����%}�3��"<�e�b80LUƮ��HsێȒ0A��B�0�@����Piᮻ�N�:zj���u� �� ��<f)��I���n�þa�r��0Q�6��%F+��o���ى���.��h:����?��e0��o�OjV�e��5��ǜ��)W��)~��LM�S�F>B`��������pj|���TE'�<I�%8�F����-.ŁrhtM�bD�k�Ku���2nV��u�� ''Ck'�j�z���,��"����EB�u���{t����,���,�5��cN;X���÷ӟ^6VU7���!���d��CX��c���?�����=���6	ak�x!.����-
����0M�9o8�#��"[c]�K
9�.C	[UV\��e��"x!W�:TF������l�9*/���D�$�4�*��BDmP��	ߠ#��S��N�;$��4nĨ��A7DIi���ش����G]'��-�B��a�m���K1� Lb�bB�xz�~�8R4K]��=�3ť�Y/*�0M�Q��'F�{c\o�zbِρ�qU�s\�Pw 6\6���ھEou���(�wbZ],ձ�SN��F�hY�f����sy��e#>E���y<���k��z^D�~]F��e4�Q���V���<�y
6�����k�V�l\(u<ޮ||�Ky|=FLڏ����1�GKk�q65П#�,?~G�Ԩ�#�Qb�P�)
ŹzJ�� C��Z��{�k���;��H�8�6�񾧉7w�  %� J�p(ŶV`��p|e(��8J�������y�X�k�������֛滜�܄�v]Bu�VEU���dЃ�	﾿I���@�i|� o��燲��5ӈ�J]Jי`��F�0���?�K�B��R�4E�� ��1��k҂���0R�b�2c�-��|:�.�g~*�Hs��S�N3F�V�|IF���%�D�F?�ix�4��ye>�X�8��&�(6�}l0��>mǂ��k��2��܌v���jdx�=F��������D�֯*�5��d�}<��8;���oG�����=z�
���6��?4&J|����a�!Xȿ�� )�6q�9�{S��u�Y/?3��E�/�q��ɭ�tt�����&��W�E����
�".�e�E�( I@T�����H�*A@�� 9JΌ�䠒��$�9����n���Ͻ�TW���SUӓq�+�0����@���Ը��o���෷-�|��-���vO���>�԰�T�%:��q
�q^AQ�=c�m�}�]s���7�#w_���	y~����
ާ^�q�B����x��]�@\�9L�03+�*��n�����Zh�uw��;��N5�f�J���'�9�]�|�Q���rT�ɦ5+���wY�^ �U�߿=J�k��rW����͝���K��v.��t_8�s&��u������P�.D�8�t����{�����OS�^���y��_���S��}��7����?�^9z5^�E���Dة�|׍�.Y˛�W
��++�.:��2��A�د�ةg��lվ�n2�H稍��&	Ҧ}�3�vg�u(m}�@�����Ř��N`���Fc������n�/�ݨ�A��,��z
STb�m~���ዛ��r�7k^�v'H]��ɂ7кn0ts�E���5�Ǖ�qu�Kۑ������,��l�Vwk򡬂6��4ӯ�o4B|�j��'�#��v�g�'�v�v�ۊ�)U�%"Dc%�d?���~�Fu�!Z'���Y�i��������}�+���%����ŝ��s�z���ʎ�����3fu�y3ЋjR�p��>�PM��mZ|�Ӓ~�G4��s��/}�XB\9��?�\�9��!�hy��gk��/p؇d_��]_��)�ZB�&���#Z�\�dZD�iKύ ���}0���T�E���Mk;D��D�_nw�������s��mY2�/<o<h��� �c0e<��h�M�FJ$�n}��h1�����(/x�i��!Fi�:�����l]%pcPDO�m�H���WH
��?X�.�����_�ig�����}kR�[�
�� /��y8��E��l��4+��w�M;�x#�f(wluaa�J�.�dbxn��4�����2z${%���������8q�����d�*����O�5���n�;�O_|�{|L(�X/��`(��b�ͪ��j{�T�L�'�1S��EE��Y�y���l7Jn�	��˭�k���OA�t(�>V�/SCS׈4�����q�7��,��B��6���I�Ш4�=���.+�T3��ZE�C��?Y6)t'FAL����uDf���W��R��=�S���M����tf �S�ЎsRV�SVR���C��A蒇M�%h�S�ZO|Q��í�e���'����@��p�ֱj���cb��ַ˭ϟl��2����h֗�;#-R��#���P���� H�e��1��ц����׭5�ow��	ʏ>w��u5�� �ho/9���ZJh35^�܏���+�)7]}���;��o����:��)h�M�c��d��h�Gtv�[��vT:��&�5�/��0�^td1{���N�f��)Q>��ҜMn����ֺJ�h�����8�W��x'cS�J)��J�v���eNA[- �4j��E���v�ւ���`'x����W��_�n�ܠU-0��Qc[���Ug���  �/H�tz9�G
�9]m�t�}��`U�뱐�~Ӻ*�f���.<;�`�������]d�X4u�=2$���2|�K`���J�;��9`_��VdZ�i�޷��J(f�nN%;H�&e���NaS����|�")�ՠƟ4��T�;X9<�u�O��R�u��/������Uϓ?_��:�p�Xp��[�W�^�acػ�X�]V��~1�o�5�y�����w�}�f��b�^����Ph�y��Ь��>;�^^f��ҫ緐�?
C���{];"Iɐ�xiQ3�8@�s���ûo��j�.x�m惥��y�}��:[=�CL��Or���8�,gz�%5����bp�!h�<������X�
kS%��V��<K�Y��c�u���;������O��]x����Cjw�+�K	�D���/�QA<��}X�Q`"���c^C��Ә���5U��3+g�G,���f<U��+rn뗔݃�МU򪕡s��^�v#,#J��׏#"�4��[#`L���+u}�f��$a�<�a��w��,a� �@ET4s�e���*@hj�
@h�M�O�l��zZC�)l�;�TӶ�^�,hz� ���㫡�j�=�^:��^*<{
������1�u] ��%�f�������op�X�7M����a�ir`����^�ʇgqm�w/n*��Y�!�N�6�d����d��@�2�!C�0R(�q��t�K@I��Ϛ��h!�n�r;1��b��	*�1E�������T��o[���A��ޠ��u���2��ܑ�����Z~�hH:^9º
3�u�,E��h^vO9R�Jn��c��?��o���H![����֛RGO�[��oJg�����oBG��>�ߨ��0�3x����k�xj�N{���r�@�-�aT�b[��r`�'���ٸ/�s H��oN:��kE *=�~dՑy
��x]Tp��gx��Gr-яo<��_,q�T�����,�V��7�%7^�ƶM�KknVAd�f��1(��l��~b�6L��C+&��c�	�j.b��7�!��|��)3J�@�T��d�LAJ<=�����Dd�T�w^^����󦼒K���g/<w4jS�$t����9ǘ���$�݀vZ]&ds�(�4���?\˅5��=t|�Y�3�5����u�qA�P�Q�6�~QH�30=������1���m��_r�ǟ6 *x����~�>ߓ�]0u��ZVa����IUN�+�U3�
�'?:F|||���sX�ΐ#٦�v	����p#$U89��r��a̙騅����2䲫`u�F�_�Aߒ����<�X����[Y�}P9�_iL�$3kDk�RH�A����>p/}�!
ȸ�&�΍�E������w�@>G��GVZ�Y{��V��ޥ���_�i��,�Q}ݧ+���44@Y=�۰�z�V��>�����k��##Ҧ*���}�v%Q��K�5�ZxM���������x ��wB��p�v��"z���
^dH�
��`j�t�v7T��'��甪��t;;m3�H�Q@�Ă�4Rm)�~�<&��?R���ӽU�� ��������a�P��o��4��Ӕ`Q;����c���8`�G	���@M7!����3 L	2̓V}�h�۬��V%��<���7ch)�e����8S�βֆ��
�Z��	1x����WW�� ��
Zz��\4Ҍu%t���.甼�K��Ѥ�/n0���(�^�N�2D~��M3�q��,y�)�c:n���F�6���eN� ��p�8-�I�-i=qWX�	
Z����z[�A�����r3��O��
`�c�a�\�~�h�C�2�/'�.�NX���9'V'+�K����.�v�X>!3�2j�dp8��`����B��P��,J���f
[Y�L#�ᢰ�`Xv"�:�c5 ��e����>��w�0Z��|ei�E�`O��qT���u��"_]�=ZM�.�ذ�2��\�`�^�ྎ�Gf���7��l�o�M4�� ȴi
�z	��t����|����ަ~�vWWCNtC�N[���{�U��	��[�
^��\���a���G��K�㟸�a�D��W��~���xo��@P�#�RQ�|R�#�n,g���0���\���ԬNl��,A�z�k�޽,-��,�/.��h|y�M*�
հ�a-�-�쓻`�^�,���;�8/WP���(As2�Aq+�[A���^��&�|� :��x�Ī�Gº��{e.�`�0�݂��z�A��<[��M�Z�`M�G�.XzGڊ>
�c�����K%�$Ô��vf/�����?�y������Ѿ���X9R1~Wx�j�p�M>�13����|��՗��Pv�K˪ǰ����j�ӈ�u�;'l�K+Ҷ����d)�$=Q��k�y �~S�a�_��"'*�m(|8�/�V+�l�������4C��h�7�Э�y������odےZfkA\����wH/t)����6��I=��vp� ���:P|;�0�.,�݉f�uXﺸ_�J���q�MgQ��i���:Пv����L�I�f�^�r��G�|f[X�w��n���H������D2��o�q���8j%�֤%63%=6�v�;���2����|�כ&��x�&�||n#&�K_(	��|�y�+��?��5"΢=F��?:�ef}�4s�ygvH�3p���|���h�Z�����s�?��N�z���QЪ��K0j�/����r��G�<f��]'iAւ_}�|×>GA�u�1h������/�U���V���H}�)���7����:��tƇ�$��n6��
����.C��cXtޅ
�f�H���h˚j�7Ո6纏��j2ɯ��j�T������3�V�ċ�U��#MP������֣�S��U��[��k[��P�8��V�Z�G��7t�E�ʗ>J�~�pd*x�CDT=�Ѳh>�����Bz[�D>7�ʇ���
y-���Ϩ�C�;�5����`G �c�`���A��������
W�B��6���=�Ǻj��S{瑭��폳��������D��#l'^$���*ϙ�1iAM�
:��3ɹ�S.�l!��V�W�� 'i��dD�w�*p}�c���Aj}�q�?���V!�!O�i�S���f��	���I�&{>0�g��U{������[v�aZ?��ƈg6��W$fN�H.����]�:�23M*hެz�#��ْ�V�G�����ں,4U��!W��s\��ô@sߟW7�����GV�=��m�t(OC~�D�i����"���c�G�VfI�$7*�g �UG����e �_���Hi�ɠX�P��=[7P�Z�&������:�� ��!�&~���'�F�j~�f���r-�3���g���<�Z!!��}v�ģ|����L�j�y$�T1V�i;P|��u�*<��-��-���<K6�J�֛u�hu�|`���
'��lפ� ��.�����K-��+;��IE�hN!��\��<�=m<������x�Bc�j��V��}HDi�ؑހ��7��3r+r�T�#�5Iw�Om�XY��!9�ܒ��L
��=� NQ�K��Ȫ�V��ֆ��.XM���Tz��.v��"�׿VL�e/���}<���qH���kH��`�g�]�d�����Ԧv�c/ë�֌�q*��{1o�`帖j���E�-s8�k���"��Ú�{�a��>������k}I3��aLe��k����������G��S���?��̤Tn�+n��l!��=t��(*M��'G��ۜ���|7%�"p�Rrm=������]����y�k�z��6/6�h�q�$|˒�]��v;.hk�os*�a�K(�	��oM��� �	}
^�w'U��̀�dA+�$f8?w?��%O\h/k��#�����Ҋ!�#[M�pX�6����&O�%̴�X�8���Y��ϵ��rM&PW���c�~�ȇ�:�A�`<L�=���P39F�qU𘛆�=�c[�0l�Cv�ap�_�$��H�����5�L��  H���"v��Y�V)b�xi%湺��x��d0t��Y0g��2��kcյQ@����Cߘ=�fa[�X���(�h>���%n��>*���:����Z9G��z�=;(vB��@��W�Bi��ʥ�R%
�;@VNU\�3��߭u|יdI.��6�6�h8솽���(�R�#��5Q�l5�y�w`�,�#��������s���X��c9x�Z����=�Ѻ�RG��m����SJB��aj�4��k�v��U�u�D���(���&����j��P��R��?X�	ܪ�@����N�w:��ܧV�������$�9�6#�Ɔc6@M��:5�q/�1A`Kq��>w`������!� UV��c�)��a���k@�C��&��U���!X�X'A��#h+dM�����|�����m� ��^+�V�yI~��
��ɲm�#�����S�M�*��Ӭ{�a'h�����{_!7[��3#�l�I�ؙ�A9Cq��[q٪�)}�8h�^�EIDHVV�;������췪NnXT��o��D�R��]�U��bG�#�z�&�C��|Pb�8�[��M�8@�ix���ۍ�݋��&Jpu��J��T�蘵S-����d�7es��N,��jK"?5��|\�!�
3�z���~��gL�P�EcP�>\!b��MYD��ph`n:���tN�w�,;4�����o9�k�S^�}\���E��l�[v�gE�oϚA�ʪ9��g~0[ëbF��]ѻ.���S+0}�Pn&�JF��� ���!�!�C+%�A=��k� `l�}�I�4{�T Z��}d��k-J����5{:,�#}�$E'y����Ǟ��/8��C$퍬����;n�>h٢(i�
�i|n K㐡�s@Tvjn��V;�qplG��áC��cIu��	�g��2��|����\>�$PG�-N4gQ���XD��<Ą���ʎ�Ab��%t��Y���h��YЀ����%v�ʹA���7����\��f�<���� `� VS	}Ֆ����~l<�b��ADD3v�j�j�V�� ��p�f��n{~됡Ҥ�̱��79\\���#�1���$E�xiS�v1��pͯ<�,�X�Wt�����HFQDM6�K*K�c�4�c��l� m�Ϛ������I+t�o��ʶ����܉��L/^�ݲ�=Q\��"H}&��E�+�Ӛ&H �M�;�]��UmĠ��9�����>�:��
�՟��$��|]J�o1RG"S���u���^��|��V�Vv鞙o��	NC]�0y�w|�^H	'-�q��C R�wE�՚���E䔠;k�&t�4xxw�������� ����Yv'~.O�#4��Z��<&J���j`�˖h<H&����R\�%�g�n/t̚��ȍ+��gy%I���@�H�|P��^�+FX�`<Ϧ���Pn���Hv�4 �W���h#̢�+˽4#aih�*R���ZU%j�&��w)A~�S��<�pw����A�#��+g˓$��3䠡@�g�{�&���'�j<6ж�2}Ը�����b�y/}�mh�ݡ�0��`�<6���Jjj��?L����)�!�%z?��^Q�������W�U�M�ʹt�3pޛ�S��̌�������0�,����_6�d~
��ϛ�d"G�C��x�����`���*��D��)d�����^n���c�0Q�Ȧk�;\�0�]g������u��̖����c�S�������`'�m�(�yi��լ���ÍY1�4�� �o�	��`�2#�Q�:��M���<�~A�)��/ESb��X�5s ��Kj�I'���s(��#��"k�%C{��PR�B��^ڌ-[����s��� Q���GG��+v�Vɇ'Gn�à�γ��ؐEf�����4��7��}k~3#�ަ�ޝ��}G������aG���OCV�)h{�;d�9Y��ڎD���y��5;�~�k�!�����t��`�KN��k��9fKT@%�ύ|����������86u�I��Gv�!Z�!9XjˮH=?����@E�����j�ƾ����|�=�`^�4eA
��BO��')ߋ�f`�pX��^�3�jy����5����$@��uy�K��j9iA(WqN��|���t|��CG.�Xvk�Ճ�b�Ƒ�w��x4�gl��Yt1-	��ٗ Y�i�*��%OU���߽�߫ۜ����E����p�L�c�%>�kdB��W<c��4�cu�Ҝ!:��e&⤫�CxVI�8E���T]+c��pXOJ�c�w.�)0j��6��4��
�'Dk+p�M����6���dp���F:=�
:qY�=Z��ԪuP�Z{�H��f-%�����fs���w҇��x��2O	����l�oq�i�^�G����C�!<wA�;�yX�Jn����)����p �����S �����=JH����P��jq_t�]+��\�nTv��,�@������O˭�9ORk�4$�,���4C�(���3���[���0�վ���H�r]2y�Z*����;�a5���T������ݞ�_����%z��`M�G7 �Wf�P����er��[�p�[@����_f�,7J�`vV:�����m��9#�W���/���YZ�+��������m2$2]V��W�'�vʗn'�ykKq��@�w\݁J��Ϗ�m�5���
d[A�w��piz5ʼ<���e	Ād�Q9�k�������γ�;ѳБ�᫢�Se���N�F��^�D6{�
�rǖ�L���OV��
nq��e��0Γm�G
Ι:�3�H�>�knrGO���WC�6	JƆm�\�F.	>ܑ�XJڙ��Wp�H[��_�>;3(��ݰ�CB��<�A�l@�76
�wǪ]]����A\Iok�Ƈ$ᆝ��?Y�t(�uS\�����\�	�Sn�'hb�M<������^K�uA�9�˚�R�ӿ��~*Qh������K
_Cy�B���Q����m2�.I��?���g��I���3~��y!����_�;��x*/�SՖ�z�n[}�y�#1"EC�i�Es#e��uh�F���-���.Jz;���p[��2|bk�(�^w�.J����v׊N���p�%�H���JՍ2�<�B�u��&�I}��5Re����hPb�X�N���Ty�Թ��#�[R9p�k-ēUFu�Ҽu1�T��i^l;X�����E�:�^T�.�P��։Iѡ\ޜkd�/�G�Ə���%�ts����?���Ks��m�\�xz����&����!aQ�^k8p�@ʨ�Nc2}�Nf�����u��|;�6Y��z�2��;d�v;[�"���Yі	��VK[���7)L�����D��ų�a��x;e6\�?�١����@��H � ��3e�͆I-���]��O�H&�MZ����V������/\�����ɍ'����o��́�~�����1S+���1�7g�K5�d������.!]�ߚ��}�k��Y��J:j�W����&���=x��\b�s[K��F#�6����;m�6ڳ�$)��й�X�#��Wp��f���t�\��	�yh�Q��e}�yv>uZ-Cw)����-\�n�q(�od[-/ufo �M��)������'���2���gsr�wN
_�^pKF^;�y���V[Y���~�y#=�/��k��Xg8�&a�Ŝ�?�K8����ĭ�և����<,��<���;u��1N�N�����s�E\�Z��>��Pi]3T	M�91�"h����Hd;�c4���>>C6���7�K0z~B1�U�R%-w����r��[�PUmE�Q�lC�MRg?�mt����{��\-�1vh1��[�Ha�?Ś�Ί�GG�.C�W�:jpH�#/_h��E���b}��_KM�ߤK�P�x�h��CB��\c�� �g�UrU)����e�8�ly�գ���Y�AU�����Uq�%+.��*몔t�+���rFx+ �1='1#"�6�!�/�#\>I�?ozģ�U�|Rv�YC��߬G�WXR�_���u�Hz�Z�
�X�h�{P5�U�ĦڈK��\�6f?�p��vp��u���{��8%��*-���~gi�J�m30f+@u��!���
W���u��ا�;�%�z�ǻuI�;
Ъ���xiJO�u�9b��]�a�òev!~�֥�ó[��*�Qy��j*�oe�밉��Yz,	�^�ͼ���߮l�`��<�5n��u0��q��r�XZٞp����~fmIF�/��^�n�y�*Y���El�)��,#O���ޜU�>��r_�{b?g�-�Q>́��6I����k�bu�F���*��ׅ�?�xW 6��ګ1��
N∢R��I��+���)Z��>?".Ñ*������G<C��{Ҹ*������%;K��IP��L>S̨�	�d� �a�/F��"�[�ӕٍT�2ˢ@�o?��%�u��c�^�񗞲�zOlĔ��[�|ccGh=�㧝bP2	�6�F\��)��>ҿ�M'Ҕ�2%��)��=����}�3�G&!�9f�]�a88;���-��B�������pp�:^�5Y0����v���aS�P�w�!��([p�Ύ��H[����w��8q8.5��?���S��X.�:�n��y��}��H�u4"�ɴŰ�bP�̠�J�^�[��)E�׉��`
���4�e�,�~;�M*��*�D��qO���5�!R����a��qeb�R�+���.%wq�g;!oiC�ۤ�6{GǠw �(�Y���f�~�������E=�p���c�m��ۈ���ד���9"�5c��Ha$���rpi��7\�x��t�ߞ�ۑ�V�s��6�6�b��k���;��N"�����L�$z�2E6KHwO���Zґ�j��N5��U:nq��z������la����U�K��!�rq��7�p���tS���Ti2��J7~�85U��H]N�'|Te����T��γ�r`Q(Os$G�����qi�LK{}��|����a�L-"�l�������������xڳ�fY9 :��Yv�f)�QB�F����+_�g�\�RP�
Иmh����CB2y���|�!Y�)��KQ̎7���Z���ZmzFN����k��}p��"�M����1�� ��T�C���/�!� K�ێ&�
��RWĕ���
f��{zEC�C��֨��j~�{�c��Mvވ�@�\̠��咰�*/��/��FE�lq
f���������ٖ�~YN�����WD�������jr��M38��j������?�e���z�"�
���cSƿ�r�3\J_����7x��
@�R)���A�9d��o��֝t��AiV@=H8^��/�Xf�(�tG��x�&�r~��8o�Ӆ������_E���'��;�}�i���MԖOM65Y�~2� O�\�84��u��sC�(d-R��gy	K/���~9#8M6	b%iP��)�����>��(8;��^d�T�UJ>E�;�[X����I`�W܊�0���3Q)��B�v����ld%z%�*�1�A�R�#�6�[T��:�0/[⃔m�qb1dMY�Y*��k���l���g�������v؄���Y��G�o5�h�+~L�G�'(��u�-��^=��B��"�R�Fl2i+�_
tts��:�s�y��1�?��o
�fgޚ�^��D:�4�˞`���p�뵃�KoM��60Ӈ�A3`�b��>�p����J.�+��Q�2���a�;�7��c�%"#kD8Y&R=T�#}��X1�$�nw��TI9�w��uM�-I��0;�4�B��.|+�Q�?dT`���Z��x�A�P�<p�3���F��1yr�1I9�Fr)��#0�N%t���_� ��J޲�!�B {A �r|��N[�kAA�� ��R..6�Lt�C$ �[;r�;�%M\�s�-PΙ��YS�%�+�0��'��s� �Hn��%�ft}��pȾ�����H���b*sSr��'�C�Zݻ'��0��l"ˏ/�|�eqW��8A^UlLh#���	���Jq���' ��+֐��m������Wl�HJD�+۲�TZ{ܨjS��5��h)�88���V1�?��B���'~���ɍA1hpV0���S�ho`;ڈ\��'^b7A�΅���M1���^���,��J��%D1C��*�g��/q�NN:M2zQc5�r�`�<��=�'_
��SX$p"�7�#	f#��(Ys����#Fp�6��:���5��M���
�3|_��W�S�1���BSн�;��+	+-�Hz�}�*�8?y�Q玖3����R�5Cyi�D��!���ն�Z��Ԟ���{�Z#�dq�u �����Ր������<��� �o�R�>RJI����+��i�E��d��V�4�m�����o!�7�"�ر��ˎ��+T�|K���H7�V9�k�%�:!�v^�����xQ��XŌ��\m�d��*�,������}�?������V����-4��	0�U�H\�.#�S&cn�@�v{v�o��)�S��s��k���B����m�=�\QG������W�il*F3���� 6F���xh�Qe��l���ь8�HJΙ�I�s�"�ܐՅ�߳�w�fX�?�ͥ3�c9K��ݚ_�ڙ�p��A(���qA�d�=2�rC��[�%6+��'��h�2�'����Cs�ĸ7�N+D�
��h�Zm���O ��F�˕�b�5m�7�ۏ~���Z�߈���.�x�x]Z��S�Қ[Te.����(RR	i{������aɪ6�Nd�E)i�R�&�VP<n�wd�:�����4g��{��{l�ς-b�u�_�\��R���r�֤2�$�")'�Fpoρ�]�͕CU�y*�b6Iˌ(�޲�Z;#�+�[i��K��|���X�e}���%/U�@ 9._�N�cWS�b������aA lsѩ�����Ǔ���xࢎy*���.{��	���!�m׺��nP�����Fy��+3��3d���Fmr��xz��yz�x�9ϖ�q.:�q����O	 {�?"h��f�����V{�V�0��S��~Do�?�>��pf�yF_��ףM�(g]X��P� ��2��%uZ��=�Uu��n�-�=?��'�\T�1�a#��sM>��6H�z-�>�ͿG���P�tw.YbӘ����T�9:�^)eRO�{8��~�y?4H�E��WX����VV��A��Ε�'�����=C6�F��
� �d�j����]%�~��-�1�������#èE]����Z�q��q[_��v�����SKM�Pm�5�zZ�j�����Sv�F���9U?��a=B�o��g��!ݺGzWg�� (�SM{u��k~��&s�bu ��OA�ow'���욭7J鼦��m@�J��>bM;�����8%��؏�h����*�X�8�j��T�uR`�bu�G/L}`��|~�S��R&��г7y�ܡ@��(��0w�[��%��Ɵ��vf$jH�b�%'�,2�W$��44_R�CFԉ��|n�Vy�@Z��
~ъt5�֜#�d@�{ŵ,�
��4�8hqX�OTv�q�rƟc|��W�HCU�h��'���Z�Ј�AQ3-�����~��wF6Ih�QB�O���Z5.W�J�eKOUq���%�)oT�pB��*�pŕ��,�8h�/��	��=b�j#�"Qn��;)п��Z��~�\��Q�K�n�U�L�A	�R�
�:��!B�>t�ދ�.A�7��ȫ%���8.p�`
�{�4B��{�5Z��3dּpń��L-�.2x�P�S���q���f��_S�iځأ�v �A�h�@�bhm�Ju��������w�E�pE8_��^����%JP@�[i�k��~"A"A�eǞ	���H��.F�n��b+��#�� s�ˇ��ࠐ�W)&}��z�Ҍ��Ҏ�a����!3��d�؛#�oP@�$��:wc��ܦ�:����Q���!PTP�lT��"�?��݉*��m����"�n��0q�M��c�ه~ȡ?�h��⦾�8�m�p��UX+��S�?������"m��t�6��{��Y�_�=�̮ߜst��P�!^�x��L���;U���������1GȓB J�*r�ða�ӯ'�SU����P�l�C�6Q:����� E+?��b�6T�+Hͧ�f*�MڠyAjEE�E ��UAE~o����㭠�g�>hb豓��]�	S�� ������N#"�:�����3�V���et������'��d"L)�TJ�NB������j73���
㻑��	�B�/����1��~0ⱽ�-�#ѽ& �s%�r�B_@�����?��,˂��V������BۜȐ���	i����gU��ʵ��؈�h@�x�����7ȯk�ǡ�
��z��_���1��՝���u����+$hU)f���|n;2mY����[`�]L3�@�?mU�%�C|4 |,��S�k��Q�l�U�NP��E����P���z������Ϭ:,{��C��F��o�H�e�0��T�D��&���q�@��T��#��Nn��� ���%�h����OW�I����~�#�W.�Ӄ�q0�GDƜ�R�8�#Ÿ���+te<peɽ�1|�g�j�,C�/��6���G^2Wl?�����ϡ�X�W����h�kw��u	�{���%w���M3R�
9�9����;�V�L���+C6����g������/�5�SCB@���\��,�|`UƔ%(г-o+bl����L��O� S����=��6��`�jëeK|*��l�D�u�{9�0Z!V��ݲi8���T���	*� ���͉� ^fZ0B����ʅ�	Ј}��2�;��-�Bn��lu� G�V�.�E�j�"���ƕ��L|U�t�_ѥ.�̰�*:��[P��m�E��ĖĈ������V/@�7�#ı��̃X�8/��#�nhN%ץ�dl)~�05�f�g@��j�	�����!\�ʎ��.vk�"M ��JH>O�}b�y�"��������!!�eT�>����L��x�i��3a���X]_[om����uE�� ��j�2��B\Va����P$ >�`P�O�����3�g��fsCTڗ��!f7m��H�?��ߵ��G߹��R��B7���_-�?1(��Ȑ�3�`ۊ����m+��e- 0��π5�by��<	b�����ܣ�Ou-��~��|/�MY����F�B�!��Ȉ[S4l�h�h�a�y[SS5F ��[m��-67� ������x������ݣ4S��.2S��qP6<f���o؀.�(`���4h�޳ 1�ԭ/X�G��z�k̍��Z#`��F8�;e�S���%Q�Z�rK'���- ��Zܙ��,QE���Y��W���aN��{��
�`p�̻�KU�^@�@U��mc�����ݿ�gj�e1��� ]� ��:U����.\eW����s�<u�t��4N�Ha\���*�KY�*sw�4J�#�e���=��3�����?�Z��(���ݧ���$)���9D�%���yt�N����W��=Q�dd.n[�t�p�V-�Xu��>�S������-n�!���x,�m�Q����Q�"tC���) ������)��h��[\:�wu��1\8:J��}���=�y3����I�0Zu0[��8|�G�$Ֆ��5W�B��bj%ܺtXMH��S����m/�*����YhMk�KO�����pe�[S4��zB]&�O3i�,��Ok�����4aM�x�#��`�����
<76;����p��K�U&f��\M�"U�|��з����;ɸ���+����X3�ʣ���1K7q4�~pE�є!���U�A�-Γ1iD��cm���h>J��=	.�l�b��*~��˃&ߩZ>UmÎ���%Or9%������*�����_�D��CK�A-����U����!��f��aL����˽O�UA�z8�&�P���ϯpd�Î}N��(`C1b���p10\�;�u�9���?#7�����2���a�RD�\�(�ވ3��y�c&>�Sz�p��O�V����n�8�ޤN�"�
��B�Xe�'Ǚ�3� j�j%kw�/�v��G�\�(�aI�����u�XE]n.j��Q<OW�\�˥�b�������P���a�����أ����mQ��ә��ع��#;��l�LN�]�)��ZΡ��ǿw61�|,U����1$컦B��ッ�s}V����&ͤY�FN<@���o�Rp�Y3h���	/ٚF��@<)�т���D�0��&+��χ����aW"V���+Ή?w����c{'K��L�����B���H	[�t�$�t�D	pm�8�%��]�߮��+W��mo���M��8�SZt�3���̠Fd
���?��Ҷ��S�ԣ��<��"BHHН=12J��.��V3�Y�n���?`�$�s�{n�y׻%�Oc�)>�*�<�\���~�!�p���w�z-���Y�~��=mf�p��ċ�ʏ;\���_:��"&�5l�i�9�A��(-X�e�He�$α������2h,�U�nʸ���(󨇥�>��5�0g�ܿ&���C:/nW,��W��5�ehЯ�C���3���t�����x҉���0�f�a]g�ց� �0��G������X�����Iyx}���Y{s̔�����犻�pX7r�'�aU^�Ē�������UM9�((���e�II��U�>�o�/���
h~�<��񳦮���7̷�$I����eУ�Z�-�'P�$`��0=���a-��q����3�G �Β�]~Wyi���x���4��X����1��JSH�4�(�f{$f���'���E�Hm. �����p@�i��?*�#�Uq��\8e�xo�����ar�$�K�G��p�h���]I{1v��T��XA�'h׊�ēE���6:��8�H�j�����"��4[]�	��Ұ����Ui]�q3`a��j����@��̞����[��N2 �'���˞���\('�O�"�����~=��>f7���>�`���pS1&c���ՕÕL�-d���Z�^���E�3��w:I;ے�]0�@�7�+�N�
�;r�@c`n�޷�Ѭ�;[�n���v4���_qÈ2��7�]$��e��t+OIZC�A�@�oE���N~��
�pқ�	gpK#.�&[��C�*Vop8�x�P�@��e
���g6�oe�3	�G�����s�hV�t��/aO����p�E��+s~��ľ���\�~�����S'�mVlk��� L����̹��wml)�ZF�I�����!ʶ�#��?�2Z����/
�w�||j;ȉ����'��].!�_]���-~��$�ϴ�I�Ǹ8�?��ߐݐ!G����̴M6}����RQ+ �|�d��/�K�-l���Yo��'�z�w�3:�a�ޜ���2�˖�������P��Ԕ��l�;��T��	�.���F��,i��xY�Ld��S� �}����J�-5��;����Ko�%��U}_#�����'�fm!�ds�K�P�}�b)A��g4�^�)Hvs9�MZ+�0�����p�*�����B����~�X�[�;e��ʡ��G��#`�8�5��AyIz�x�YIj11��`�֋���eYt��RWU9��I��/�@�pX�$������J�|P]=��?�6߽A���P"���G��ey�	,W�= R8F~���� ��y������Ǟ2"f��m�X�#F�ڽ��Q�ꣴ��[(�vݩ3�1��nc�Kzv�$1e�( �a�X�w�2�^��\��$s_�g^胢֐�~"ހ�S����aW�
y+� |]���%{T���h_x��x'��{�¡���a�/���{N�����c-�{	S��yW|`����$�)����5��`��<�f��}y�/NEU�]!G��3�~qF�D�h��O&�#��i�	���Ͷ"%C� .��4��{Z�pC��o�����k��� ;8
!(�;s}�&s�����a���S	r/]�Q�j��4M]]|��XT�?\�o]ue����؀>���JY���� ��"���PЮvi*�a�=�_�L��>�#bI��Q'
�,�|�yB������PQ��s��#�+E����*fM�d媚��tS�<��HH.������Ćy��$~ڸ	J*����Pƿ�2�̽�q7N���\~E^ޭVe����% �\bt�@R�]�,qϻ��i����a������a2�5� Rd�(Z���Zx�b�p�>��m���7I���C�����\��p[�$�@�����&g`���x֤��0�ܭ�	Q��̮��cS7hQ[������K_(ퟱ�$ƈ{|n?�$�M�;���	& �d��\c��_�>����\?�;#~�f��	�e 0YwT�^�ۗLCxn!A��#�3s����O֝�#F��2�M�>���ajʽ'���,; �e��-�}z\�,'.�ZPlh�~P��bx�. �oS��m�R����A���L'CrD�t"���{E�����R�s<�Mxp�����Ed�!���������D��蝵���$�5e?�g\}������"�/�H�,P�:9�{n�w�_Xu{��#q�,����<�����u�P����ఆ?s�p�/	��Xº�Q��ѩ�IG��編�\`��}fh�E��/A�"DV'�Y!ｭ�
yt�@<+���D[�qcd�'�"�I�n	9��oV��W�ЗJ�}��@��2s����l�G�i.�笓xW@�`�vc�}�biU|�K�/N ��j�����>Z:�����?�PI��:B�*�<��M�؇�'��,~>/�����
������&��<�٬Q�ܭ7�%h
�u·od�� +:�̋
a���,j �'B�{�ϑ��BQ,����v)�� � �^ �~��lİ���Vf��-J~A����L]u@T��vX0 �DRR�t¡$�K�Nghp�I���J�J9JI+ �R�1���	�?��}���|���n����Rʺ�B���a]`d�9W�l�9����-�qr��DQG���_~�oXx��(c��%ٗ,BӢ�vP�� �/�f�a�#��h=���#>7�|�>�l�/D���{KvP����L
�RI��[d���bo���U�D~e.��Zwy؞�{�A�����;H�H:N�؝� ��-Y��62Ia��Qu���ٜ�t'�)�	���S?Q/b<���T��WV`����_�L�U�m�r�4�˕ %��<<3֩�K�w+g�s�Q�?A~
�~j��؂��&!X��.n̘��ӿ�X�9q�m�� 	������Q�W6�l�H����w��jNk�QO�h�PXe(B���/V��B����P&���Ax���{�*(������s���������!g`�S��q��s���%1¯'�	a_,8�Hm����"4�Y߷-m;/�����R�������C��y.�D���Y�?�E����P�؂����|*2g~j�2b����)�P�m[�t�0DFE�';a�����U00���o�9�a�M\�YS�&�-�C���Dq^~�/�vp��!%䍬����C(#ť��3C5@c�;������KDo�,9��%�_����Im�E �/�1%��-W���|�a����vh��~y\�U,���|�k�E��ge�R�D�Ll�;�5�j��֭�>��0��-�����:}?!]�X����e���6� �Oӌ���+�?3���C�ߞ��S��3�J`�z��D���z�?�L�L/��-�$��^͌[�/��c0�Y�U	f�	�/��o��bo;/o(���D��+�Fj�OR��0����c��*?��f����� �Q9b�\�C1��l��wz�f4���!0�QN�j*�:�s���"̤��S헛SR:��9��}Z�&��bA�i�$��m�W�4��q�VޡKꖗ@�]�F����������Ì�N	X�w��cCܠ���τk:��8�5TTOgf21n*]
��7��6��V9�BUM_�t��kG���>��RX9�8�Q�Usv���[�Ч8s��i0���A�:�~��߲��B<�[�g�Ys�O!W�Z�� !�/�
)P��A\C.mO���fec�3�ÿ$��2����Rj1�&�u<� ���R�&��	3�iĖ*��p�� M.��)K{����ɴ�M��p�?L������+On�����ު
���t�;�A>wД����"�@�/'W��*�����h$�{؟V���$�gc�~������"�Tf��b6�|�,��@�'y�����V�+8�u`�C`߃0O8Y2,�U��"`����ŗ�>_֍�Dt?
$��v�"�/��oA��&
f_�8��H<�ޝ�fq��j���U`��F_�Z�i־T5����wP�S���/�O��ւ��a�~�1�R�����˺^��=�կs9$#r��_�@t�W3n�J��̏�����g__8��t��{~&&��"ࣗ��O��6�)W?�P��\���G���G�ɑ;��
��?n�ɱ��p֛(J~so�S��vn�9�
8��!'��!=�Hz�*B�n�jt�*pΏ�'Y�9a*)A�o��u	oPoh�a���"��KT�;�x�=v� ���X����9�cf͌,5$�������K���/~�O�SL�|��]�	��	O�[_�xs��\37�(hH��܁�vv�@�����p���W���7 ��9"����FO�Tn^�[�m���~���N���'�,.Uq�1v���u���;M�Ф7�l8�ʨi���A���7`!q6G2�%�4G�6qW�m����~���R@$�=ZZ�Դ_�Z�<�.鸀� 
L�y8vX1����<q���Nz#羏��da&)�~�&��O���{.}l	�WaFP	��p������iPM��C%�O`�p���n_�[Ҍ�$x|��Y�uj��bm���ė:&��g� ty=$<��S�LlnB^��&2��Oc3��������t�_�]H�D`0QY���gc��ܺ���́� �X����$8l;C���@3����
Ǻ���Ӽ�4~�ơ1*%W��YR� S�������3e�����4B���o-�O5���
R�.9^	���5N	��M�~���WYW��|��c0V̚vi���$v���#�M|��Lv���7�X'ر�ڂ��s- @��]��~F��N4���W���0�IY|`���O�m� ɾ��\`�M�`l ���`G
�[u��+�B3�q͌ǥ�g�r{���EL9�&���K�F�rr?+mKmC�(�OgKjAH�\�5�>�D���$NJ��]3
�6i�6�mA4.ǟOs�q�&*��ۀ<^q�>�yJ �;ks�b7Wx�p�� ��/�М0@��@���$%t����uzv��7<�R_(�+��H�Rf{2(x#�b]�rNKJq��W�D��a~����]+��!�Rc��\��}��`��X��b�Y50ޠl�D\��b�#��%6�|~�W�W�P�^
:�� (K���������_4��ȬK]�řH�1�1ߛ�<3:~:S���!^p�e���1�6��r�b�?��$�ucB�d#	��Ƴ��1�3��fu>���D"���wnճA>�d�d7(r��y��e���ݏ��Zy�oH����*�Siߐ_f�T�����?{Fw��D�,;�]Rm,E ����b�O�ϕ�,m	nঌ� �sx86�{� ���#.�-=ҩ�о�I�+��aﺤ�k{�����@�c���fu�a�?��P�en����jOpM��=���A&���m�I	@�a2������Wx�_�������`����g��	�U�_�IQ����,��P�'���r] ~��#!�։��[E��dn�?��IP�����_�����J15�ҳ}�OP�1��_�fr!J� a�Oi��ro�R�8|���y�O�&�������j���l�!����3��G��U���w�M#@�	���m�L�O=���)Yۜe�Hztu"-��>Ōq�m�)t�K�t 9�֖~�Õ�4���.7Y��)�Z�2�><�wm�v� �i蚍�7_m_XW��U|\Nx���9A��2�}�f��)$��?���X!���G|��������ng٠%�<�[���W�V�ߑ��^��)6�}�L[��
yYy���`6����"�[��
ӛ���O��5R��P� =�Dr�|��'6e��,߰�?�<�ݲ�~C�=+�N���_
��Z1#̓���_���(��.�Cϱ�^S:����G�Խ}8�q�-���!2(hq�̄�y���qi�@�S�Di���`����߿�x�K�p�8��}����OϿ�L�ކpp�i��2
ZR�]=zUwh�nnM��;Es/һ�4�
ή��p!>�䗻��"���w���R�,�A����~��i��No����S^�Z+f��I�C
�qT֘^^9���*�t	`[; '��s�g�hx��,u8t�9�0u���_���=p�}Ph��`����d�Z�jY]H\XuR�da�����#�u���ƥХ���������BЍO�����E�K�ߗY{���`���[G����eZe��S��%���y�-���&�,���ss�=��gC�!�ҭ�j��8�H��g����F�9�R��و�i	�<��g��h��oIIP~h]�B")�����b���1���I�b����s�}�2��b<��IV�;MBc��.��)s��с�\=S���b����́m;�)���'����u�������Z�c�I6�!1b�Z鶲��H$�J�ѯ�cV�eĶ��S�r`da#���-�v��$0��Xr�W�N��NIf.�:�̼�Xd����!{^��V.y{��6O|T �;��l^�,e��]g��1������n���y�����|��C���	�W��W�9�����U�b�����p��
����d���Њ��Ί"b��G�pq������n�3%�D��zMI�
cZ�H\�$��Չ��b��EͨS�	��5BYZ�Z�*u��U���2��ᴕ	���O{�i�S�h)�p0sCG�����𩍚q�9l�%C9�&n|sd�_��$�:+ځ�eo�D|I\JQe�&7|�Z��t�0	���0y��і�.� �=�}���LY�/xx�����{�A��Uj�\:5�w�V:(�x�LW���|�7�-d���{�/�Pu���$��6�b��b.d�C�ӣnb�U����}%�*�5���[�0Ã{��b��,޲�v~:`��a]��W�J�Kѵ-�0/ר>c=�a�(e��%���qӵ7�|���O�F/F���_A��L����P�ְ����XSM��13.�,��kJ�X�=�^�Ǵ�u��`]+�N�U��\5��{Ey�,n�=w<?�E2���JK��},{��;XW���xW�����x�����Ɔ��"���v8�,�^�(�ޅ�Α)٫V��tt�V���y]>�Ar$T�$l���V=�i�����1�|C,٩3^�������V彩X�0탦����?/E�GWs����v����+ޮ�t}P������a'n� �g�z��WPH�)G���ٯ\�c������ԧ��M�#�m�B�{{�Ge"����V&��\v��6n�H2�[TZk\;��Fd��G��祐���_y���,�Y0�M{{�k&���/N�,���Okq�۩u�q�����G_
V��$1fKu�J�4�˝9����QE-o���d�, ����
��OW�/7aQn7e��O=�ն}{'(HmQ"-�`����9�Y�H⛀m٥d��Ecg�l{����Cn���˸�a��'�.րxt���� ����3BB���h�w�VHa~��YD67�F�~:���}�Q���ۂ�#"�Lqsz����������Ci�����տY�;y����-��H[I��J��N�	��&����5�c;�S�ʝ&�C�d~N��҉M��C]���z����F��0yb�i����H���s��fZ�'��1ہ�����˔��[e'h8k������z2N�(?��!��`���<�Q�MS{���[���e]��o!3��I�����c7�!��G;.�� �*�������o�MzN���2筱ԇJ�2|-�<4v+���󟌚Ǔ�ͣ�<;���'+O/ϔ0�!_H�~̶�j��n�"��6�<,��J�L Ǯ�p��V�z�D*,`FeZu� *��F~���X�I1}9y���Q�D.�V�v3���zdb�i�����f��Aj���bw�H%������.A�1��ei�.�N�Z��/�6�4aI�`/�fwV6X졬	f�ae�"�6fJ�dE�dV%�o�;v��o����e�6��n�0�̠s�IVo#��N�z����V�mm�33ҥ���^�ܕYv�ϝ;�4hB|,��o�`�#��♙i+��*[��1���s���xo�9�%�{��5
sα�h�;�Egp�[?`� |�1��|}�HJ���?���w�J5<D��:���,�����2|2�� ҾQ�$}���H}oޖO���AP��%V�Ud[)���ze�S��?k��p��=t@էp���p�>b����	��9[�؇��o\��H�(L��}�d݊��o�#�!�sc�s�����i���r��~��%�%�4eK5�z��y�EV�k<%��P�]�k�>ǧ��3�% ��� ����Ǚc��Ŷ
�	��z��M����3�� ���D���n���\)p?0\���b"���:j�_�����v7j����?5����#6k����N�z��������Ԑ�<��8
}�q{�sdax�5�^���U����jքӊaoV��Ɓ��|�<:F}=*E��=$��2�Ԓ2U��&�߱��)�$�]�I��o�A�<u�x"}�}�Q\��BtEjz�`Q�����=�օ�<���VX���w@U&�V�љ<�
��-K�ו]��؛��c�׈�;I��~0��'�z�7����B\�eҾ����Atc����S���祈��f(����u�=�1��������j.�5�}*��p��@��7��2/�o�܇t��IVla,���>��9	�w�7���|�T[mqAEk��`�T9� �%�4�X�S��\�1=�����1�@�Ȣw�T$��b;�����ň��Q>�����z5����}�����jJua"1�)9a��<��CS)S|��6��N�՚�AK��MG�d��er���|�}�e9z�ক��7��߹/$5HND*�j�I�l�Y�
��o�/S�b�^-���⸎:oU�h8�K!�|�1j���>��)��U
;��|�nm$����̣�+��*`��3����u�*m��D>�z�;�bcm������#'��u��aoR�L�M�w�/���t�}�Ƶ�݇��2�m��y�ɝ=��H�mjߍ�t)(��{|�v.�$�s��h�R����D��,�l�X��yO
�T��~�A�U��X<M���v�/W���5@�+u�
*H�@�F��U��:���P�}�t�0e�u�������o�Bg���7nSK��!� N�*O�m���I�f� 3-����5F�a�J��)�=�����񙙷�70��F�}�k�����у�E�����X�_�OO����-Ҷ��${�<0�����s� M{{�����|�T-������"?���)=��/h�kKm�S���q���n�O�طy�,9�u���d^�Ǔǃ<�\��d��9c[I�j�J�El�i������#P0�@���DRC$@�@�v�o�U��Bt��M��Ӕ��)�*՗�MK`(�6~��$Hċ9FU���A�j�Ȗ����� ��C��6y�6]��qn�N8�Z�u�fv&jɿM��V���ci*��ذ{��ٰ���M�t�I�����KΫx.��`�F����Wcp6@6%����@8�DӢ�@���?t����xO{쀿:���-���?�ȜE�������$���������J+b�F�p�8V�34UWw�c���sD��̰���� ��~/�t�+O����M�\�v�^P��]�R(���G��a�64�(n��"��t�A���$&���̹J凗���n��sq~�p�L6��8l��K�����Rڹ��2tԽ{"���V�5�y�PG] p��%P��*�]��_�tyvb%e�l2,�4�nz�J�H�����O�Ɂ�y���BS�lt{���{�W
�#�()�=B��!����k��7�	� ��϶���a^�ߓ��:��!���`[�k�o���'�㊵LÞh�j���
_u�f�	�fF����"��!dB_��X�m��M��>�i�ݲ&l�1�^�I�X}�2�2%��U:r�����'w�om}n�z��D��;�e�M��U@@s _d����͏+)�wJv������3�i� S����,�͖)��5�{��\b��*(��Sv�@��&���%�ߕ."@�.9�4.� ����I��TS�7f�v��&��xp�7��w�!�5L���Y6�O� ^��/tH]��ur�q��0ff�"�f��n��h��.x��W/�����I�>]H�TM�Z�IZ������O��nMD�8��n��K#���(w��� ��t�z�|� ���ľ��U��/m�;P�=��_���|���2�w��b���+�i�v_L���'<V��9������]�!��x��n��T�5��l�G�z��c�_���y�w�������|�}�,��!���F�L?}l��;��=c���Q��LS��W���^2�6'�M\�F(�t3A���\Վƀ?|�S���p͈D�����lI$��_������ܞ�ʌ�ݮ�#�b2�ko��{��I�қ��E��Cc�'s��n�m��`��C���I{��[r$؆g���΍Nik*f�Pg�2�g\�Ūu�x��2Ew��֎�������wԟ��V����5���nh�U���ů����ly9i�����[[&is_�g�*Wn�)��ˑ��Y��8o�g��:��Ԫ������7	=��-������f��8�����i�g���#�ә��E��F'��^~��d� 3���D�(�WTaBf-���;t�+;�x�V?Ih�����AsL�s��ڥ�/��YF^ޛ�&E�2��`��#�ڣ�o�2� �0nԔ]�U�9���k9F5�^ǚ��6[V�
�fU#�-ON_#��thY��P�EB�S�J�����dN�J�ч���=����"���Z����R���2���a�<����'��$:����bA1F+Wu��n��h;_M?�>�u%�����/ q�U��Yr�%�r��OZwȐ�#2_��C�4�3�F�[ /��E���{�wW�����F�Kx'y*�^�;sn� ]v즶\�go�	�+z�٥k���`=����_���!��N�S��{��/&�����[oR�z�.g�t��mp,���*ն��$=aA�i�wz�p�ra}G�p+=�r�V�;��V�8s��%�Ǜ��d� aS}W��m]���d�1g�;-�s��n����rH������n�PHt���`���['�nW<p����8R3A�������������4]��[i<g���T�����w�3����[11�d�}��mϒ����=5cg�2�g��*/7��$v)���"�B8\�b�+�txl�H�\�j��^�j*�]�h��eC.�� �2�Or!���f_�\�"�h�r�?Xa�����i�]�X��\/9 ���3��,
��R�<v"���a��kJ�x�&��5�UT�
ǹ��9�cQ�dݥ2��D�K��	�h�d�;���	^��KVk��>����hIx#�a:����)�m7��{-��+m!u���c�Au�		���,Nɪ�@J�`s�y9�g[��lV:�H���qj7��#���,6i��w/�*�1oU���缑�?H����x�& uK�ɗj�+?�Qƫ���=�V`�]-´N�K`�����p�6Z������	�PD��D�Z���d#-���c��eco���hM U�𬻊G�c!"B��=�_`i����xH�X���^.i:��2����*C~D�F��MO[��3@z��I������kݬ�������Y�t�>)�
ͳ����t��U�YVȭ���ο��O�>�ok�ǟ����S}U$}���`f\��s���"���[��^�8�Œ��%���eKN��l����"8�V}��Z�14e�K6���"�i&��E�<�	�6;%X&(�/Ye�4��th�P�����µ"Y��DI�p���������=z���g=n���刴hgo�5���K���9�[�9�-s��Y��P�~��"S[��cN�kI}��	R�)gU_��,^xlw^	t�T��;��_3꛳{$��:@ċ��r�{����mz6}];�6���#���5ԈW�7���4H��D'�A�=��~��&��M�T��l�4�/�~����T**�~{Xd�!�z���MR�h�k��\���	ګK�ު��*,�/b��(��'�.�b�Uz�����l�	Z���;�=U��`[?`�]8$�u�}����Bz�9��
;����})O�C�]5���5�1u7n�+�;No���>��tb떣̿��C�V�S?��6���q�Ր�� ���}r���Mኼ'q����yЄ�.��n<�6�?~,WcI���a|t��xw�]<i�Tl�(.�	4:�@�`w�v���p��=��m�r����O|��k�1>�����ȁd±E����i��@�Z��HU�ܲw�D�swγ�0�'/�uו0���s1�ʌ�>?�[m�,���	�jeM��wT��$-�G뮪×ɏq�o�
}~���0_�]���;[Kw~��V�N����%�Ծ�O'���v�d5�����R��l7'�E7�?�z�M�wG�N�В��ho���0���5�x�e����΁]c��EHºɛ�k�	���Yp��o�I�����6��ͼr2I�#�D{e�ޖr:�j�B蜜�N�i�#{��o�:���v�q� ���y������|�`W磴�U�%�?6�.���WR���C37�����sA{\@�lmR�@´+�a�?��0oVDk��.P�\�[M=K�hY����xix��y�H�R�h��s�>x�LI�f���Q�V�;h��J,@Ih��בx2�.�9JJ�j����?��G�~��2蟲y�<%�䔅/	��am��!����S��c�U�w�n�.p�\8D4�G���k�� ?������*e&�e7���_�Hz�����b�\+V�.��=UE���(������c������X�;�L�^7�|E�X�i�6���8Qf;t2(�[�T�2%2��(��w>|:ڞ��]5xZ@�� I��X-��T�����R�Ʉr���gLg���|��BW�ܪ���cP��	m��'I^y���bP&K@�t0��:����Xh�����F��ٌX�p>9�q��c�j�j�_Kŧ�u�����Kz��f�{M���'9�b���̹b�2Z'��3�:��I)�,����cE�0�-�:	.'b�`$�ѺqiZ��	\tZ{�0�r��,��Y	�+K!ǂ��L��V�%#���(§|��eo�sV�����������3��[����5���br��c����Hi4`�ד��!Z�K�%<���E�Zc=:9���}�h�c��	�l� gv��Y�e���6��-3����'���bRg8VE:���az)�����i*���z�1�:~B�)���N�6��,�i����iOc��Ͼ��E�]�w��X �qy���R:q�� k��f�0�ܣ��Xsϔ	�n�}1�����a����K���� �.K�tզ��v�۪��3dŤiK�a��ǥ%����a�5����k� 9����0�p�[L���-	@��O���2�)��1rG��a� ҂��~��
�U�'���un9B�%I��٠^K��6���÷:�	7ϖ��:�u���o<��nV��ô6k�)V>�i%�?�m�W҈�V]��ꔘu|��B'z���s�D�en�q'D�Bn���83�_���z�,��S��=�������s��sb)�M�*�x�)�E>a;�?����NU@0}&}d��.���S|�kί��
�5=�"!rv����j�<7#��x�#�D�o����7�ky��y~����rm�����x�|:R��?��Oe~r�� �I"%�2���Nx4�ѥ6DDFz��I�\����ܜg.qK!�
��3���lМ�t
���(����p��}�qbz��W��-ۛ�C���W(^t7�a%ÒW��@uC� �jo��ѐBB��4f�ƽ�����#����v�#��w�,L�֠q�{���	8AB�&�G�kl8LT���Jp�O �x�\U?�*/bK-ʪ���cD�G�|�{2����:� ��s.^�ȏ������	��m��J��*�!�S5{\7<,���zb�;<��<�0L�� ���?u�ܼ<�G��W� ��FD�8)U[��h@����۳�_v���/� T�./�$�h �z����#�?�P.�_M��]�#M�2dq�N]��{T�5��|�?Ȥ�^V[^+a"��*B�l{���ح���{�x{ ;���=�B��T��c(-����Ӿ�~	�Im<��h�q	�
Z;�L=2�be͜X�PyS]��d��!߳o�	��B�29S��𥇩[9VZ�'ۛ�I��ԯ̬�'�#"�.�k]F�8v+>�1! =l�oW˴�;Æ�G��3Omv�]EC>P��kC�xKUǠ0��x�sNZk�*����+&>3U���E�K��6�+ˑ�����p�
a����Y/�uWk������d	wqaB���AO)1�*Ջ��}�1��Ȕ�x�66�`�� w>/�I�����y��T�"XR���^e�����gJ�p���U4}L�C���8�͝�q�]	�Ұ��ؘ(�?FX?��~hV�>8Ь�@�0��A������T]W�-0��K2�� ���pA	(�����כ�F����ן��lV@��-�\��N�:>PYI#_��[��sjo�.fj�i3�Ġ���ZHPGw?zt�d ���\S��:�:*彍��۫���i$l,J�%�a�_�)B�Qf!�o�KQ�m�~0Q ��Z��DS@������!�B6��2%���+��ª�\�T:sk`ux���l�Cm�8nW����q^�b���$@Z #9��1�Yۜ���^"�پ����1��R�&W@�j~��E�M���f��<z����ˁ��h����򍊑��sɓ����א�!�ֈ����������;d���rD�-�h�$��!�l__^3r��0��z(�ʇ��>4k[�9����E��d� <br{�������2�2�TIj�Wx���V.T�r�X]t���M��<������^odߞ�~쐃|�,=�^��A�Xn�{�+#+��S��#��q@u�#��� #��A+��� 1�O#Em�W�x���t\ĈUFL����X:FX�1��D�Jq�H�FuU2ti��%�V_H�]=z���+b.���n*ׅ���8�9��P�_��O@b&4��:�+̭4�&��c�U ��E q����N]9T�m��4�Qv��UC�j�դ�!kfY�Qx�;'18�0�)^��len4��>��&�]���s#���p(7�H]�r�1m�I��Ğ�z�3b�M9�(�Պ��A_����5"VWwـ�%s��x���ݹ�Z��-����F��"_.�#�NxpЈ�x[v�B!'�yp1Nl�>hJU��}윒R�K^�����D�s����q�c��qo��-+���T/_��m���֌Nc�B�����mBL��%c�AF� �������|��^
�U,r�����(\ m���!{ӏ������'O9X�����]�z���ݙg��{|����$�I�S��D�� �a�ནGK��'��-��3���8_yEp��3�/��q��Bg-�9KL,��>�O�T�l�+���g��l)g�$U�}��rL@�F~L%�M�{�b���=�C!jo�����Z���1�=;��I�1{%��;*�����钆"4E�\T�=s?6���t�>m3\�sG"2稛� ��~�3�<o�"�ڷH���ܸ�� ڊ�MG5���������������$
�+^�	M��k��Ȥ�3xKnߐ�@1�Ft���{.���W'��B�Vʧ].���Q��j�ԯ�8*��YAn��}m�AG�1I�����Wށ�a�^M>3%%pJ��2�;�B�ǰ4��JjS�b��eѩ��]K"F|6Tq�s���k{�xо���7��?YI�& ��/�'ܐ�2-��ۺ��[	�,{�mݛ�>�`���%��e^;��K��|��e����&33"V����~k��x}9�͵}�m�H*��lHP���ݦ��؍L;�Ħ��[���ޝ0�Z3��S�Dco	����Ġc��DG��u]��J�V��I<����jK�^uM��+(�G�E���K?2��qǸEFK��և	(pp�g�\�R��\�8�80v�]��[��HRp�~�E�������ڲ�C��q�3�GZ����)�秺�y�:C5��"'>8���EM��YM0 V%c���ʭ�����k�����DSE����j�"�va���w<�-��.�>�+���^�>�o�1�k^�����GjG��l��6� �6zQ}#�F�X��}����T�z������"_Dk�CK�v�q�6_����F�F\��s21o�d7�]xڔYP�#���1�՟1D���]Q9�U���c֌⡽8^��9��(����\/��s�����0���a9���Ps����r������U�ZA0��o�ോ�������|�	������q�v:鯸8*]�2��Q3����*=Bp;>Zb���͂NM|����MXn�6,�<�_JK6$��b�d��w'%8��Ob �?��\���}�d���8�A�=�,��T�l� �iۛ���7g�k�˭��o���"+qe�����Q���~y�SH%8��"�]�X���&'#m����B��_�+�\�G-9�0��>�$�9�3u6���k��|u93](�/���;�p<�@�eT]��]�*��?;�g�<-^��I;@�rwr@��M�(��X�[�E�F�SVT]�m�v��]/�$P���D��5J3]{9�5롋�ѾV3��*�J��{=�~�i�B���u�7r vt��_��n�H��O9V��̩�f�݆�Sۣ��ec[�A�!?W��LꋖӄP�z�Auz0/{�9JC�8"b�9�6>ի�3���w\bG��m\K�	�}P��?�t�f�;O�N�F����� x�v�ڥ5�`�Rz����+@K]gJ:����4��&��I�_ A.s�{6&�!&��-�Ȕ��d��i��#͛.�-���&�f�� ��_}a�3h����wE�,�3j�d;)S��|�&W:c�T5���1�̳Z{�š�ʛ��/�"���e��E־K�(��F���J7Jl �ʈKf�t	^��o�B������ �yt/�Z�C���R�Γ�h��نF�ˋ�6�`g>:w��i��o,*���N�*�*`ǰ�Q��` '_���������{���	#CN5�>=�N�ex�\�7j�}�AD�:}ѷ�+�2�%We�7Bqى�RW�]W*M�(φ\��oC��������=wƉc�X+�fbZ�z�b����ȓK���ס�N�Ԁ�uM�˘e�G���l̷?�U�mL�����y�Z�L���-�؏�BV%3�*�ѹ�a����u�0q�0ޟ�<�a���˄�/���@�#2/�8�X�^�p�0)�t���y�yq�`��9dF�R��3�ڟ���	��=�ʀ�AK���6�@�E�9����Aӱ/����l(��ᢙ�d�:�\`>	o�A�U�V$Ҕo���tj����g2���qT�h��:�z'��l�fFd -&�y
R\�8e�?�9
J�]�4����o��W��#r�>L�S������5��0D皼�S�	s�Bk	��Bw6�v`��B��c����s��%����}}��lzp)���b$a��5d�v����Rz��Dv���O�?�3u��Frf6�kFx�l0-�*�'���$���znӇ %�^�ɺ�[(C�o�����i�h��c�{��iזu>���?:�6�z�"g:�p.\���=F������ȉ��"������ƭ��}��;�<��"�)7@(բ�$����@*V��m74ᓅ{=���I��@�����3QC�*)�مU��G�_c%�����1~.�yJ���U�?�͑���wE��-��8-����yR�j.���.������5�UR{�SbG���l��fޜ��ߣo+~n]ٶ���l��qYP��w�;���o�W�x=r��*�%��J@�C�?�𧅶�caj���!֒#����i��-\e~q��Δ���MV-QP��;ϻ_4�Y�-V����A3Ci��Xi�0�E_���|����Y�U�
��@7$�AD��j;�lO$��=�%�?�M.��ɑX
RD����^z�32��J�77?2�8ެ��R�.��PC����֤(q)옘<_f���r����].l���Tg	��x��I)T�K�y�M& ��Q����VBi�x॒ޘ�N�k�/�Q釿�N�C����75������X��](�;���<�Vn�v�?�;�ٝzWәs��������'"Ld�;�Y,�l���ˉd��\�`% U�Br���;�4��`O��#��Yg5H��Zu�"2S�7v`�E��΂�A10`Mj����"uG2����j��{��%v[��j;�g }���?;H�=��0��j7�J��������?\~ɢ(5����r�ٓ��4��<�
V��Rɾ�=����NZ��.2��lh���]N�!�����C:H���$i21s��}4Z}|G�_ܲ�]����?Mg�i�N.��נ{n5@��A����ILu�!�+;8����3ˎ���#�'���A�N�.W�Ճgly��2Ơ;�u��|v�H G��ʥ���,X�1\���2��}��	�$Sx�v�͹ef�8}eզ$p�r- �嶷�����s9�^/�9�N*�����A���x
?�~�f�x�V`n3y����+���ǣ�ڮ/_���F����^�������k�ǩ���;U'�(�{{�D}����n��C���M,�:/J�V!�@�h�i��9OY?��;�����O��'��2�8i����'��+�����L���mU���+q�'Og�8��%v���Qe�8�pK�ᬛ=�m4�����|N	m���ԋB�Fb����*��f�X,������x���8ƙ��u��U�W���f'�JG�:�G�*���F��2u�F���a���芔̬��}\�MnƲ�
�Ik��ݶx��Q�[��d^�|b��;����I;z-���2�ti��sѱ��p����0��6���l��)�A��>:��ѳj�n�fC��6�~vzi��KH<��[of��R�j3j�h��Q�Xčn���L8�ǔ�BaX[��;ϐY
�]�s�BgF��r�<Lnf�p!3�<Q�z2�mJ%{?QJ�Q�k	U+�vs�C����Ǵg��%z��:����M߲�2#�`A�L����$횑/���ma�@?��ɑ����!ɪ�r+9�0jKOUEl��Ą�^|�5�؄
p�;��|�����)V�Pe����[����x���d��O��x��b��N�R���ﲈ���P'G�a���f����	5��V�����+^q�*���tu�� �ϻ/}�ۺ�D�����nNk��1�jp	��Ț$_��i��y�n���zl�D��_1�r�ܲYT��%�e(9K��^ed����x ?w��ӽ�t�^���	�u/6�C�DCܻ6��Xz�q��ڼ����,�đqs�=|$��҈�[��W���W�k�|��t8�+� �)q�E��g\iu3��e�����!���F����7�7?�O��DU�jW ��J?�M��>�
"zHlt'�Can�
_@�4�IA!W#�9�\to�,r�+N���m�����P���'����6U�(C�10��q����%$v�Z�k����?pIv�|�g肃�`�3�q`;�c9e QQ�9n��׍]�89�o�F&ȩ^7��a��,�Dј٠�jP������*s��k�-\:�F��Vz+] [�-k��!�9]��5�||g�=�������ug/��=��`���Dr���m�׳��r�L3A��Y�� NW���T��MP�����Y��K������@�c�j��h�����ч��ϱ�qhel�ոV�J����;�
�,2g���z?���R�m�����d���| �tj�Afr 4iz1й�b|�9��H9
Ci�9X�'�[��"Hrʁ�D)��[���'ֿ�{��EN�s�#�nmy���͐U��G�>����� X�s�)�����>�@�jYf�c��؃B׭��*5�LP{�j� s�	j-��j�Yf/�� J�Y����>�^����V�Qбi��_��C����[��8	 �V��0)��W4gG�|����v�Y5����.�K���4����075�x�yn����M=�{��G�
*�HIa�/Z-"� ���VОY�Ym�LS� ������Qc1:����b_�����N��i�	(�<��J`�Xs���l��+��lk͏;�,�T�u���T �W~�S)Ӵ n{�����y��W���m���A�nṕ&��
�����ʀ����Q��*
W%���5�TRD������(HHw1�PC)"��9��s��{?�?�E�<g��Z{?�9�Q���m�i�3-�/����p!����ᾲ�!��Mԫ��;fq��N�?�1�˙%/���z0�;���д]2}��ήH���8�۳�^[�xWAK����ٟ�:�d��'gC�IX�Oq]��@���P/���~��Cw��<��j@r?}���qI�U0JG�z7*�u�8��a��Q<�I�\�r�3��"��TIG���%`�^Z������f��G��'r�;����~�u�+�O�v��g<"no�P�QC�����P�KLDx��F�W��Z�-w��ɻc�����d8�����v-":���aj4��Z.���?�U:H{]�S���&޶(�����3.�\a3��>���N��$.��a/z6�t5�z�EN�XU��&aY3�tC/}�_�9�+����)F�uW��sU���𹃓�ZanE��	�Z]��y�0���� �=<"%�Zk�����Q���Q=.�h����,��Ŀ��?�:��g?��� 
�-���Z7�H[�C��>���<�2�D���d�
�#/�ӸS��u�W��ˤ�T�q�G��$Ao�z6G\md#B#�6�l&S�T�-Z��A��`V�WD��+�3���[�.�y�X�#�Hl�"��v����"�8�q�"z��jk?��~�.�f�f~P��-�*y8BY����m�E��(?�L�	%��y��%��d���s��]:���CkS �v��c!�����rn����gF��2E�J��5s�g2�!Wk��A8���뗿�'�^���=�8	\��.�|���F�S��u�֍\�����,�UfE���&�a����Y�X)�v����_$h��w�r��� �-�u��{��Е��ɱ!��~Gn]2)�pټ�]b�Йi���q>��Q���UN�	Ug�ɱ�3���nP����}�(r[��9����¶tBx�������H�P�� |�#��h�<9+P�l����(]���M��6<�&���r�R�8+��cĽ���<��q_�"B�@��KMOO�5�+����KX���ݜ����,xG����"xZ?�_�v�����P�1�L��'t�n���G
aM��(O���q��\�����z�6#��������f~�-q����'R�G�w���3�`��0!I��� �����5���~�)��y��ێ	�Z^#�E˸��%�_��k�x�B�̗��C>T�~�rogk6��������ݭ��ǅ��Z�yp��G"[�i��0)�(%�4��ZB�]I�;jz&]�5	���m*�l$���ź��{����і��0�����i��H��?����@Ka;���Z�$��<p�V�<�������>q2 �J��`2�.���N-d��ҥ�t���������.~��uQ6��G�Q~ 7O|���7ż�h�:0$_��]1�t�`��w��_	����Ec����g�3��[*Ą�fb�Ib��O���(�z�qe�B7��1���1���!��D 3�a�������/�Ϸ�O��a��r�N�/waYt2}�¬��(v�	� o�Ϳ�r�Hl~��dQ\\ njA�����2l�0z4�р�y��_P��c����(���,��Wի�c��kss`�2�����K�$y�!^�����|":E�n�>�b��g�>=1:x#ۥ �ـ���x�<IIY�Ŷ��-8�PԻ�ט��.
9��RN }�)ͩ&1��F���uօ��n�����1u�b��q迌~�����h=�u�i=��,���OȢ'�Ѳ�>+��=��Y�x�ey��I�7;Vz�l��t%=����Q���|L-F�%�:~�H,�[��%�K㤃��?=̀O����\�]'}�5�����nzL\m�Q���=�0��Q��-5w1X�b5Y��ʶgpi?C���
z?��I}�g��_�;{� ���w����Sa>�B K�s�oPW�=͊~��CL{g�m��~AC=�}/�f�����np���i�5-4}|Q��pG�g�d�jZs^��ۤS=?��أ�+�mԨ��):L9�~�>:W��_��	$�}�WP܍|`zu��s�%.Vc�Lt~���lH�K���[a��Za������l#�qOJ׏��cdl��6p�
��l6����V=���dE`kq�W�v+���F��ɗ)/��-��W:�ˢ>Ua]}�=��߈����. ����D�G�Z��P�Ѯ���dMv���[=M���3����@��g%���~��Z���{ַq)(Z��
h�#����|��R=�k�J��(���*��d&fR��}������a{�8�5���R�x}�%��˸)��=�×PT�<��?�F7�C���S^B�*ب31%��"�i����Ti��J�c�nw�:�1c�� ����~�	bt�7�M��,���z,�7셁��3c
 )���3�|�������֕S��XG���2���8�:�L' �Vވq���#��8c��ɋ^ױ*Y h#�@�K����c4/\L/`��~~�@*d]'h�V�������@��b�ź��iS�^�N��z��6�̄��I�K�l;�_湀*3[Wvc�b�:%��*Mu����gg�C�T��s�|ڨ�uN��1ʣkG.!�'����}b䌇�\�f��I��sZ�ɧ��U�{$�a�͕�R'����_��nڹ2��~���ie�;�7<� ��!�0��Ԏ�*S��-��!��8n@�>��R�	��gip�+�4���N� �o�3��c�=���{8y�h*���*������e߿�d� ��K@��KF�r2��qE�(���f��J�P��&������#t\Z�}��Q��[�jx	+�AYu}�m
��;�Jd4�S��Y�:�8���>|� 4L:�4�y&V��y7K�A�F���Y��_�q٫����-uI��uLr��=FJC��7�����P�u(��7A��j���Z����м��!V�m^Ȁ� �F�ٳݎ4���~V��Eb3��x+}ǎ�A�=��_�/L�(kӻhxX�p�'��F�1��3<'c*��7�|�1��*�+��;�l�˿�}Ҹ��H�7�Uă���h?�i��gû)ᕅ�\���Yz�ߛ��t�� 7��qp<��VK�]tk�G���A�x�K_nR[,;�y�a��!�� ;��uȭ�S�!��]��ǁN�ue ���9 �ЏM�_�w����~Z�U�F��E�R¼�$�|4]�l�)��hV��cѪ|��O�j��x���Wl��;�o� 3�M��~�:�}���^�����0չ��vs����=�̈́��0f}�*�<q5�[1�-�YFUd@٬���ˆlʌ�Μ���U�^��.ܼ�� ���yȳ����	�y���'�1�}\���V?9�p6wqi}����aw�+_1�j�J֧�n��UU!�����<�ɧ�v����FW@Lf�G<��Ak{9�!�^�� Z&����g�P����<�zk�(o�ӿ��3K���
�����Y�^��Ex�������
��q)Cݞ%_l��X h=,��	�h��5���7 s��!q�l��v�x 5+T\e��c)���J<*��E6���z��\he~�V�X�H7�$y(�����Ou}1�΅x(�*���ڜ�Ax9и�4�����5���O�
q�8�"%�m2�~��'�om�M�ߍv�_}ոg%��o�3U�m}?�Z Z�X��

o�w!��� ���Ei�@A@`�������_9����ˎ�&z��5��)W���G�8G
�r���_��᥁<�:�um�� 5������Φ�y	��)RB�~�����f���ӟ�\xs&^�����1�A߉^����"�N/K웰��2���Ԋ�O�5���y�tqyM�5�S[9�=�N��٭�tm���h���2NK�~�����8��ׯ��.9N�i�#ݥ5+VK�7:�ê�`p}iw:��i����8���B�K=�5����
��}�I`%�C�
��.+洈[u�zJufi 9����j���R�槰Ӷ�|����Kz6�e�"5��X�)��X�zm�1�F7��|V�A�R�NZ��g@�Hf@5`�l�3_E����3S�O�hٱ��}�[���=�4?�UU� �Nf<�mVU��|��������т��J��ZW����Hmb�A��y���)Ν8a<�4�5�Z�iH[ɦ7 @�K��	�����q��!&���w�r^]p�|8����������'��p v�c|������W��6x�_���_M�Y�TN��g��k��RX���$�{v;Тa�u�{pH�G\���U�m��a�ݴҤO�y�׾��s'�䔥B45�Ϛ���<I �J�� U�
��0��x}읏kzdh|`drfƷʶf����½� 3�Xx�
8l�>zY����t�����@��z�3N�A����Y�{nFt��@bFU` SR?�1d���;��Z�!8��p�?̐���5��,��j��7��k=�d�/~��� n�RA�����*�������>`r0�lTQN4��xb��p�� ��z��k/OJ�Q:�Q=>=�v���i8@�K�E7��ی�..a�R�)e[R��B(�1�����)�����bk�\��_����*�+��61t���1�e�%� ��x+C��`t�������y2Ӹ{�R{�'����.1�扰�����I��~$3���2��]��K��s�Bzo4���ח��w�P��|Hb����6v�Hd���#��0���f��|x��'ʫKirc��۷N��e5s ��m7�aI<�'���$�9I�9�ҺW糺�`O�քJ.��~�x6�w���g�����8_Z,��ޢ ��y@�!���v��(.��7�|0ٳ�����t3*@n(�Eg�)ݱ�j{�׷�Ք�śI�e ��h.[��?��A^{|Z2�c-��I#��[Req��t���EP�<����d�>�jF�
�^iz8�,�,Z���NΉ3��ss�D̥�ENW�W�ͽ�~x�!��ؘM���a��䓎uCQ���ğ�H�|�h�K9��ٵ*͖���� �*��ݘ��*��=9�mѯ��[YMD1�a��?����D�7u���ݞ�g	:��)ҳ�d]�˼������\�a(�ߐ���Eb��$:y���ɟ3��dӃ6� �@��?"B�iXu0!��Y��$��l��Ѐ.T�.z�ELK���E����B߶�8��4!�̄��ՐCn�Oݗ�	'�9���r9�wȽ�=��|ݎ�}������
���i����[����j�cyx��-�m��e�I�j������a�
/Wg4j���8��8K!2g`�.-D5-���ժ4�T��5�[�&)��@�>ݎ�ji��m�/t���5G:H=�����pog�7��϶p�&4�H��V_X����s�>�~���I$!��l�YS� 2u�`�����v5~�?}0:��j��d��]�W�u51�w�����쌄�"�b�y<�H�Rey�_�1Q��q�dɓ)�#�3yfx�6#"��r5+t��̱��f.|�o��7�a�O�GRނ���V7|��Y?�u�$����]�g6E)gD�k�̿�u��9Ȣ���ޥ�+^W�f��I6$d�XN�e�B�,��g_P�Ud�{�����w��g��x��j��t(,�Yh����o_���k��mg��.ГB����E���}zF��`��<p��-���I��2iG�����L8��Y�¨ƽ\Y���4���c��qn���p���F���u�_qG�厀Yz����L��8h��MV8JD��1��.���=����Y����>_�����p�Z��wN�'��^�tΧ]�BcH��52-�%	̰z���f�Ftʕ m�ĳGj&�1J��R��g�;-	��p~h臟�?}j� G;��E���=bae>x�\^'PX�@�c����l�ŷZ�gǇ�<��hZ��e�)E�V�<�ϑٯ/�J�|�P��*�����'��ߧ!z�ٳ���R���:��)�o[<��~}�VT���ı�0�0���OIO���'�R����6��V��E����9<Ulx<W�����~T�f�fP��{��X�����%`{Y��\m�X�0��MNw��`A�@#`�f^݊xм=�4�hXʆ�ݔ�S�Ef�������&��ieIK�%�u���K�{��������Op٬�t��:�RaJ��hN�����Y�A˳���~&s�UE��DGOm��E��71���A��R!�r�g?�<OU�*fg�Kʫ��^�1���5�v�V��Bx����l����c��^�P�?���`��o��:M_�0r�l9�*B�Qz���ķ�(P���8����j%�~V%�|��6���zh3��b�ga�I�;�rt.Y�Tw{��q�|C���(�$��Y� _X�A��;|��M��v�u}Tߜ�q!#!�Yd=%�l?���kT.�e�x�I˨�"2���=�]�B�S�N�K7j{~��R�Js��{��������:S��e��iDK�#c)�͞����*7����Q�6�#1�HINFx:,$�9�.���	�j`�gM΀S�YF���u�oxQ~1���[QqA꾜'��=�O��͍k�On k%JNu<���*WK��M��c���.��(�cM������0���^Q-GR�Rv핃}l� �J}�^d�U4�M��A�P�R}�P(�dF�e��.��C�Т�äXV�����Y�L-��Mx�s'��'!Q�t�]E�<{{��GxN�^��BN6Q4�\g��,���1��gg�lrP��=>�,	�<xP�RWǐ�Sq�%yg~������x�y�,*��iD��b8��<�,�(���H�nL�)���蹞��K�̅�BĽ����k&�/��8`Rh��N��gN��ͻR�u�\K=��:R�x��̼<�P��#�^&����>$ �HG`p���/}Y��r���#H]�$ [w!�Y�%#�������0�
 �);����C��1�#�ao�
�~��.2%���n]�\�2h>�Ax{��n��4TU����fL����=;��o[�^b)�VE�	a��������whʹb+��f3�	M�f��$LBu�,yRBL"@�I<7���/Y�/�=en#i�'竉�~D��877�]�M+͖��;�!H��q�:���[{_�U�!��q��!��iE86���?�ʮड़.ʔ��1������!6|��$;<gNV��x[D]�@�fy�I;�����W(�$}ヨ��ȿ5`��+J�r�����qJ��>����\���7��B���L%18�f�%�������l��ɭ ��e:�.�?k;�^_�a�d0�]�5Y>���i_�B�j��IGl�t���v���p�-��Kv�(�j�_ɷ�·!�|Z�/�+�^�HX�L�W+��c�&��Ck�LV�:�Ph�u���@���ډ��T��F�D	8��
���˳J�����>��o{FnǬ�ȩ��*�y���uʓ�*���������~
X��p_�Jڻ�nc3��df��[K�ҰV���G�*�2^��S���cu��b��4�q�����@&U�AwK9��S�<��l�v�7^k�>լ&�j���e��.y}���K�)̎�����z�K����B:t?R"W����T�S�Y��aqB6p�f�u� �E��ܓ`��%�d����������S�i5� %5K��t��{b��꾂�s
z�1�cG9�G�H���u�P:�ILd�^/��+}�&�w�⑴�����76Ny���_�G�D"
���{cA�����)JHe�ښE��E�Nn��4k�7v|(r�~i:
A����͝¸a�E>�U�z�O�)]��f���d�(3C��F�OAu�Hʀl�ա��1�0����!�ooh������VO��rs���d�ʢ���:(��&�'J/�gr�c������Q�*-����H���|<}%$���>��PQC1i�<����*k����[�{	����g�d��1�C��\�*����M���S6�P��b\^���9�>�~�c�̫�G�Ê}�1��W�2��OB���:D��S�=�zt"�$�{w����.7~�H#��O��x�_��kУ�S��ګ��ԓ�&���L� #88 �|��:߿����'�#tdƤ��tb##7���^�9F�ȩ�h��'?A�Á�Y�3� �� m��ϒC�`h��^J�+a,7.7�[�6=���
_�r�1�1��6�a��li>���~kb��͛j�TV�ʹ�i�nl������̥�H�(\�k `�1���/�2ۊ��?�ؕ��=ü�Y�*]I����X�V��<<��o:�=R��ɥ �w��qm:�ž7CD�Go���yS�`]"�Uޚ�}^����5F�R��y�-��}9�`�����M��#;p��\9\��zz\�6���p5/1Lȉ��gNDjB�C�G5E^95�䔁����q��TW��dC�32Gnf0Hʎ�?,"��.��c��44�%���SG��g�'��_;V��*�g�$�>��>��������(U?e"�T�'
M�ì�@�B7�u-�;dVR��?��&�m���>̴�=�yɒc�V�幋phy<�>�����g�+��Q~�K�f�2�l!Ʋ����bl�ni�Rv����>A�:EVh���n��h�[�܍*;�C��h����Ͼ/r����TP�{T^@���I��:`]\��?�P�
eT�G�U�~�����L��~�.��! �TК���w_�S�ʴ�J6%+{��=�Lc���"g��=	��; 2N�O6}�N9Y�I�e?�����AhFG0��9�]dd�ڜ�z��n	�*r�}Cc)����R#��_������KӸ>��4泆����*���PA$Yި��c�@l�YQ9{J����k� z��US�X]*���b�G���cS&�JΟE�Q7�����(��MB��!&TPM$�>U�ďT��R@Q1"��������'Y%Ś�46�0�-�=����� ���ݓ�g#o=���9X7���Nj۸�O�'�(�'����ě���9\�����o�x���j��b���������5��P`� ���Xz����y�k�&ʵ��)'�Ŭa��ù(ޔD��KN�nT�K햋7�U6FY������s��`D�l,��%1`�R'N����|a3��Z�.�v3WkBg�n�V���%2���]AW���]z���Z.���J�����T�zO��H�����m*��%Ge���@�c��<�,�b��P�a���}��q~� �7���-��MdvJ�/b/e��H ��M�?(Φ������Q����Y]�`��k��p���K{>��;��<+��n�E�pu����>"�$�~�r��p/��I�Y}n�R�B�s��j
W;u�z��X��|�/�����O[2��;U�H�p�����a�V͠ AV�S��}��ۓq㮺jI����+PT�:z&�RC`��qL>a����e�Dx�a/W>2~�_��	��ڳʯy��>c��V�O��H��;ߊ��� $C�bo6� $́�j]�Ǭo�[�Sep��|w����MC�LM�EYػJ'���2u�P�c��⧟I��YY�,ڙ�R�B����u��6U!�����w ���E�|�q�59�!95����L�jj���a�	��w�a�Q��D�W����،��H)9��5	�9[��c1���ъ�.��g -��D0Zs��3�Y�����#JŁN����gWD	A�m^�Ī
�o�Gl�w�=}g��b�ղ�ћ��>ɓTd�U�8�?z�c=�&;"v��������|��O  ��Ж��MFe���}��Ϲ5�T��xiR�cI�:b���cb��J�ԸT���'<����9TP�x��q)���D���o� E��(���*�v�/uw��0���t��p��P����Os�2� �k�
 �U�٪��'GR�(�X�:V��3��ʆ�/��i]��ɏEY�hx6���3���Җ��F٣S����ɏ�B����o��˧̤a����z8�8�;�|����� կ�C��cDB)��yr])� QXu�԰E��?j�$:$�6Vݧ�w�ж��������'��@��4��5h0��
<\s�,�"�=�<�%��{@r4���5�N������H�.�ǐIJ ���.�lһ%?�͵��|��f]��Ĩ�K��8[@�Kq�Yl�%�ɂ!8϶���g�:pF�
��
о�Zw���3�N&ԕ�Mt"�a�r�#�0�P+�ME@�}��Ia=�˚���4ݟ�~�u�A��YG�'=I���@%�+Q�h����,�O�&�B�,ε��#����t���)��������~|h�^J�4���.Bx�MR��!���i�o�<�%;�K���q��d��>�T���,�
�jX4���}|+����5OhAb�񈷥.�@���4�G�B�u�-�
[�ξ���e��c%Ph�����)�T����S��홺Ӕ�/������4���c[��}'���Z�f%�l���\����彵���C9�Ȓ��`�x�c����kc��x�v�/�,��k7Yq=yņ��}S�1��t��C��f��^�o��J+��=��}�g~���T+���?�C�S�a��t��r���&^ۇ��Q�4�u�_�w��f�>ʯ��	V��f3|rJ���d���3�R����a�{�e���9{�E�����ܑo[�@�,�="��걺[D��]�Kk�]�Yt���S��糇v?m��{k�[�A�%f����t����рZfa�iyZ{tX��x�(=y_7�^����y��r�� �V�d�Z�.GIAQ�6C�(勯U���^�g���h\�Ҝ��Pg_�l��4F��mɵ�b��%�����i��jy�aQF����AC� x�I�	�A��U�^>�+�W���P�G&64ꂠ��&���]�����&J��j' �Φ�lreg�!�Ks�Md�Z='�CPK �E�N<��:�٦�`���]�nfc�&ﺥ���|�{Ub�4Q�@���j�%/���v�~bk�A���/��]:�S ��e��4}�B�4,�xJ��û}a��k�����;��j�q���K�5�^�Gw7�ݻ�58��g�w�h4�n�(���-���<K�C;�ˋ.u%5��:E�[���Q��S��1��8썵(�V��7��rg��{uKC�����+f3w��Re�k@_�����oj���)vtZP���w�+@n~��E�5Au�E����]�s2:��|� �e����T�>`Є��t!��L��4o��WT Qrm�h�^V���<�6)�M!����j{ud�u0Kf��bW%���\r��� �@�=�|��M������YC;����G?:���VN����
�r��>}6���XNPY �4���˓����(J]THs�zN��{#�_��w���Um#d�X+��-� �:�v�$Iw��\a�0m��!�]���
���%_y����C	��a`kSF�m�/l�8:��!��9����2�I�������]"�?��"�)����"i�j�M����l���]7S�>�� �r��� �*�] ��_���coaܯ܊eiʟ�,1��Yn�c��3�����gL���R�%���,�z��r��0&� .��<Q�~��@k������y �Z�"o�n�C�yqHŏ���uT%@�n�T��v�G�'?�Ss������N�x�D ��� 7�*�Vg�X��jILt��z���׫F"��aJ�S �T*��yz9�WkC�Y���l�{!K��w6��nv�1��U�R��Z�]Uu�]�^X�I��[)��ݾh~�&�!��#@�so���ԕY��g�Ϻ�5R5�1��]E�l�������H��uH�t�5�=��R�rs^���p�h����T���61����i·K�B������n�Q��,�qҗL�dᰔ718��ۛ��n~�K�o�.`��>�QP�j���J	�6H���m��Gk��߆9ǰ����+i}x��i5+W�"gΧ�TL�	�
�gR5��/�K���/�"�5�(Q��'�������R1p���/�rL$3l[*2jv��$rF)5n����|~��|ﵶ4hx������޻���h�L�P��M+� J�����)1T&���5h�8���a�z�QQ��(rp��Ɵ���I�)Of��F�����ĿIU4g��.������<x�l�x>�s�����/Û�f%eo��}f�'/�E��V@������T9�K~2n��<�th�����H}����ܙ/y�b9e��c�H���s�����0Zꡚ�;N�|��^�L�mh�~�\�'`䢋/l{�ʻ�d�>��N�sPpK4*�3ˎ#��j����G���rɢ�lI�[�����N�đ4d�� :�ڢl��u&��r����� �
�X=�4�Wݜ*ѧ}Bhԭ�� �E��W��0��饡�r7i�k-_G����<����n}Z>��B�0��e�o���p��8��p�'3�J��I���V����+N?�;≭K��p�$�h/7�cs�dvp�N�U���Hb(+I�̙� KC��9����h�R���{8��3G�Ym|�.��,��H�Iz��Y��-�V˭!����꾃���k���#Hp0���P}iJu2����j���/��M���u~_ݖ�\�GLt���?�\ǕL��G(����>/?i�#�5#GRG	�.�Tw�<�螿���R�&]X���r|^T_��&{���hS���3@���f���c��O��R�崤I�)��;���F�'�|�SSB���
^p�Q�p��h���S_��D��;��!�;��s�2!�zߡ��l�;�t����ى���T�V6�p��#|�:Yo����m�>)_kB���k�\X�=!����*��,��ߡ^���	t�֢���kRuu�d 9�������R��w<��o�[j�F�c�����1�P�U릫��`n�<�t"ST��1��`Q���6�L~�R~y*�%����P���&���5�X:�Z�Vqkw��"�S�*�P�{K�!#0�����	���A8����;U泆k��s��)����%`���������oũ������q��ђ�s{rK�F7M�0I�n��vn�4�^���?�ׁl@tFe��+�Ŋ��T��*��>�%�+��n_mn��p��L��ס^u���g�~�-7^Lp�VD|��fM��£��2Ax]�n�e3≜ܲ^��������Rۡ�zzc��v	�;8�w$�&�zɹ�#}<m+H�l%�q����Q�I�����$I�8:pl���>b���ikq@y?�t�Ω�h�i��-�`Һn�d'
#tݩ��fc���HrM�=�1b�l�J��O׻49+�7ŭ��9_�q�&�C�o��+�*YK03�Np�bG.���&\��t+�y��7ۋ�"���PPP�p�����P�._�fc���tݲ�Z0�NK +�բ�����h�(�ԛ�Y�d)VF�hMY���1B�	N&#%mM���(%z^� �`��R+��x���ᄎ����Z��v2�C4�>qs��?�!�~#��ϳm�R�ڰ��/�Wl��V�����9L.p�=(!3�(1d5��6,�>��%�������L9.�o��Fp��s��RdG�$���R�A�d� ۠io����x�\�e�����$��`�ɑ�Z��q��vX$��/ܽ^S���HZ�r�M7{|�>�?$���g��z{��U�a����Ma�5J�yM#/{T�|X5vX�8s�l9׾��F����3���!������|�5��pz��2��˻���G��L���!@� �E���d]�j
F�i\˽Tx�@z?y"#�P'�V�Dr�A�"����ZZK��	��P�Oh�̡�6����s��{�r3��]�㧷��uG�Y��WK�\�C�p��6��)Gb���`w_��)��~`S�D�z�m�l��,�}.�Z?Xqpi�%>2L��6_� ��+KV,#K������o���7�˯Ҫ���n{!����H�ҜU}Bܐ���G�q��],>��F��e������n@��/'��Եg�~4�
������䊥�`�V�u7��
���QF|	?�Ûl���h�����/v�1���ox�6N�<Q��P�s#j�l�|�ܰ)˘�O"Vs�We�f ���Sf�շ�h�r�a�Ks@�3���2�X/#�ܞs==4j��y�4)qimq����	t�w���������p���n7�}��4����=�ᒊ�5	��4�RXZ���h�ެSh6��fʅ�C���;��[t~�Ī.�}���[�AB�JƓ�vG���=�P��F"avq�b��;�u���\"�Y��d���$�l�}sXK:��>Z �bT_b�:窇�F��p��H�?]�_ۋ�}�����G͞nJVX]�Q�/�Zfe�|Z��������+%�M��w�݅�}� B�C�Ն�}	�4=S��r]��C����$��������q��J{�Yb�������Tl�q��\�$V��u����\}5�+�K���uh��+��(U��B�R��Wj-��(�ä@�\FL. 8�vY~��������^����aA8kWH=���� ��t�y����W]?�0.�4]���1�U��Y��
1q���5�g� ����%�Ҹ��8�q�:�����*��^(,_-����p^b�P�e�/C��t���b&��V�kڢ��?��!��L777�iJiq�\���	DV����w�W3��� ﰑa��O,{�I���I�*@O0�~���I��#�7>����Tͨ�h��d��vi�����+���N�֍�%� _��ˠ�Q }S;D^��^)=y��!�%MY�[��Q�Y�)��=�cE�g-��+H\�{.�v�_��˓PZpZ���z����]{�1�����LI�-���]#�fYJ�t�����{[����VM�!@��|�mu�uf>�:Fɏ���ZoZ��+O<�B���E3w	>�1�v�	[	�����K�1����pz��wmyT�F�m�{;B�өׂ'�d-?������i��C�w�i��V�	��N�T�;�$H
J$��cP��3%ˬo�f�\�?]MqyA
���s��-�#��hC0�|KWy����(��#-�Y�� w���)��Q��P�����,��QP���	���YT�,�`���p��;=��?�J�EQu1�
2�E2��Z�2�ֹjR�W]Wm���A3�QZ!�\q/�a�>�HE�2uuX6g�Q���ִ�4r�]PՏ�G�p�qH��4��{?K�� ��T��TQ ����#\z4ׅp�<�Ѡ�����̠$�wV��cy�f�g[����"*I���(�(�>�aj|�gؠ*C���P�,u��_!�^��T�U�͟��?�+&&Z�䚳^9O~����<���`��5y�B_ -<���૨�E^�v�7-%����p��5�,��x�,m�?��	��;��G_b�����ʳ6����4���۽9�%��iCq�,Ν�x�G���$4�Uڸ]D]0ݢ�%z�e#FQR�-��nm��>5Q�rjq"�(�d�P3��ld^~�d#�1�:�9R�c�<.;vjjF��6�{�R�I��aɔE[��8'VBn�
��k�����a�U�#ul�����u��,߰e�M,�����UvO��"×tCk� ���¬��"�;��!K"���:�	c���W�Ĵ�-�:%�HW۽G�0)�����,'�-Rqx	h~
0���I%����k�{8�y]��e��r孲B��K����>/HYZ��DS
C �&�)z�N��l�Zih#�ޏ�U$� ^cmj���TN�'��w T�.y���d괹k<���SSĔ>��L�I�La�I%am4��ު��6�PA�f��K�u�>���pEG���Ϡ�{��H��KI ]�w��;Ǔ��~!���.�lo�3\O�Ͽ3�x*0�������K'�fH��D��	Y�r�S�f��� X�D��:n2W~����=�uBڮz�8x "�V�%G����+K�@�e�x���ͫI��7-H��'�]P0�,���@EkY����7�?��,��0�Qr�����2@7m���n�B����zVm�T)��dQ�M').�k\���;\'��n�[e�fa����,2<A�,uӦY��X!n(o�Pxw߽o#1�����A"P��u�InL\���.�6����ʜ���o?\؅E�
[K�a�'3�������v�289���Y#�����'fI�(C�<����T�#���rԜ"�8 k�����%n���{ޣ��{`�ϱ�]	n��˨c�:ol�2*g���y��}֨=h{֌�"�6w&���2��w>��H���$�k�����c?#��>�����}p���j���找v��-��)�y��-B�QZ��{�X�V�&_��� Y�Y�C��?âx(]mXFr���/{�.R��B)aH�b��rV]�����kT��3��D���[��MU�b��ŉ6�ʱ�|���٧6��׵�����lU��j�a��<<9H޹��ړ��[]��k�K/?�g�W?� �9��<��Rv��u�+k�o�Lx.�X>6��w�5�g9��a%�U2�4�s1�},dZ��:M����&J�E��zlӮbI����7�G�ֳ���7۶�@'ݯ��Ul�?;�ݓ�hl4�"�h~ʝ�4j�q�(Z�q��yXPN���&�!p�}�U���X��ٜ���[�)�/�ӿ���[�ve��������v~^r��C0"I�K�t>�9�����U���i�l�HJ�M�P�����I���dC��zT��@�8@:̭J}���X�c�"չ���o_:7�0"��h�qѶ�:�1f^w�R�i����(!�1:s�5�j��h�)�g��x�c�e��I���Ŏ����h�#Kp�G[ 4��c͡4v!�.:��
����ќ�r�aOs��R1����X�k����\F���v�W��Qr���Ob˷SN��Ngʈf��^��������C߶0a^u1 �6@�;�Y���βJ1�6���5�u���jKCc�	��2�M� ��|���X���(n�s0���0�gi��qE�������t~{z�X�N���U�{�k C�H���4o��Uu�mq�NP��f)p�OdXs�@����E��Η6�F��CK)��*Fџ������=���/ZB��DO��A����}"�{e�	���0D�����=��;3����߻�͚���֜����g?�{�3�[��8@�Ѹ��N�����\;󈈂,��n�}ZA�L}G����:� �~�/`���Wө6�h4�z��Y�K�p!��7�SE�����P����B�٦c0��R�]����D<����j�9O�J��a�蝥8>�iG�t���k��"Ü���ln����AC��M��kdG��L��+��������M'�i�Ñ܊*�OR��i�64���	�.�;q1|͖SV��gM
�ufKi�E)�����\�|ٗ��C��!���My�o��)-_%���w2��N�)r�Q����n�!�I�5v)��O��ۓ%���|췮�ܺ�4R�bm(]�%�ta1;���� �;�{~F�1�v���*���P���g'k���9jAK��jr��l�;�eN[�E�9��9&���x��T�[EiN����РG��b�Hs��-���1�Al�:���Or��L����V�o�l~fx�ὄ�e��UG�����������P��Y�7�������}n����p�����Y5h�?�u.&Ӓ�b,x��A��`��E\&��)ZO�y�_w
6�i�<�� �J,F�9U@Ǚ��A;q�x�j��u���L���3���C)Q�>����=ظ�vE0��ei5�VA2�9b�5a�b��L��
%��A'R&��}iM�h��z@�e��@��@�[�,��#KV;Dd�%+��Ľ�z����t� W�uuUi�y�C=Ck:����sj�vd:-�{4���t�7�p��S�2�R���szM�'0�~��h�j�$�U��&�hA,&��7�,;T /Eq�O�`��k[y���0%`�2�gf���[�_y������w�����v0�\+������ۺ���<̃֠���	Ʃ�U3���Pv�w�Qd�&�E�q���� �Z�� ��"b��L4��@t<��&,���# �ܡ�o�5X���Au�2�-�b�?��P�����¦�W��1�pxXb��ޣ��-�`�BteX�oZQ��Q�87;;G�i*�~���w�ab���b��}���C(`�ؼϕa;iO�O����s!�,J�`c����m�B���Y�� +��?�a�K�Q(Ts���(�����֪m�қ`3A�ȯN�Ϟt�̩Ҧ�&����P]:��X�w�2/ �`��?.d{oH����Q_�Ť���b��q��8m���b�a~�g�3�Je)�
�,��`&�@+�NB�%e}�bu>����_�]|�0-1��K������K#��$�!s�kk��؝���뎏H�/UVZSO�`+�u�n��h�;�-�^�}#6�Lg!_z��^QB��5*!���[&�:f�e�]�%�a�m��.E��C�����|��x��@�DJ�3Gh�}�^�GL�S���WJ��\�[)�<v���&���U���;8`u{մ���c
ω1��6��אs�l����˧B��
xTM���SQ����KS��	�PJay��>�ߟ���q��L4��U�E�\� ��.� ��jqJCy%�c���"mfj�~9��%^w��#�q#�a⹻�.! ���|>�T�U!��mI@Z��Q�|���IB�~o$Z����uQ�ޗ�Fו�MfqsY4���Р�c5�Dw���O*�	E?nb�k���[�{ٗ��7��{��tuU�՘'�ߢ9}��A=�=��Յ;�,"���N�z�@0���λR�u�$����5��h�1{.���Z#��5ź�j���V��z���d�d��++'�,��K9c`�?_��]n俌��Ւ�L�ƝƸ�gu���}c��r*q���f��k�e�u�@[� ��!��S��!՚�T�wT
|�*�;Wx&�.cb�1J�k�>y����f�N��~]ʤ�&�z��հ��P<��i K=�W��{v�{�_5g(9�&�6��a?�˗��|?�kɣ�v��jbQ=�L	��2���׽J�]6a���.��E�v��CP��-��J�v_>�ݢIh����1��0��Ԯ�K���EJ���T��(כg�'4��۝��_���m�"�V��мʆ=f��+��e�ຼ�R���F��"5�K��2�2r}�͸�G��y��E1�S9��˘�T���jR��z�e4�2;G�N]�3'99'���?��gSf����� '���h6�{��t�ϺD�	RIO�i@���CS%.|�M����bL�s|�w����!����s�K�h�I��l��K�}E��H71V>̕��u������E~�(2� 'ac���j�(>�H5���1���OJ�����+�º_^�1��%9���@%;}A>�-7�@ �Z��?3�p�SI��.�n��:Ԕ��*u��H���+O._�<Qo�&�i�����K���>-D��Nr�`�'�V��>ޑ�#��7˖��b���s�ð�����<z%��CΙu'��,yV�b!x,e��+���Vo,�ǳ~Y,K���@��*}�g�( �ȷ*�:�\_��5�>����٦�p��;�[��U<�n3cתE�C��
�ēr%Hn[ոN�/�|�s����E����H��C�USM�lI§%z:_gQB��|B���b)��p������X�[{���3�3Q�U҄���o}�%X�I�L�^�@�l���w�a"#����sU^3����a`;R0!��ٶ�2��+%�5B6�w¬N�4�;<҇���þ�s��-T�+��t����,�%N)�E�O���<�
�ؒd���6�̽��ᶽ��rn�!��:]���W�}�p��6j	5��&��� Bs_�����̃�ً�����|����&쎏�ܼV|z=�>�n^�@:s���mx"���=��U�F�������*�^�,�d��Tȧ�p6sHC�ښ�J�j��c��P��_H7n��Mo�ؐ��m��<�N0�-���()����o�[4HI��Ǌ��L��=Wj�[<|�����	��K� 
�ֽg���æ�tE�R��|������\�o�7�7���}�läRP�0Ffa`*��aǷ<'�H�$��D���}^��@T��Ka�{��t�kBK9���+���`j��JRtm*�<�y��Z��d��uJP0�f�ペ�Ⴍ��L�o)�b��Ht�w3���#x]������dj��԰7lP�&�۞�^�Uu5��}�Q��gi����C��,�V����~�`���xv��;%(q�����Z*���'��:�Mps:wz���	ww��3�kXb��櫎21bJ�w��]&�"��I��VYx�/Kè:v�߾/w��V]��(����뉣o߸\)���*��=�Fɟ�L���.Mؤ���N�Y*����\0��l��P�a�Ob=A��چA��A�<�?ͻ���fU�5_0˷�Ȭ\d��m;(w��|ifc��R3���a�4���4I�K.�Ʌ��݄O�%���q�~� �v�~��ܟL��|�ǜx_����y���L�m��_
By��btN�=¯���� d*��V\5m�n��mS9,)�%�y�alXm2��G0�A�A��b�<ޝ�(��3�/~��� ���J���/`�������uO�T�%*:�E��f��bGEOD����*�B"��7��r�J���\�7P����t�Yk8\W=��ܾ�+����l�r��m�*��ꚟg&>�9�����%&5Iw���RV��b��3z&9X^&t{m2�K$��o���m���ec����r����cD D�����C/���5H��*W4�,!�S�!�Y8yP]}��QV��!�U���%$�w�R���0��-9�$8���)ǰ�����f�ꍹ$�H�����a+��zҫ�s_3J�?�B��==��QJno@K���3��q��̃A��GG�V�j_��;���I�F	l�r�G�М�3���I�Xw ^G��yQvqE�M ��>��T�G���ݕ~;�����Z�Z�^�����'�J��1S�k���Q�Yu�|_иp��d7' H�WT�ڹ��﫪�F��5�d�������6¢��ӵ����<p�\W��|&�5�T*N�v[�b�V\_���O��h�l�O8ܶ- �%t,Zt	�[X+���v�����\?�= �u�(�T������S�4-��~�+^ա��~�����ctO�ſ��lc�z���JJ�L��kEO.v�����#<���u��$���ݚ����O��G�ie_���?�5�|�*��.�{d�[�O0��b���;5H�WH�	1��w�]�'�l�ȷW���kI�0���'�>2Qd�y�����ǒY��y���rD*��<~v�� ����Cd�#ث�f&rb�Y0?�hL�ި�����<f�����?,%n�����ߵ&��-�iAz-M"1%�x��8DV� �m�nJ�F�á����o������N8��f�]�Mk7_R/z��Z{��͕Fx�������b&r��+��U��ǽ�z�ܥ-�'u܉��Vs	˿�MƬ�&�pYl%G1���cJ���L��	����l����W�sR���D������N9J��㬹� ���)��z��=n	r�t6�&|�=�.��n� �ͬw���Z��*�uz�j�"qK�v���M�h��@X�ǽ�׵�o�TV�szZ]R)W�8��,��TWy<��;e8Uz��W':��!�P��0�hgۇ�*R�EI��F�/n��̖Z����K�N0���ğ}�ma��R��at5~$y�7��s��Eq���4��_����.OE�<��8E��YJ�nȣ\�D57�k�W|�h����P��=�J��PV���:Keh�T��6�TS�7 �����/���פ��*��rfPi�L��l��{�^\�	c�2mour�Ѱ���M]I�3B�ϋ&�!?��h#�&!c��e*��OgD�4^�J�����������$�jW��$p�љ�%���ü3�n-��]�mq�IRLUQ�N�<8q�#�̈́���_��_���<~��M
��l��_�C(���7�>�V�0��*?�׷g%re���6������ߍ��3�"��B� }�Hb�����a��Ǒ��z�������EY���&��`��ٖ���}̊:-�LƫyH�`��{C�l�_�׽��e�8�G(�0jSsBto���jk�	D!��=���]��7X���z��9���f?�fw�ɯ�-��B��tƐ���v�ߨ�;��ڪ��IB-�*�I"��AJ�&�r��6������oJ�ZL#�[~�C�/�̕{r{�<�/�|U*���\��'��������j=�@_�����0����ܰ�e.BC
?����H��4i��M��S��X�f�82���̺�6q���>]�v�$�-����X�]�U^�����|��d�z�I�|�}�Uw�����W&	�X�%�w���#6QlˊK�t�[Kƻr�����u��Ԉ�m��F��kZ��t ��E�ʐ_�A�a�AA�7���Ӹ4����~ޑF����a������#7��aߔ�x��z������(�-�tl�7���`���,�b��P���F1慭�b,5�ݳ�>��O�7FڏWV�S���\ZXX�0�#��"*��~��ƙ|��x+���,\Æ�c�K�Z��&׸�jX�]����� �_MԟM2�_��#�u��Xث�ǆK,
�����wO�HmH|���Jw��rf�����oe�}��Ȭ(���xJ�hM�����$J"��aч8�<\�Sؽ��.�9nl1X���@df��o&.���l���{��Pq�6�2����Gx
���n��&�����1(J�0���1Qlu���l:�e(��ak)*���&Q���#_ӁEǂV�?�\��Э��
��9Y�~=�p�l���q^]��~�az������dvT?��,x/!���/��<��1UUcee�v^$*�[��X����j]Xۉ#~-%תJ��I79�պ��Z=�.!�w���K3�Xy���y� ���/��un�Y\���&���X�Y�4E�����cu8�-{�`S9�������Z6S9�����3��S.U}���݉y�	z�^��k�`)��8�
>�ޚ�?��m��~��������@A�k�<�U�5+�1�*�=#D�}���!�,�8�s|�i�D��VC��j�ԞUt����݌����`�^��s�� YOY`;K�pФ�CN&@sAt�%@�5� �;~��DZ�iI;�����Ӻe���g��{�N�S�[^��x�d.��LDkY���M�\��>�������qN���&8>X����V���T@$�٪Ȃ��O�7KJK��Y������
����������1��\�����h���Fգ�v�[S|�J���j�U�����Enf�G@i�d��ԃ�ݽ(��J�^pF9>�L�>�2�eJ�=�<���ka�]�J;l�dK�R�\�Yb!�a� ?Ĺ/__����UӜ<y''ϣ��(v��j�є����^�O� � �)�ég̚��g��Q)_/�m��y�]u�mT�A�ˡ�	bQ�����u{yޞN�|�mS�d���꾋SP|H�0AJ6<̴��Q4'gpP���nj��mL���I�`�=Ɛ�ͣŖvR��"��`Z�n�M�v��od\�fS��0>��<�I'<�����I��� ����#��<(�~=����w[Z蒰���ܳ�a_��9��]ɞ���wr���b���^J�,���l}��z��:1�i+��t9��qdq�5L5��/*rk�ЗdhV���(�d�@�H4XLV��lQZgs
bE����>�}�=�����-��ѿ�F��6 ]�'����?���Nv���~W�tz��֛�}ˋ����'Y6���o�Ȁ�fS����?����s����8��r�غBi���q�B@��@���\�;�n,Ɏr\���W��K7}����,�~���Z˛\m%����g��,�Cwsu����^Y�����9�8pc�N}��żN�-[�r�����L�BE�;y���"�
PX���B$������Q.��6�6��+�zi��.�+˙3�g�+��Y{F�/0�� �Z��"GLt�����_����ln�O�Ξy֯+O%���}��[�>%AQ�����ٱ2��L���MI
pYC�sȻ���Δ�S�m�[O� ;j�bD}����6-_|����`�Jû�ire�
�X�z�eQN�`��c/���=X�)�9��Z#�֤A�����o
���zs+�e���D;�0�t.������'3�49K���+t�Ţt`%�Q���ZO~P �f��k��R
u�u�M�W�i./f��4�+�"5CY>��DۉM�B����4g��G����m &�QVX5$~�~|�ָ�X�y�N�)�L�ԂF���̨��n8g�o��U����1�҆l���<���E�m^8O�^��m�i}#n�ڛ���Z1ڬ�9��:�4B�b�r8�֐�7�ˡGv�sT�-(�U���(l���\�
�'I�UɬoO*��ҭ��q��gU��M�b]v�Ӟ[p~�b�@�r� �C�QK�j��X�4q�Dj�R��6�*%2�$H-�/��*�F�����+d�_�fS���dy`%����O�wY�X�ų��9N]�UYI'.�zeE�����ӱWڅ���p6�G ��L@���w�]Y��o�r�(\?f�.t�eq�2�]'K��[������s��%�_~�Q��<�R��nU+�74!�em��Cp�ⅰw���j)}��/ňy���TI�>	��]y��?�(�E�$�pK��ؑ\n�I����[bEyW4��,�z{
'b�Z�╔��z�;5�JԙMN��6�J �ejV>o��&���#]@q���r��6�I���_J��H�{���b���PӍ��W��*�Ӯ	1�4mVz�e��ë�o� i2m��,ߡY���x s�kD���]︪�`���W���*�^�-��0�F�N�CV���_E�!~�m�U.�3��^exU�nA䟸a�C��Qt$em�}�c�V���N�SG�Keeb�K��n��ʩd��핗y�,�O+G:^�G��$Q��s����Nǉ�U�)���(��#1���*��H s5!�=}�{C� Z�Z�R�<d6� m�J h�A���՗�T���:nؿ!L�w��>�-2����d�.î'+���A;M�o�C�'��*�|��m:����a��S��,���IC�����xNR̔]R�n��aE�� +��|�!!u\�wv���2���b����Yv:��/���u/�#v���;S�T���̇�<[�?/[Z�v��@	�����k.�m
�N[j>�d!F�P���`�aܠ���W1^�H�>&�{5�1C�p);E������g Y�\&�r~F���x�}�Kc]ڢ~J�N�X<���Qs��g{�/����TGg����}ӡ7~؟�a����F���M���DK�:W}�v��kpM[�w[�Y��B�&�7����V��)#{�\�����%Lg�$��d����	)gZ��+O.���N�� �訽��\>5�Z>��RG�RYpN�@����mv���k��Hbc��Δ$����(��7�X�P$�����fzs��U���z��CW�ݵ�f�Q��~ܦLE�TV������oUcl'ΧnWk:��$�eq�����5���ɴ��T��:�䊺�s���3ފk&�F"~�{�{����V��>|���1j)��7fP\=���Y]!������y>����~���I����b��=:�s���9�2���A:�ؓ��W�l��wܭ�]�S�i��}��.՞��Q�+������3j�&��Q�N�_E�̟)ڄ��ǫ�{����m�.ͭ���D�]���DE0��"�N�I���L�Y�<b��!��¯�S��y0���'��L��ލ���^�Ma}���5'�j��M�����kw��~����I�M���qg?a���Q��4��|'Lzwn�`�{��|��<;ۀ؉y��C���(��w����YxL�Z|Ǫ������òjֆ�"�ۯ�ϖ;��P��C<s�����uu&ԕ|�6�πƲ��q��P�����y��P��w�e7���`5Jes^�;���m2�T��j;;������b^����I�^�ގ������H,��/z��,3��I�%$?�+K(�~���{3=	@P��ю�� �w[�_��o �s�u>��DM���U��<3j�!t�g���d��29���YG޾�/�=����ek�6h/!����RpNN%��������5N�]m#H1��:�sD!&N��.��pc�?��^R��äH�S�!u��ABϦF芠w�����ɝ�L�o9�}e��9��iP~�x����7��wx�9�9@4��]��5�\Oh�'A*P"����h�c��)q�aH�y钲�Wl����})�[=��zMq��VJ*m�Ϲ�]t|PZUf���.�?ҥ�wb?�&����e���9/~~�faHLAge?�S�
hKZ����^9�":�)e��D@�vr�d�g��Q<L���p�>%����ø��v."��=��A�",̍0��uM¡i�UC�cɔ�~�ܤ������a�֏���W'�൷(c	�G7H2�B����S��Ki&l�}iwD=;栟Q��1���`8]5u�ޤYd1(\�T?�F�ȓRЈv�r�tS����O���1�X�1[y�5������}����5)���+;���Zk1n��)tN"�l�v����m�̧aʵ�[9r������;�ߞqr-��R6{G+Zq��ɢ�$�����\<֟��P��PK��:�kC���&}O�E ��=�[yQc�h��ǆ�]������C�n�O0��qR�����8们�3��Q��j�d�M�Rd𾦲���%>�0��E���]��y�<X�oc���n� >�9𥘱>Q��%���f�����`�O���������b	UJb��jd�VI�4)@�?���0xMo�ۙ%�~��x�
�0�ݲ��-_�\�<������y��J-��AQ5V6�Fs��-�d�U�e! ��x_��U�+"!y�t����$:J����K*���O�u�f�edul�%���o�z���C~C�L�~E"S�����cz�����	�E�/���	z�9_��c,rm-�	��lԘd�	|I��2�IĭǹNb�/.-)�H�ke�����!��b2���`��0{���`y�
�����NDx��s�-��XVƧϷ\8N��p���cNX����L�}sE�I���WlN�8�z�\`�����?��
G���G�ޝ'g�^����.g����|d�z8����}�V���<Y|�����<c���X��bo�$���hT�\���2��M��	y�^��V���O�w���Y",n��ts�U�A�n���m���dF�
��ۥ�.��	�mz��2��/��m,R��_<�m��K��9T�I�ٜ:�������S�-qR��������L�����3(0����P����;mN���U��G��j�o�bz�	�P_I���/�<�}���� X�E�o���楕ɝ�l�23��,f�~�'��<^����:r��G�]�u�2�k�6 �?̬WOl��K1�ђan�[c!�0,�� �J��	�c���T�B_l�]b:PZ��Aa�,;(���7��6��I�7��;<2��`:�:��#�$*����柝�0���ݮ���1��2��B���}&�m������GX�@' �V���gYMر�Vg������=mTe-�8Y�@$��w�w� ���W��I�\[]�=n[��y5)�K����5TrӘLXmWCU(�z���{~���b����?��n{F��b�/u�K��M?�T�7��ݓ3��<#TP]Qj� C����	��m�vCj\�©�F��{&���I�Fq�|��N���Ft�+�̙F����*+̦�i�Dt ��βNg	��u�N`V�_,>S��Q�:ߨ��)�SN���j�Kkf����%���زm���,��|�α\�@���`'���DJESr/��㬸�"e�|�'�����],�[*V!����ͦ�9���Kg��Su�3��F�3�!�-A�bG������O �4�o��� pPw��
�<J� ~|�ۑ�¦$���^���c��FX���T�Dd�U�����)M�"z��C�-��J��:&�0�F�������z�����<���Z��(>W�f�����$
6g2�y��4D���W�q߸�'�Z?t%Օ�"��� �s���2#(��&~B��ͻ�t�Xz�6�8u�����7G��OT���!�.�O��;��G��_0h��-�5��=�n��<�ӦB^��R�Xq�X#�C������@��@;�w5p�K��\p:���ixzy%K��~���=k�6�%�6�ib�~��T�����X��˗�ﾸ�򞎺`��~!Л���Et0n$��AL�G6��IƊ!f�G��?w#��Y>M�?�cӝ?\���ʩ+�M�,@���Y��J�{�m��1�C"e�r\��Og(��96�к�Jo�lŤD�9�H� ׆)7V��w]s�Rr#��n۩꟯�'��8��H�]�Z;
-���ҏ��a�r������������;����GYb�&gG$O��G#�g���$ ��ba����n��cO�/�k�<�mX�	yq�=��T��ә�}��������c�F2�K����bcm-�u�eA-���xD�p�|�-<}w�FU�a"@���4(�^��q*N[u�$�����J$F٥X��=����M�:8x>ZQE����Ǩ),lc�?u�����H拰�N*�a�t�s�t�c]/�2�t�}���88!�����O�	�c��TNn?E�<�`h�4�Yv��m^���h^�iL���a�XlH*���Ӿ�_�������蒝���u��+�j���Ot��O�C�Uc����`mG��w���'N���}�Α�|�R�t�N�Tj7"�7�m�+o5H^`�~H#,B��-���>��7��-1����6=��}Qg�J���]#�s��;�ִ��L�H���SQ'G�V�U� ��>�6����p�l	����X<�B8��7�H�8��h���
4�f�3�m���j��fڔY�c���6�V�e�'ǯ@N��W�7L�cA�O� S���`�)>�)��u��$��Q���C��|7�#�Ϭ�E d������nX�h���q��v���B�3��E�O��u�ylݧ�������S|��e,TZ�zPN,��lw{n˷��Pf&rf���nS��\+��--`���O �=ʎ��6r�0��B^���bb$��7|z���-�3�5��"��H���[ۗ���l���KQ�b��g���<{��y�Q��w^aUA^�׀���u@=e.s��>�o�q|Jr'��re�����B	�^#v��q����Db�K;�J�G�CLI_Xh����b1  hFw���%�dBb�\+��o���f�jQbn>�ޛ�����t@
�����.�g�;{N+�B�݄�lh$�?\��Q��VuAq���N�x[d>�ز�v�%up��������ˤ�.ͅ���ls]�4�mƛ?/��k%�E��T��f��yK� �?������0n\�n��r��!��(���yR����7�Ĉg~���a2����s�5먑�j�̧$-�?�]i��/���eQ�30�.����f�����麼�d�g"�ϲ����M�~{Wb
=t>P|��5� �̎7�ۯ�n0�m��;�+�[& �y`?�:ۻ@S�J��M@�gx{,�9چ�u��k�om��	�)��C ��e��Ϩ�,��҇���#.3��@,U��|@oNf[�TR��f��P>���~.��< lΞQ|�놋�M�,TvJ�Q���H���`�V����mg��"|i�ǃ�4��� }���x�`�gKZ3���f}��?�,s�㵋~��G��u�{d�no�&�wL.q��Rxp��@�%����t����t��2��ϓ#'��4�M.xŴ:�Z�]������]5��x�*���'do���v=��
��q�q�5(��m\/'�&;LB�HM��T`���󜏇w !<J�%���_�/�m���e�l�m�W��6_�x1I	��[�ls��F�e��*��0���?�8��wM� ��5CO~�4�_����P���:�J�����5�0�h-n��W&�>v#CȒFRT���FJV��:Τ 3Z�}�~�7�3�ܡcu���	G��&F��<7��jþ�d��	���!@�:�)İ�r�_��~�ָ��_�r�uw �F�u#ٜ,�(n��|�7I�xv�ʼoe�7���/��w�7{?�� se�9��0Sg6���`�pA�(������G��r���`�M."�g~�w��?�j�H���4�ۼm�J���L2F�"U!��]I�Q��5qj>/�$��9b�!���t|��,����@�Kj*H�4�j�\(����ܖ,q̠:?iN��V����e5��xh�������ve�N��S��߯6��f"�=(S���ӓL��z���3��<<Z��{�s�O5�7k����Y��J��[K�� �oJFL~涹rZ)�a�BL�ۖ/ct��)p֓p+gh�Iw`��+t�<�j�q��A��^���+�|J�;ĹO��M���%�VS��\;W0#:M���}�BF�Á0�
c����;6Co4M�� m/��F�#����:��<�5��KXl8�fb�Tj�4q��m�!�f8M���G��mJ��c|�'_H`�_�/'�OtAΦ6���}燥�����_}{����N.��.h>*�kI§eup���<��+�,�b�.�&~�z���o�>[%nu0���q&ƺ�GQ\^�l���k��N꿋`����,8�cOL>5���������������=��~R�.�Sѕ!��Q�Z��w�r�͟�T��K A%Di�v�ȸ����P�4O�e�)�Um�������A7e7���Z��Q�x���w�4������ן�L�cS��67��/�
o&��=�P��X�'*}���Ϩ���n�ʔЇ�	�v[�q����
cw�{1V"�Z'����=��U+��v*s�Eu,��`u��D��>��-����-<OQA�R���>�w���n$:�k[[��D����{�|
����ǅ^���`~��u�GU���(=�M�d�"����J�o�(e�v��y�6�G
�N�Iz��;�v=��~j��������et)1�,eI�<B�*ԁx`�3
F��PQ��#p�"b��_��Q��Bל���|i_�'d�E����:%��'|2�f�{�u��ӎ�t�1��J����s�5�����l��"�)C�K�5��'˪���M�s��to�D,���s��r?�!&���M��ڕ�_�>5�=�G�.���	�\��'�%L��o�`R���F�q��r�%�QI��7Jk�D���&�w���B���I��i�Jt�>P �mA���f]��^W���o=S��Sǧ3S������J�e��}�ނ�_���; (�M`M���?��?�,:p#j�Ika��Uu�{�� �`�G�xa��b���E*fJ� ��1>kZL�i8��Dr�5�2���;�6��&q'&��u���[�Y�;}�I~�GT�By=%1�����q���wO
]v�e����t8��x�H�^��F/�=9�&��~.|��͆�4�x����Q��4�p*y���(5�6S+Rx9�Yg��*fKp�m�=�����`�jquK�1P����şg����sE�)@'�h,���I_h��p��{3��	��{�"��n���6d�&r�k٭v=��X>D=V^b`��?�ƿ����(�"�ֺO���~��� �,�N2?O+�˓J�bL5$�r�|�}�#����=X_~S��̜ Mb�P�q]���]s�]�u7��������.�S����UP'
;�h"�M&{��}��Q�R�Ƀ�:l�� 
{^gC\-�n�}�F��Ӂ'3S�A�v�D�k���Ɨ�Nf�O�z=�1S-�X]��g���ӝB�`m6�6�C��S�}��E����NĵNoԢ.�z}M[�0�v�ݤ6�`sp�T�I��o#�yWB�&>rw���V51�2?t#���,�Q�Y'[C�x\Bn��+=֢�H �����~�}CD�ݛB�h�'��Q�1������_��v��Ф�������s37� ,r�^H�r)m����������Ӛ?������>�K���s�nr�޷䣈W�xő��v;���	�h)8�rX��Z��?9��y��U�OX��b��0�F�lF&��	n��X�	W��jt�t�`$#�G߆�	�]����=/�h��ʲ��]��fI[>@Pz?�:!�bF��ڍT\c����
7bm�$2��;��|�/������ș8a�U��U��*)�/���G�B�,uQ�s�H���5T>�5U d��!��Fv��/�0-�"P�{����$� ��6��]B&�u'+��)�����q�X|�Zxo�Ԋj
D��m��L(�`�.V@����5g�_���^�D؟��m���%��g3֛D�H#dWx~h��6ݼf�.\��v�W�c�-��,~�EU�>�WWC��0N0Co�sx��l���f�l}rI\b�0�l�,�&�AW�'�/`՛� {�*o�i 9��8j�����_�a��lJ+U���K&:���VA���<�S�lҴgB��Ƨ���l���K��k���N~y��D��5 W����6I}�@i�y�x�xŠ_ �L��x�^�U��˨?��HB�+zs{��̓�@�����~Y���c.2��Y���UllY��s���զS�<��=��xt�"c3����i��^Ƌ�l.�'�@T�p�������-|gެ1ߵ�"'��)n��V9�k�E�@d~��Z%4�=��_��2[��?"?1���Xy�1#����~j);�nV�6���ߎ&�H� ��r$��X?�����'�qҚ���v1����e��Ԙ�_��N�Ժ²�����[�@��~��~�s����%/���0\4m���C��khb�*x5�pR��	�י;�]wp_4h���(��VZ�-��������3G���-�'�`�*�(/W�:�J7�2�\�������[�<ֽ0w^�E�`j����랬��t��G��������d��p�yy�aS1h�_b|�ox��;t5�PE�n>��Sx{p�j ������V����f�5���ss���'��i��`��py�B��41�	oX;%�A������֥��I3�I��pv����,w;y{���0L��ؕS����'�w��zWCan�z�B����+�n���Ƒ����6K��=�o�u�Ko�=��k}�����1xq�R?+�E�<��6;���M�������}A���EGe����Ȳ����#������w��m� !A���&���0����z������R���b'�ͺr,m�8-s�������b��&��6��m��#��iA՛!>�D��mL�9�3��h"�Z��.E����n�����Ƀ�����e��^m̀h�0C����yB�G������h��q�v��q��ĩa6ԥ"u	�8-�A�rv��x�X�+ewE��W�����^�������<|'k�����%u��λ&i寂T�
{���Z���ƭӉ�23�\���jK����P����"�c�dR/=�ߜ�6T�6����$�%���ɔ���*���Aa��pY�!�!��)�K�ϟo=-bwf|�t��n�᭦�α���<��k�ʱ�c�x,��-��1'�����Ԍٴhu��G|�����ՙ>�>�A���h��FG�[���IsC���7��S�飭�ed�e��=!:?��躛�)����C�w�5u�m�Z�V�R"�
��"#�
����
**� �VA@��T�2e�A�=��V�����|���}��O��Gr�{\�u_�sN�3N_�M�'�[����Gܶ�ͤ��b �M�����Q���Ƀ�C��ov!��g�yt}�Q�sxo�oQ��;�˰���G�������8��uKFS;S[}����(ë�fPh���D��/��e��g^5�5.J3K�~�AP��P3�1��Q���gY2UVkZ�5N�G=8�>��]TXK|<��g}
�B}z$��R��{T)
|��7��\��o��k��-�c�7���P
j���[��vd.����~��֤��?����H1����2���8���]�kc&dwg����O8�?�:�(��/����T���v����7�����?Ӕn�nu�3<z7�SK�O'ӗ�"��&3���l�/�j���ƺO�k�@���'(��\U�
4W#	T���Mx�g�|zj��4uR�im���=�/�O�Ĩ+�}WMb,=n������*f&y=ƒ�]�."��o�ٽ��"�"٣����e�ј>�UU��'��o�k>0[�,8>�Rx�z�z�� �3v9�>:yu��|�.�]0yw��Mn�\�����X�7@}Oؖ��ʢ�?l��ڷ���e~���+4
�|ha>�Ac}�f�"��A����+`�_�:l�H'�'*�?K�GW����ڨq�"T��ff�F�*�.$.���a���?+nL5�p�OɌ��U�"�V!q�_O�����g����?��
v�����a��p���� 7��V�s�
�{������XI<�_�Q��-�)0���*Q��W�{��7�N�H��QP����(\�N.p�2���9����i�WiX@�6n�U��t:�BN�N��}�a��ċ�z��=�6�`��Z����|���&���k��`��ƞ��N�<N	��1�د�~��B9lDN�q�W��%�嬠A�e��qD�~��ÖW����[���F�\
���k���D���5������11�Ig������|�4J=�!*� h�IU�c���Q��4�B�`9���,��*�"�=�C�5,=c~[#���r�Av�r�t��-CPJ�n�!cqjG���o6�dV�D%���'���e���G�9����ŵ�	d>��~�0�u��k�M�Ŧ]]Z1��t@�$�8��Q}/�\'��ɵ�� ���aa�S��#�I�kl`���A�&���E��bY��
x�#�Dgǩ	�98+X�6=l>p�8�`�{�뾕3���m��R���AD�}˙��4)DP<Iy��S�W9n�����J�o0��4u�M�PC��|r��3l��br9�{I�	��·�~�Č����O�����HO�	TC�>y�o 2�X�����(|��W*/��T���/�����k2����J�T�=���m=[Hf�NйVX����a�9���	��"�]Y��o��{��UJ0%6C'�������>>z�S͇?x�fg�z����}�"�g~է�οd�;��>��( ���3��R�PC���~p�t����T�,9�^�}��B�x�Rp���.k-֐����:�m�;� �l?�600PI��d����_c���Ke�c뱜�����z�<@��[�d�`J�1Pʞ�cpG��8!A�+9��J�n-�a��g
��9g�jT<��U�_r Z���e�����+ފ�?�S�ey����X�|T}2g⦱Z���ӗ+�(tk�,�hc"��y��>��G�{Sxs��(�]4yc�;�>C��w�=P���p�93$RX_E�:r���+v����J!��wx_��آF���;X��D�/�����o�%U�4�,�v�����v��eņ7�x�QL�	��~\ �AP&��&gv�e��1��ێ�n*6�ԯ��������a��[��{w�<t�<ZnL}��|=y��Y�	~$��\�����+t"� 3X�;M�m��t;��7jS)y�v�k�S9q{-% �����g�}d�,���[��6��:P>]/�}X�P#f�V�4�ZL+X��w���� .�&�%�C�����W=UIp~�	�+k��N�I"ӆ��/˙ga)_YL���i�������s��u9A�Q�sG�7�s�at�{�&G&&�10������{��,@�����?�~��Fd�b��ẀPT�P3����{���շ�Ru�|��gzh2�,1rY5q"��M�t����Q&~�ʯ&��B���~���g�>�̇O��e}V�2'�YW�A�{���{�`ZI�F��ӂϢ��U����ؑ
�*�Ƣ�n^���~wh*��9��_��}���������o��ć�jnmF��:�D|��We
�D�P��w��:��*"�U��2��%���U�nc�MK�ح��^�q��I���uG� �^�hX+�a�������]E��$��<�6�R�ɫGz���3|���K������֯��`=]��mD���i�b%�ͩJe���rM��Q=ޅ�;Fc	M��kgO������QK��d�J�X/��x�P�D������T,/�*���%H�ϰS1?�wpC���c$��.Z5��F��k��7^0z�@��i��� �m�ZOH�s���<�do'H�8�{h
�+L���l"���UD��mp��w~�dT>O���}��΀�t%���附���Z{���Le����w�t��e��@3?S��U+KtG��jHY-���ihHb�c�Y�#�ذ#,�/i�v��و4�\ .�z�uE�
��q���T��v��i���}�q>���5Ųg�� ��Un쫎]��l$(ץ����:(�2q�.�?�D��	{7U�Yļjji^ș�i���é��s�)M����M�f�O��}`��܀r���~�p���#ܩS�_B�'�B.�:���:h���rz�P�3r}��Y��2��)��vJ��ЇVǹ�ꅺr/�Q��ca�o�ԙ�M4���ҝ���y�wʧ�f��֖�R���S�^�%<�
�"��v���}�T���q#�5���(�Gk��RB�ڪ���k�>�O�� ���f�	u������t����ky|@A�U>�IWe�5�b��JJ,�j]9�$�w�#�6��2J�Ŏ80�#ԋH��"���%�B�P���6���U�J9(d�˱�V����6�}�.7�MJw<�3c�I�9rKպ|FWz��wh�Ц���+�Ğ�i��
�toF��*�W�ڴ�@@�F&��aT-V�h�!(%��X9�lp���I��l��"�f��~3Z�UM��%4�(���:��N>=�h��{QA�Z�K�8���0�x�A[��d�(��K�>�Ğ�)�˛�t]�,԰��@�˝��~ܒ0�p��%gil�]C�Q1p�Ɇ�F�k��H"�g�%�!"��N���+�U����D߉U�^�yAk�}΁�z�dj���F~�O���\���!^u�'��0���^Ԓ�r�� g�8�9^UEq�D�r������
����K���<A��CWA4��ze 0Y��zw�fZ�
����[��c}�&�[JR�Ry#s���s��w����4��4�S��H�t�U����	87ŗ����c�'<�Yj?���o�;Eo�O@�P��z�Y����,q� nY�ǘ��ۯ�l���kM�(P߰�����d� ���u�K�]d��Ʉg`���I�2��u�m��O���r�py�t�#��ˇT�=T���~���Ь��?'�bϧ]��:�� W�)V���f�5�����cxfbe���)��Q���˩�Y�8&�a|��o\��2f4
|�,�	uǘg%f+M�[Z9#i �Qvy2��䦕b��:A�`?����ѝLW��(�K����`�>�����uos�,}�܊zHM�� rE��ruHN�2ٔ�n�y<��l"_��xd�S�����W��=�͎�@YC�ƨ>�wl(��<��Z����Z,���qA�����Pp[E�h9�[Y  �O�����fq���{$�����r��|G�U�R��z���p���a̕A�+u<yF�|�e�imoF��9�0W��]9v�'=�Szp�~�JG��e�X[���;��HFi0��C 5��.�$�	����a�<�?�~ �J�W�8t���SU�������H�W�<kӌH>V�� F��U�X'����qb��]��w#�z@��f5�����%���{��O��d�ꛆyL��ZD�u|����,'I��0�l�q,F�2Û�u ��&���kyR�ֲ�ˡ�2@j6s�r`��ﻻ�z���,a�4u�<�E��E����]��:R2:M���]]JN\��I�h���^�'�a}����ac*z���oMmq.�H73�j����dv�)l����?,p��k�o%;,͊��Sb����p�U�G��r��&~�Jl����G?�D���W0hvs��p�&�E#��rh.�%�g;�`�'^=�;�U1�����Ϩ�-Pz�7=� >�d��A��c|ZB��I�e`����uD�/�����JƼȜ�VO�U[`���	7B��Oϸ�^Y�*I��}w�޿����޴����&��>*�ޖ��;oI��+�UW{-L��`��D~~+�R�~D_է�	�'��E7���[�*�j�˧5=��R�q8��Sl�zOĄ�wk����5"c���y��-�#o���C>�|��|[�����[F��䅓��I��r�jߏ4�Ӿr=KB�8P���S�I�h"�4�����V�MU��c�;��3�/q�9��_ }|#�%���䷩�8���^���G�b$ac���rN��RZ��L`M����dUTx���֐��R���JQ�D&c/gtٷn/N<g�D�e�҈��{�Ti�wM�! ��GU��9V�ڪDU>#%#
��9�$�暛�D�XZ�����^P}PCWHw�n��Q��|����l�Vp�)���P���{d�!�'��y<R7Υ�E"m��]-����t�o>�]gt3_ڛX,�@
��������[�ڨ��(��(à6a ٝ߯���]e5[�"w�#&���OX�5Erͽ�C N�Y�g���]H�������Kɟ��+W� o{�hY��Qb]�a���/c�~����,s<4�1!�9){8	��YoE>r�n���T�����zeJB�p��#&ng뢈�v�q��]�����z�-��Sg��iBl�"�Q@)���gU��f$���}w_��Ŧ��(b��g�H�X�%���V���@�7��Jq�N������%A����u�2�F��+�+|`?���~ĿN�4��5 hb���(���^���h�Eߡ�\3�LS�3�|�?o�!z���h�H��.?���7AuwX�#NV�Y�,���|�0��	˪��Ikau��������#A��O�d�y�+,]S^]a�%y�&�)R2�z�r�(�#����Z� ���kA#��m��BC%�2�V��P/�X�t�l��O�G��sE�Xye���ҁ��Ȏ���$�i��Ώr=i�{'��v�Q#
7Y��:w�cѧ���8�=b��\^�-(um�std7uA1��d��t�MVD_�N+�Nq���k���XϖL�q�S�8�>�,:�cߥI��N��Q�
������+C}gT�|i1���|5@��D����:��#�w﹙z�!�*�*��`�H��x[��o]�|���l�
�+�!n�� �{B�|I��Q��@$S[h�fh[�ai�>���B���:���u[a�)���rh��L�6ϭ��9���i�u�7�+�G6j��B�
�+`���-2��W�����z���؁B���lp%R���>,L>�U��琹�윌��(hu�4��툶�ӕ>2bҁɯ��.�68f���>����gͯ�[۶�A	�]�ĐGk����\�p#u��Q�D? y�_g��ܖ?�����(@R�i�k�l
5��
�
c+����|Ŀw�P}jv#�U�7���m���/w7�q&W���M q g�Ip� �OcC��go��V���	cum-��$��K������8{.�F�����L�hϺmk�8X����چ�+Jq��|�O��D a��6Y=ۆd�?���	�.����
�����}��u�C�3�N�	����C�
y9p��þŎ$ܯ2��=��J�fK�di^����ƹ�c��� 	X��W�o,�X��ڝBF�N��K�x�|�X�<&��>!�_��+�b?�.~WZ��N\���6�ͬZ���`$�ѹ�X��4�(�X;�����B�`&��N;��^�acԡ.�Z&��������Z��T��dO��2�Iu��<��h�S۲ᡸC�-���g8q�M8��w���΃�0���+%�c�����e �V��vm�[9�����i������Q�����V�I��� �w�9�s���˃D�����������]�c����?���e�����c����dtO��:o#��	�z�������JQ8�'IGe꿙$v*.a�x����Z����D��:L�-+ϸ��ʹ�l�LPp)w�	{)ly'�/��C��"e���797�/�N�W(߰:��u@P��h^��@��]g�7�Đ�9ŭyQ|�f���sKM4M��w��t�n는��݌Y�-o��F�r��p��N�f���^����������7�8�J�IkcۂD��������"��}���-R���FCC(�$0���\�_6�*~'zs��n �/q��̣���?T~��E�UD�"�>Jt�?����L�4�nuT?~ ��Ð^���u_�Y�,��2:�uѦ6�+4 L�,�h��y���IM�Ҫ�w����]%���c�8�,�ןl�O~1r��e��L�方��{t���w�Ƿ��d7����X����8u�m[/Aҧ����1*g}���X��M��䳖�uq��H�}7j�/����Y͗�UE/h8|�0��&��l���eh%�����DϾ('3���������Y�u��1ߞ�h,e�����G�HN���#�gá�h'��� ]������h�Z8�Z2�飄�	����[�<jd�>���>����t
>�v_��U��:7�G��Q�o���c�����]N�R_�˼�r�:�Rfc�qaywM�կ��T��Jz�˖I���(�l��� ���%8�n]h�lli��5����A��;�?+�������O��m���VϬ<�N>�ݼn�{��-m��̞��o+��R����VA���WxP���f��cS
qu����8��U�,��^�4�f�x� �-N���������\��[�@��L��i�M���V�B\�no�"c}!k���5^H�ɪ� �F��-8K���>J�W����y��M�����Erݷ	H�|���Co�}�rK[�����(*��#�dAh���s-+�&�F4�X�y��NB5Px
�Dq�'"��?�Gb��L�#����8����΂�J��q�E��� Avj議7xȁ�i�C���a��l���n���g<������#�� �7�%*�0ͽ�[CnKo�+Ă�8�&i��>��M�)�,��m{�-�,��2�$�	&g.�i�0������2&�o6ik(�L���E��d�u����ε�ӑ
��[�<x����s��k��G��cK-X�W��[m�=�2����9P\-�V�� ��Zk��Ҷ�ǯQ��zﰱ���s�q}̡�A�l�JɻV:��0^��X�ndO��6�c�n�1|���e�t$*8��r3!��߲���E{F�l�k#��P{z�:~cN�晙��y4SQ�[I�1�Y�R�m7mo��u�u�RvI�n�U������G7XO��S�B {6�4�L@���nM��m�|���4%Ӗ��h&�4��m��3�.���de���VV{��	�(8���xV.p�")�(�h��e<wX�i���~Y�#8��N�y=86�E����n|�a����������L9��f�I�O_9�
dr��#u��Ļh�����e]r�Gh���2H�G�F���+��!�T��%c�q��ضy�R>�|tۤڗ�v� qX}�4����t����έq��m72S�0WVz�&S��E���2Qܒm�TZ�%l��I���˔�۹}��&e�����d�̒���B��*3�]@��=M!�mK��Ih��qsq#��^�6�h��� R���Q?��i._i��f�}Et@����A ����78C��;�V�b�'��a����`]�*l�9�6�^���k~vP��X��Y�r!N3|��4hMc�̰"M}E�Aػ;b�.���<܉$���x���7�7J�s��n�r�����U8�Z�捣5P��2�V�p�k��N|��N}�J����L��Z�X���6�B������C}���䙊��k�\m~�%O�ȅrO�DʉԆ�;nq������ۍ}�e�m���xb�Ci��`6^��rJ��9y�������,�4��*��ݦ+�հ>���h����/�r�7'a���[	�@�_� {����V1�ݦ�H��/�6���4��o����Fz��j�K[��&���]�#oa�u�����_L�)ڋ�ℨ�������և
n���8���>���!��;�!�嗪Dwo��A����ӷ��b�n����FC2"��t�9���a�0�׼58gZ眈~~�Eҙ3��Zä�I������qI�:,x��>����f�J��>�<7ѓ�Z| 0`$k0؄�˥ �'W���"��+���\S˅g�Fr�-5$��%��#������6f��A���?{�[��e;�Q��0��Z1+�Q�ޭ5x��[�(.z�I'�I#*���*$%ɉ�v�\[}��l��y,$��8�?4v�O&ƽ�p�d�Q�P\�m!#&�T#���	y5�T��.S�Q�0��� 6�E��V�2�?����d~�~��Ȱ��jz����ǯ�XG;z�=z����/�|����qr�S�KTe�8y�����r��l�|�	��:�������M&UU�֐_��3u�U�yY���x�I}ai���h��r���9C٫g(D�m���^��(�u g��y�G#�`�a�S���1^��ȣ�o����8�/��B����2��}^��ϰ��eq�<�����w{���ԴG���=#27�:�57i�v�[/��U��r���з3�׶��Z^��8�[i�U˝��_O�Z��EZ�̭�1Z�Ü:����ۼ����Z
�{��&Q݇����:0f`��X�g�6=W|kr��Dq�Q�^H��\��_��Q��m[U�'���	�O,�Or7�c�����,���/�(:9��ӗ����e�X9�.Y������V
�ܠ�{�wN?\m�Z�w�yp��='9��\��Δ"�_�H^���J�o���fn�61�|].�R���'���n���*KH�¼��jjk�=8��=����S!�k��-[
o35�����}�͠D��ʉ2:ͳ��N�S�N�1����U!x�ݪB��Ҧtc��`��ŧo��A��R^7eۜF>)�u����cKo�zQ�2��P��P� ^N������}�_v���c�[�,�����y�W֚�|iWr�ջ��3޽"'3��KQnS+V����z��J���\�AF��L�٭�l�@.l����ܶ�H/�z�k�loT�X}(D(��#o���Z�~!.��]}���zG�M���|k(������{�����Q��6fd+��3�$Q�����݃$�d��dKЂ"�A��C���c��BE=#[\)12�e.�g����֝;u7Ζo4�`Q�W@)�}���,��u�'q�#��a��[M�3�zȡ(+�6���%�V��Vx;��x��dϠ���o��P���a�.l���?��ۗ.ig	�}g�8kx~&���t�%��֫��lg?�:���jK �^߾�5���r�������b�
�Q@7�N�R��=�
Q,���;��������<�l��ߊ���W��P�,��C����ɓ���&��i�C5^�m��l;�j�C;	fj���@o�'|����2��Zmn��C�H �W���o�$O�sF|��������-1֨�o_�X<f4S�ߡb��ײ�!A���9��S��rԘ��zD$��]��i,��z�4���f����C��Ed/�k�>�-�B2�P�}�Fr��Rm9�x�J��1yW���o�C�J��MѣqK��u�cjPs9'��!\,��_]L�kÃ5��iǾ�@A��&�^kI#r�r���9I��S� �]
���P�j�Y���rtG�.����h�y��Iy����㓇IB�Z;T���S?���BQ�h��h6� ����5qn}�6O����"�;��T٣΀�ɸ/����@���^К�4��yﺏ��ٓ����mL��<����9%�
;;,v����G�!}۽-�L颅��W�/ |�Q�N-�Y���dה��t#��KX�'V.)�c�{�Wdz���%KyJ[���Akcj�J������i������)2�H6��]>��m��${���(��H+̠���Fc�r/s�xIX��L�����ְ�b��D��^�JAf��&�
��������*�O	ޚۿ�+h�4G�Z������i:�6u7��/���M70R2����(p�����B^(�S�q�k��`���Xu q�h��M�/KZ��Q�WG��2��&s�'+�k�ڄ�w�2o���@�/C�����m#�֌��&F�Xi��[���`��fa�um���܅���08:��.?�Z��6L��W@!�j�@����Nd���#�iHh������]��'��@��M�������D1C'k;,�m7����'@<>	&�d}�=^(�U´��"���p�
��:��	�tW[x�z3Y���ff ��PZ⡤��D�B�w��� I��"�j�0�����dݹ:{��:j���������I��_�Mӛy�R|��3t`��X�91<⇳' ����g]00<�Nl�d'��mp���r��?��%乙<�Tzf�๭�V�J9�={>������ ��y'O�j9W�[Şw�������\%A/>u��?�vǻqE�v�Pd��HBWu����YB1t&���]�f/OWcy�ipO�|+��ig��\��"c(-�h/8D�#qʖk1��R���P�HI���u�%�%��!��
��{���)����4��z
<W���f�ڻ��օ�*ۉ��W���7�ꚬ�
��<��'u��k"6w��5��nqg3x������$��*�~�%ry�v2יWq`���څ#�8��7%�U���N�J��3�Y��uy�7kA�#\�R���'꺏���u'+�ߨU6�p�^s�V�E9�L�?�L�"��:x(z���g_�N�<ߛ���'ɿg^�� ��;�'s�n$�W�˽Q��@�$��t�'/�C#��+�k h�=��FsS�k�sAjjf����r]�Кᇠ@�˓Vw�f���z؝i}`��p���ډ8L�NQ-i���,7 \�D�[2Y;tA!�/�4>SV��=h�}®�e��׀�O�-��������w�p ������V��O�[j�L�˄�+����od��F����*�
"o1w��b0�tㅶ���w�/�'�qY~S1q;�u��\ʬ���9��}��+
W���U�/����J�L2�^]�?P����V�Q;��-z��ܲ{�ѹ:���2X�i�
t6���1B�����K���9�}b����%Wj6xw|��m������,�|9Kg�Q�I���4�Q�]�y{ΐ39{�CM�����2�fCґ�d�;dgP�|�B�H�!-<������g���45i�l��H�nri������׀g1U0i��&��N�;��6�&C)�]�ֵ'K��n�Љ�)�S��T�c"&>��|�@�qe�,Aj�kC��/_fk���6oT�9����M�A����RT�_�?xvLxӸ_���hs��ݻE�������T+�Z'߾v�|����Wu�2N�ޓ�5+�a��zծ�lb��G|L �;�xEvǳ�n�`�0l�ibD�o�{)w�`��c~���kd���t����5�y���D��)�g�����[�|�j��`_��D��MK{���eV�H#Y�s��.�}`���.�b%F-����h��� ��Y��('�p	��T�i��� ���@%�>��~٦�����y܊�r�r�N]t���0Hcqv���߈ͦ�E�^,��SR�xW�Q��o�xn��9�c�tA��lQ
�2)��=B�1��B�|Z��f��\~{D�we_��b���XK�ڴD��ֿW>]���>1y��_��2Z�˚����4˷�'������QC�������I��"��ٻ�}�	�>jy�ڟv��ǽz�7��<@]\�O�KW?
��%+<QN�V柚�1:)l��7����ӶO�Y8��,ᩎA���	5'm��ƾ�ׯ�t>������ӭ��Ԋ)�2�����z�Pk>�^�ͨҞ��\Z���ȔOQ��۾kw��$" 0�)�|f$^*�7t.����z�A�Hd�����m4�X߯x�TL���!��I��|�^2��p�����%��vu)x$�|ɦz^���{�\��N��@�u�t�o�������*�"��'U��9t ��5�븷�)�@�@Al��	�mओ���}���*U�5����N�g�Cwl��ulZ
I�c�Dc�(;%�N������i����"��JX����L�@�<�@Z;us�[���E6C �2kq����$+�(�ߠӓ�gH�1���"Xk�MuN�p�&�y��äD?��.'�93�x��)�Z�WnL�M�=wO{}dtz ��d!�y��Fy�r�w�̬��9����E�V���`&&k�p$�c��=�eN�0c�\��s�v��"����/#.~l�ư�� m��B?�3�4k��ٵW���@�x;��8u��ۆA�9XA�W�n��C+�t���>��z��bw3Q��w�a��fQ����zd4|%�7�Cg-�iB_�n��Y�cd b�2�=7k��y����b���AjՈ����T��5�Ơ<��|C�!gNV��5qWï8�s������A�!R�cz3)�o�C�B�KX0owN�(��×��T��{�AK�Åsg����������VI��)#&�V��Z6�[�u�KB!N�i`E1Ndj�$��p��<8w7���Ѳ�^�c~�b�=�WB_]�'���KJ:��.h��ɘi�<���^0<k2��$	Q8u8�϶J��*��|�B����ň�fö��*�����	�/_>��ج*�兔�xa����������7)*�o4p-�|xȱm�����d����H"����@c�u���1��~�x�haXDd�(tZS�>X�?�Zƞ5V|�.:��Gւ�@N��`��p���E��8�ۓ��$�=�ȁ7�q���V��R��(�BK-���C��o~�6Ԝ5$빼����\�0�	9xt�}}�u�u��A%���L���	,�<*�_1�ѽ��hCW�>�<�@���B�T�=��S�-�9J|�MW���ct�OZ��m��������ʒ��>�l�k3/��t���M.�FJ��#�4��
=Q����-����:�Al���W�h�@,�l��aZ�����ƃIX��Sj"i\�NS��%O�rDߛ1�5	뼳 �ZC9�4<4z���r}�ū悎�B>��� �$�a�>E�˴�ٝ&�IPeiyR3au�C6���w�=m?'�8	0��|����͌�R(��RSjQ����vJ"ynz�Z��ۜ���CC~���-��%��C���-ȸ(�P��l�ffGDP��UMɔ���4
A�d�
W�4s���Ӎ���@�*.G�h� 4�T/@\�jX��vnz����C��U�S#��>þ��Q;�j��> �V�mW�aF������7��uG���3���B~�b{�Oh3ӣ?��r�DUD8=
j�倴)+�$Z��w��c�zC�8�aF�'��R���r=wNO:B���E����G�z� G|j��i�{Zˬv�rQ�N���nH	���w36��Os	���Qj6E���	*��i�sj�F�F��{Mߤt?V�#-����Vu~LEX!�]-����w/Fʾ�$�t�bR%��l����)�w0���	�[�e�F`S��C�Jtα,K�S��B6���fJ�����_�TF[_%XX�!���>:z�GlE"P-�	��c�ݥ�v������?�� ˢ�R{���MM�]2Q^�G5t�i !�j�f�d�1 ��5-�6��������֪��zX�Ȍt��#���v2�G�x��R�8�b>`����Tp�C��gdqs#���%�M�����ʆ�c[��F�MoK!�[(��
T���H�����o�&6�1�*}�8��b�pV�q��Mk�V X�_���U��:��F@�~~�cԛ�����8�m!B��x�N�%��I�ii�Ii�h����1��eF�~(�h����hϤ�W;5Ly�E�􈩻4$�9��M��hK=E�NSuAH����-]�α�~'�qx�U�A����t�{�!�)��R�6�x���V�ӌ��-NSZ�Q����ٟ5btN�o�pČi6�gb D{�����<��Ԗ����I�53�9�`��lAk� ���7���@�(GI�3����O@��C`Z<T�r2�,>��$�<`a��d�h����K�]1�*�C\�����*ņW{S\� LGv�Ak��.�2`Ā��~pO�$�,O�ʄ�A�GdXyعk�Pn�܀�#]�9���٢'5�'��6��	|B;$J�t�b˺��,T���#,ĞL�.�*w�P?j��DQ8�v�O���3ɋ��t�
5������x)i���~&�&G�N�0M�z�z=���Q ��:�"TC�9P)��������c�C�T�z��~�����T=\
��Wݲn�:J6��q'�mZh ���{Z��Gߡ���ꈯP��#�S��4�ۥV%�@ o��yO�qxZU`j0���h['eX��+=v-��zo���b�P5�͈��Ix�ă�R��'Fr��\��V>�	���ǎ��5�|ݒִ�"q8�43�0�G^g�$q�zq�|��}G��>����Ӎh�����4�J��P˂��K �>��n!.Ƒ����i�L̟��#�3䃮ټY��C"�D`��!NQ�)������Ѣ$5�HQr��ߟ�(}O��NZ`��]��|t����1Ϩ(��n�~�jA�0ҫ�2� �U��� }y�G�&�;�#6�8	(�[�ux�+)�T�>�$�+7U�d/P�N���>���a���V`DE����ݼ ���Bph���z~����3��U�1,�w��S���~�<S�~�O�#5�m���N
dm�����	4�獀n$�5u4�tt�Rz�5�S5�k|��&��ϖ$1R�O%e�<��D�G�vᗦ_<2_5w�#�g ��ϴR��̻�,R'��,�Z��d��J��H�����pqf$�7�(�&�X�^D�m:zCX�γ3�(Q��(�l�/i3�~��ZS1-E�V8P���r���$��BտOwo:l�D�`�R�ʡ|�Ł�T�1���ׅh9��E��e���]5�ħ#�r�O��{S�v)|�RWs��_����	/��Л~k�����u@���:�UCۈn[�Ղ��F��ʪ.4JGX̩ԥ�d�+��9�h�3�R�hA�vSN�eΎ`l�ڭC��N�tCO5��Ε"�=@ԤE���7?��H ���k���!p�x��Z	�%�7/�6e[
gīU}u���?�Y5���R�Ju����c|�*-�?�g�+�'��R����Y�ow/�-�~�Ԑ�7�X9��q˥E��XaU��0�J{n�3���t?��'oI�ݖf=���Ԫv�%(*��Wx^��z���ϓ�tnI����įCP�ҡUU����2��)Yaxd�_A��e�\��Q�	/>`���М}aKMհv�!i�e`��#(a�' ���+�U�I�)�a_L氚��Y/܍���?�z�`����x�0v��ǰim���ds�\[ �SL#*}ӱ9m'��x��ؤ���@u�OZ�n�����s�_ֺZ�땽=9���Bn�������+�FA�궝�٭�{��6ջ4�I�8�Rd�u
 �Aٽ�� �AF�5�Yt�>���z�R?b�y�\D��z�  ���ڧ?��H�K�H�٩�}~K�4�|B�O�}� u	�_yC�M��"(Nc��о����:FZ�����߹�A�Z�E��[�%J������C�Z1��!�� ʸ�Ȕ��'�#����.L�%���{a��nAǳZ�٧����4c�@�%�.6&+�} �Z����h���"����_H��%�x���2bRE�&Tӭ��#�3lL�pq�D)[���n|�m�ן*���XR �}���=��s��R:p�^^����̽���p�{A�F��n�'৬2`�����B��i�҃��y�׽ �����Rb�D	�Rŝ��SuKǕMf��"���I|=��%X�]�L���İ�т<�ه��c��(6�"��.�ߡN���\�cX�MJ��B��55B�d\�y�a��WZ(��{�z� �a1���9��U?t8��=G�xk��ZG�:�X�.T���r��KkR>C�4)]ТA�P�u�4�9i��i�����Ǫ�5�15�`5�g8P��
v0�8T�]@�#�����3i�3�/K���:��PLEE���ao�=;��/> U?$ט�d���j�v����H���K��gl�]�h�ŶwYaVq��bү���Q��/�Ɯ,뒘F�D�Q�_
V�%���W"dwcJ�Ӌ��$\�߽"8uK��bPū�1W"375V�"�VA$L-�1(�[ɢ���r^舻j�4�ܗ����͍9�7����\Tt�\��FU��W��̝�s.�3�w1 �z���J5�W��L��W߶$Y'���{�C���)�^x��W������A?~����)� 'Ѕ�)��Bω�K�j�qp����tD�0NiÑ~��^�O���w�G���m�Ì�R�~�D��S����ғ�ɛ��f��oA��n�&��9ո�k�Q�<��o��¬��{i��q�*��H3�EI�$!J)[�����Y�K�	�s�2�`{/����
#}J3�83rM_Z's���HJD;k��HH���HQ���t�!A���ם��C�g(�F��>���S��Ӽ-iZ�pm���� ����@(��MU�����]�����)��^�e�"��]l+:�u���.�{Z�P$���Tl������aM]��hZ[m��� 2���Њb+�2*�(c�A�[��(SdT1PQ�BPQ�QE�0	B ��a��O����������}�+�Yg�5|�g���I��?�m���4F>%��ܜH��=�Bh;�ejmY}����7/��O�[q�됪��
n�lP�ԉS��m�h��ڛ]�7w�dk��׽|\貴�Yd��U�@���-j��C�e⠅�й_u�|28�|y��S�}s2���smk���e��:�rvHTy��g=�/��(�ʬ��OŊ.�kyw�ls<ӫ��/m͇c�Hq�j�EG�Z���lֽ2'��o� (;:b�� k�p��@�vߏ9�#G��rx�6��	=l�B�'��'aS����h������8�s���M��`hQ��J6�J�J)�1��l�D��9�c�qv�L�����������ϭ�/v�/�r>��i����9�F���bi��%�zƙi	�������f�����,fgm��F{4�[�$����wD��ԭ-j�Vv|��\��ݦ��.WC[���y\��[��_p�*߼��ě-S�����ܤJդ-�E[��Dq�X>����L�;�ې��W�<N� ��U�yZeg�ޕC�[�
����T̏���7��h�f?3-|��@�~뒔v���L����e�s��=��1�{J�Y��U��AZ�OK`��0�i��EO^�������l_�4���ͻ��E
:m����s'ֆ������ZG�$fc����O}��{y1)\�%��{0|��&�`�y��Wɜ��6�:�z���d�o�8s��0k�k2��x��s�ܵ����6-Ky� ;4SS&���,�^殝/L�����{�%jߩ-�a�u:��ȑm�ʛ♃>���9���������^%����T.���,¿O0�;���Ж��33EPĞ柯z<?�2�=s���v�Ѱ��<U��"��Q*tXlp�+۫��4?�!D�[�6�Ŗ**�}_w��۝��RO�ދ�i~I?d�Ie��~v[2כ:��O��i{-�Ś���}i����u��p �_כk�����O=����/�&hs�ν���}jA��p��@Q�v~j��h�1d(9�;�nBU[��T���nm9��7��`���#�ˬ��]��׾�������pq�Hv�ýYy�����	�l�W.�E�8;cWMҽ�of�w	9{~�DŰDf��~r�~��!��y�����u	�Ԥo�b�;͹{�_�7r��{ʾ.����V��Z�t���]��u]4�^q�`70λ�og]_tF������Ӆ<��;�.�m[5�8޽'ӣ��2���o�.O�jf�0P��)Ӎ���C��'�L�~j(k�}�}�77�:ER���~���;�s�����ǜTr䷩��F\J�T�ޮ�����-yS3@���+cͮ��S�N�8�q	���5{�G�Ή�,J���4�j�T�v�"��U���xV ��N
\���R��&l(��Lz�hUJ��#���;��O�+�3U��Q��K�yX�|���!-�
�ڱ�'jS�g9���>�{��̥v��q�J����Ɨ8�֮��`���_u��d��>���gpx��+���\�l٫޷��dC��EL��5������g�n�����/��uM��ph,�S���+o�B����qM���������vA�o�dR��K��)���;�|���t?Ns)���p���;.<��z/��i.{�+�}y;�7���~����<�bx�^�H���r]����.e!����Z��4�8�^�tk�I��r��v����mZ��z�K�ք�}ג<���潡Nm/G��-ͷ��o	���r��hΖr�K>o�s��%�ʉ��-�Z�g��l��q�~�K��ŭ6���s���Gj؄����)I���Ι����)9�)<14��z���ӷ��}i����]y����H�H`^H_E��D[H_�&
�1���Ɉ��iZ�;��o��~%v#ʚ�$� Mя�2����oP��m���K��\���/�~��˥�w/��qBO,P��d��OU��|;���Ҕ/��������Wj�7�Y��/���՗W_^}y��՗W_^}y��՗W_^}y��՗W��yu�w.dK!GdJMA�KS��{�2O���m��K���.�k�����?=PY~�ǻ������!L�����wk�����k����oB~:�����L���Y�~A�����I�Vao˴�̷Y)�)m`�]��qj����}y�˛_����7�����/o�?��?���&?�3��x�3��?z1��]�$��#����X�/o�������k>3OE)�-z"���g�������շc���|֧zr�����8E|�Siy�E�vI ��	������2�DԾI\JO�<���k9t�,y�����p�h���s���Ѓ?�Q�"��C�R"�PI�\6�(�<"�=���g��ѣס��m����z��OD��&+?�<5'���[Lb���;i��Į[HE7�3{S�<:�^���i��m޼9+��f�\��Ku�&Bۜ����N�/�8�$C<xO	]�?���"7��\��g%2�Se��hk2�������n"��ۻnjj�[�siR�C޶�:2N�Nh�:�?��c����+n�W��}p�$�������������Θ�����T/
]7O����p�4鈕���F&��@�/��Z�-K7K�}��.iߖ��Hj �t�M��;c�*X�l�~�\S���ay\$���br���w�����c�}"�1A���8�����pKb�[�1�R��M���J�}��t����oi$jW���g�E˒���^��[D��Ik�=������AcHl��U�Ħ![E�hS���h���2�g��y�s�Qe]�(hI�1�1�q?7���W�g�Æ�>��W�|��pV���^!�m���yMϠ��իW���5�˰�+z����n&,>D���FE2�M�pd	s��1s>���<���tK�pw�@ø����4C^[�*�~ല� ��Pu��}������"�-5 D+w�6T���X9�����ACiP���;88l9ED7�w9,[�E��E��2\�Y�-�sr�ख़,~�DTم[��[0V=K���z?`�}u������-*��*�ΰ�.Y�c�+�M���R����g���g��/��u�~P�囦�2D�	=��,�4%x#��f�<�W�5�K�|�2�y�񨻅��s��!�_�f���A�`�/iPAN�^��ж���$B~��P�/o��L �B�b�m�&��q[kk�E�. �,y%z��U<Wy}�3d��eFKK�VQQ��	�����p���_^0��C:�W�V��߫��<�E �Й�}3)��?/ ���\ ��2m�֣p��D�U��aq%Ae���8����!e���A)nO��2÷~z�����������/�C�e�9ro���x;��t�ޞ�@�{���M�Y,��k��̹�*/J%l����D�����nT�Bui�Hӂ��|Ցp;&���KH% ����ew�SN�*����-(��!��K��Nu���.#c
p�uIII�	i���pDn;�&�Zl�i�71�NH�W�~���l HЍՓil�v))/��B�4���(�[JDK[\���m�oVf���3_��	8 �ն����7�.�$PR�����ϻu+���D�)�%�
�]�?6��;*�T�\��>��!@�CDn)-����@0����gW�^m*��,�#h)����p��❽3sD����Ÿ61+�|�/%�8�ŏ�E�QT�B�܎)� H�{co�-�%�����'r��3X�O���(77^� +��řC���g?��&�q��DW��g@��h�P9�)�-3v{�;�mZ��v{5튗�ci���UQe�D�7^ěj��ڝ���`V���Mgl�WDk��R�j�cuzL1,�+KO��j��}R��g��sZ���ۏ�22�#
5�!�w)� en(R��f��Гu�?��x{-~�?m,�v�l���b���p����ɪ�ʁ_��|�r|%���&�}b;����:X�ܮ��y'h�_�݉���yB�(�����񴰘G&6�+���,�!B`c$r��Q�W��Zʒ�y �bD���V��+?��͡������7),) Ȋ�*{	h?4��$���o�=+���޶!�o��8j��k�!��W���S�� �} ��[��m�����
kjfP����x�X�;��Yb;����I/@$���.^�i�A)��scN����̘9������"D�_���9���/�-�R�[��r]l +#rǵ�^5)�!�V�,_y	�L�������N��>��ծ����;�-h=�}�X�R��x�Xg@4Ʉ�N���X��!��*��M���DsCh�^�Kܜy�Z	r�$�4J����B�22vh�g����U�"Q;��X%��5��AU�e�9)�D�� ��k >�����z�F�N��u0��B;���� �ʄӕqT  ˣ�v�yg���"�Qɋ�:��ٔ�Q�E��c�hY3;�n~�F�^�<9��K��4��u��E+�5�5�u�����)p�d�M�)��׳�3��Aa��W���5���H=7������4�؝�O��>}*SUQI�D��a��iYY��tT⨶��g�H���jK"����f�0��P�ξl�΍k���y@d�|�ȉ�_���IM��=k�H�r,��	<:�<�,9{$"}S�����+-a�6���Y`�^���X���
k^0�x��#��0�1�����C
I�~,�l�%�
���n��	E��Ak��1Z� g�.�����PbČD�4%����G��NĮ}{�X�����y��%�E|N�l%�"�)���Tu��ح�|�O��bQ���Ot������������c�&��?$���[��XX�D �WOں������?� ���YS��3*+�EK��� *+1**�sx�$���&Q+��2�$�W���i�풱���ʽ�!���^�F)�����m�P��u��G�$�"#��+��(���BX�$��>�z�{� K�� ����	�BV�j��ت� x�2��#@Q�o����`e����xG�:�Y�Jeü��	է�#x[K�6�.�>S��X��m��$���E��%$�猱�����ߟY�C8���ХK9|F�j�@~˽�$,
;������l�M|W׿�.�������&�A}����زjϞ��2���p�a}i=	c��o�v��>�X�ϙ7I��Ą�QE�٩��k1���oD�w$�͵Khx�Oi?��ϟ�8yYY��;�x�}#3p}�J�tn}X�k�����п��HƺW�Q�_��%���)�������f:���)I���������r���LE�!Z){��p�X�_�r`)��4T4�������������K�u�@9�U�dm�(�`��i��4RY ��3ǛR~�ʙ�����ދ�p���x�;�)3��,�KU���@`#
��ƅ"��}a��^��˭_Q��3g΍�V����~UT�&̰�> �q&����7n���,o�Q�o�3p(ח��Z�c,�E�^��x�ňr b��m��>h��]	����0k �V����y.�?6���޵�n��૓����y������0�	r�.,�Z^^�.��������l�v��/�����	��e�a��v���(h�\%o��9ɧz�����(���tJYRkZ�1H��j������9 $JPe?pL�M�@�_@�\� ��6[;9���k
�D�Q���3snu�����%b#i��c|�q�G� f�N���sXfN[�~���B�� �JtV���|N��q�?9�xɥ�˨�p�v���'�@ǟ"��V����ʃ�1��· $H���k�5�U�s�>�l��Ǌ�8B�K�^z!%�!vV���BA�#h�^�i:���s��5Jr��_�e�X��!E�w�Ct��t���:��1]x'����8w�1>�:r
m�*��x��/�BK���KIl0M~��f���	+�x��g	��o�S����	cbtS�'_+�!��$^i#3fsH�;���j��b5J��Ή���"�C(|��fl��׏�:�DԠ�?>M����Ud�U�!>G�'3�x2,�� 2��!S������W��Y�X�V��X*�9!�)[p��ݡ�i�SB�YgB��8����WCͯ|��ٳ�V;��2�xGGo���ԑi���d��J?R�� ����2s�B/Y��s����y�JW�X�?x1'M�T!$�m� ߬A��O���y��R�f���ި!���z���Q�C*�i�A������'�S-}m}�"��B��=���<U��o�
���ȡ ��Y�F���h�x�3/4�g'�Xi)(SF+�F�K�ĩ��8����  �`���Ϗ=��%�{}�@~;-X��������
iT���2��]��cn.䭓��ݲ�-PMޢ Ʃb��Os�i��
C��|���\& (���6�*r�m�Q讁�:-���9id��"����w� ���X�7ۇ��كB�1%�J"�g��R��:	�yj�T�Yy �]��
��$��	5�9���J�1Cyk��;�y�o"�M��Ӵ�p�]d��9���O�рG�'I8�I�-��A�J�`2���ƣ���۱�L+�?��t������)۴�u?GE�q@r�¡0F�K��y0�"<ŭ �13�ʼ��k�Sf���p���b�#+q��r�� TZ�f�O��v� ���3sn��\�Y� �.����s���[PxӮc�\j���RԐxPN��Z�k 2uE�\��v�VE�vKu(6�z:��F'���L}�WD���l�Ӝ;Ϙ8�,��{���
�����o���ݪ Oh�u�^�n��O�'x��}NA�~ϤAM��7��� 8Ib8-{Թ�b��c�SE2"9	-�=p��
_
�/��4���-���E~�\�Y&xdV����"
Et9��^��Y�e�u*��6�Z�	������j�vN�0J���g=<F���kP��b;�LM2&F�C/�����	��6�D��{D$T�
:��#�i�s��Ȣ a[�wk-��?c[�#�5�+�!q0��������$����o��.2&����?\�z�汧��~�ƣ	��b�K�H!@%��$3�>&�X��fnȼ���IǍ���ޭ+�k'���S�ⱄЩv���HF!(J}�GǾV�ZM��>x�ђ��;��~�Qil��1,|�����`$�u�K򮙹�'��J�?∝�{$I킶m���`����#wza��~�}�&	�����W�q�S8�j�8�V��S=�y�vd�|�d�$2��̢�R]�cP(u��|����'�q�c��g\uYcӳ!��)����Og�+n�ZT�_v6�%M��Х��Qb�L�~E<�au��ߊU99�!95ɪ���a���8��m��V���E��S���� ���I�{�ә���8�>�$���E;h���a�OTYW�ObBMI�\&*��u ���f���\x*]�i�#ր�YV|^��-3�geI�&�?|���'�>�Ǌۮ-E-Cb,�;��]\\��&�S�r9q�[��Y=�:ۊ���Lԧ#g��d,�4X\	8qA�TTY������qMd޻Ȯ��
Z��dyRR��2d°�Ȅ_h?}����c��q¬��A�"g$^i6�
��K'��(��ޑ�)�����|,	�@��kwm)��nP`2233�P{;�ǣ/�C���uH��n���TUUec礈Z��2���yYء��$1?��YL����U����z�V�Dab:�^�#\¹4��be�m���R��@�]��(hF��JD[ʔҕ&�h�ÒQeC�);Q�$�����,�9uD�u�f̃:������� ���w�7oN[�0@l��������H��]sXy)��XZ'�𡶟.�����T��N����J�*��?{H�v8��^�N�"��=��h�>�F<~sk�ʂ-ʞ�/^���ʚ��W.�
~)�|Xgf?,�)���e�8� ��8<!��g��1��̊ �1
%�;�
�xC�U{4��?��Ђo�9�Og���C(NwJ��#Gޅ\dp+��/̜l�-Z ���J�6���a��d�� 3,,��1��5і���o���'�Cv�梠��?����$��Ц#x[���Y@ouT��_���\�R �מW�,ʘ�m�|�Q=�\ҿ�T��$/D���,�u�4��\g;��Q(��)�QjE�K��W���tf�%F���_e���us|�}x�����Xm����W��b��J򠏘�4Xx�ر�_Ѵl$������D�S���Ř�kʴ?,(�\G����i�F�㝌����L�<ʚ��k��dD�u_����Z�%d���c�Eր. �a������ أo�|\ǌ�b��G�Nt6���b����ֿ:ˌ�}��#|ׄ}�L���<ب���t�/� z�i�m�F���~0܈����z-w�\N����T�{ǧg?wN%�1���J-?Q�`�G�N���FK�����7b<�P�M�A������^��\�C객]���*�v &�_[#ʺ��z�����1q�ݻwU��ad�}�+�qX�}�I<EGIA�$u~��װ��&(U�	�<�H<��_�>����3/`	�>Iq���_����3��[3!8���C!�U��#]e	�	UR��U��nD~	q~)��
n{��N l_���u�9�(��x���K��wiM���o a����T�5�+��P��}��	V�-GIk�툫z> �P�z媉�/��%�!�-(�� 0t
�����GQ���O�+4�Ϫ�A�C�a~��몪*E4w���е CE���o�I��!4���:+�� 0�~��d��(c�9�&%ň�-��Z~��1���G�t��m׃��a7�N{8%�5��R*\%�?��+���@�}9�gb61c* �x�*/F�$Q]doŸ6���ǎ
+��̭��:��\��:���^�ԾȐ��U�g_8�
*��:2��AČˎ+I<*��Z�"'��/j�֏���B�2���(n�Zch�|�*��K�x���D�R��#��4M�d�#��kkʄ��b���_`h}cu�� )�߫����sEd1<�W���OAg��v#�Lau����q�?�@Kv���i�-���)��ege��[�U�`������6��<m� vSq��֋oUP$��lK�ϓf���V��Ȓ��#sss���A�[�7��#���/,�ӳ< {_4�������Eʭ1e0V7�[�)]�=�@��rUh�.�:�!�Vy�wK��D�g8����̜3+��-pe����`����� �A����QQFEM$%�`'��<��'���u�D��m�W��}�0�mѐ�����i�ԅ��`�%�W%u�̐~V|B�[f���I`��8��\�h�H�[�:L5=-Pd9 J�=�,���`pʥz8��[�>LV"BO;:NI;�����:!��,u$Z�-C��}���+%JXt� �y��2(��Q�є�h��B�R�1R��須��׮���}�ە���3ێ�I����3 ��� ��Գ�
��<Q:���kx�K�;s�LinhJ�[GJ<xp���쟌�0�a7�Xz 	=B�9�=�픒Č6u����Ð:R�����'"t��[M��
ނ �L��K4�"g�XsΙ�Z0��p�m%�R&)wլ�Os�5c�j�>R&w1.�F$P<��_[S�䟢��yk���>#����~=%7w_��O�ʡ�]y�>F"M���a�T^|�>��8�RH�~5/3++�ִ���uS�$��`��)��1�:�E���?2+l��Șx����3�܀�������bј9��()�߄1�9fD���v !�׹�	C^�n�;4��m��)�����n��t\��1>EdV�����P���=߇!{�G�������.'Ģ�W�t�s!S�Q
����cd{n=�Sy��Ր3��uT���`'����������D�y�_�CJߋ��?��P{�]�*�Py�L�t܅'��@}qR�����Z�i>�r��;c+�G���\2�$a#N�G	���`���9-�y,��/�1��v�'�e�*��
�h`�X)�����</+�����Q����>ϒ��l���g�����!?�n�٧V83� �'���W(~��Z�s�`d�u�A^�
���,>گ>B�Tr$�L+��~)<R�GYp۹AAA�(r��E�j`����?�T1��k��[�Mf�5�3����;��A��.)�ּgfК�P�Y����Ϡ�SYrvY�E��s-6vo���vx�絎6���T7>��^��Z��{&s<�c>��f>�y�PUEE��;��(��xVC��:RhU_P0A��������$⃨G������.�)#.B��:�Q^�l�
��c����9`	��cS�2?e�m*K"������`0�>�?��:��w Eb1f�*<Ƞ%�s*B͖�2�]�09�|���
l[�X�q��}�����^�z�F�t1<H&� i(:�������E��P�4�S����z�f��)N�{q閂�לɵ�.���*�;����J��Sr��0Q'�r�cA�bG VsQG���
����L�#�ŷ=H��2})zC(q��uf��J�ݘ�b���΁.k����J�6+G-�f�e�3y��1*����JD'���uFB�d:*@y����kP�5a���^�\�p:�]�o]�,��ɿH�o��6�#�\���S�6�X�.RS���d�w"1z,�V����k���h�1P� �\F�*k�w�ތ���NK���z�6FG���~,؂���QG;�Ӻ���T���@��Vw�@7����;�7��p�2v�=
���a��ۚ:��������ف�X���e0>���^�da,����u�9���� 7;k���J�x���t�,���sC�M�݃�s�z��ix�Q%rV�&uɹ�r+~�mì/̗<
Qހ�4����r��o� (�H�R�?��񣖆�F�jj��U8C��G�Mq��O��e	�M���G�|�/YL��ŀ�2�)]L�<��2��N�梓x�P����T�B
t%�3s�H��������7b���>p.����*�6�otLcYr�DR���~TT4���2dI->�@w]r�`��n�(Z�斖@�V���RKU�pwI��ӤqBB��ȞF����,<���u=���;K/&��F���~��.ߝ�ؤ���R�*L���8��nd�]���q�1��Τo3L:ۆ�cH9[�ܝ�ױ��"M��:��a�y��<�)yf�������
���3��⏓y����t5>m�6O��� �L�ݧ� `�_�K<Me�#��d��d{��"�����M�w�f����0�����M&*�K~$�[�VdPi�/�c�@�_dh� �2s�u$w�]�w
[g  �:i)���Q9bLGÔ�o��D��9�q��� k8n�x/j(��Gw�:���A���ۋ�,�\]�c�mD�t��o,lP���Tw��0��6���dצr]=]��5S����$Ui�n�w�P���_��H�SO��x���7�%�K�0�V�^�����׫V=_��ę��7�ތd��~%�����"��{|jq�Wl�����ĶA�#]�4�	���(��61M��'O������8�ba1>� ĺ�*t"��Y%A�4|C;�c6�t�����M0��]�!|��v�-xP!0G�eX�i�g�?q���i
}�Li������̪8O�e��A��X��g���Ǟ��F)lݪ����q2�^��l�)06j��r�J�y�s�o`T�1�׳��JSG� ��b��bv>�ϟ&�p5[o`a��L�JF�.l82!3q7J�),��*�}\����y�hzv�0�"!}��Ҡz8����ݷ�p,�KȜ &#c����&\H���0Nr0w���"=�VVw�8i�b@
�m�݉Y�q��X�m*��O�5��VW�o4�F�e��r �+���$=�����
��3��έ���ȥ�Nk9aSSS,3��	��f�Ns�86����Ү�����1�U=���'��rUC����BG{ߙwӓ��s�:�!���%��[�-W��2ʰleUUfUuu�/�@�����! u���܋��L� ���j�Z�P�`�Jy�����ׯ_'U�$�=x��^ۄ�ȟ��.��k��ڙ�;�;5�_JQ�ͳ�4%9��]ۗ����� ,Iwuuu�����(iP}�����"��p�s��eJɞ`$��
�d�bU�3����35��v-�ٲeKe�OY�]�么"���[����j/
��B��5��o"	}YM��A6�rK)BS�P�+s^Փ��S�E(�|��
gy/��g,`��o�1	;�/�a��O[#u:��D��<r{�;�^m+;��?�Ճ����/%�u���о�{G����(�eUT�l�ښq7�j�q�^В���8� ��j0�
�a�0�6�K2q�q8K�����K��)��>(HN�%A��v��)^b�B�[M��,TUPPؙw7�ϯ��cV�iu���4�>�~}�%�D����� ���f�{���>��'�0�:��)�:�25��G��w�.a7�}C(u'w��E�z� �,�z����e���|��G�)/Zt��0��X�>ۆ���W!5�
�$��l�?D�}�M�z��B����T��I���8�'*C�����z�Yb 
u���"c5����s��ˮ5޶\�ޙ�����jqpq��O���G|v��mk�LP�f� s�U �P���;d�0��ka� ��]0���?!?�[p/�ӧ0ȸz���aH(>��m���Ͽ�� �^��0��Uc69���	AE"|16o�Y���d��h���R�^����W] .Q�В�-� _��qP'�E׳(�nI�꧌��e�̲�D��@�B�f) *�b�����������O)�12��󇰨�d��2���T\-�J32��̙�cL8V��q���"C��F�*	����7��t��tC�tVf��M�|�"G�377w�-�G��5����� 8�E8݈(A���x�4i��vڡ��}#7G����Y6�����N`>r�ǎ��\��S�	v���~8���w�(ۅWm,_�N���
h �q�4�/��F���t/�3	e~����[!3"Qҡ�v$U?�i�ֹ���716��:�$�A>R��SC����Ū�5����W�ԙ-}T���o���|�����z[6#dk��O5���"����H��������sĤw�E��oC���I�;|�5̷��ѧ�ڳ��M��k��yI ����T@y���K�c3}}}��U�䩅�<�ga���Ls���Qg;+++��r��8_��pX�~=u�л�D��C�XX�w9bd����.A��F�ڰg����`�sc-Θ_--�6�:�e���^;������r,��>��y�����VB��y�LC}���x�eGG��1&��Rv��i�7���x��;����?�,�W*�FG�Y���l��y�
�1��;>�8zX�)��$�{7�L!%O�J�s�ςjbz��{	ƫ��)��d�oI;���,���N�5��BAp����\�+�:��:VB���D�,i߭�3�ԑ�gϞ]�:�Va�Sz�1$v�"_&B�kXs��I�|��h��=�`�Z�o(�VGO�z�q	�OKZ������o�������:9��,�%z�;���ob��3� �Cǲ]x�"��d�Zd���}(xE���:��ͣ��;J@�}�$S1����9s]z�z:3��A�7]i��Y�3;̉5I�X���tP���#�Ģ�I�MzP����W��R��AR�333����L��������x$�*�� ��^�Պ)�O�w��Y�����`!����^ŧA�姡��F~�+���M� �����?�c���CJ�W��h9@�7����������d�c��@x'���~��u@�E�M���ɫ�_Q�-��Um�4�!�Z����\�^���؍�r�@"���ȃE����[X���%2�z0��-�}d�8f㎸\ޠ�~�a�)Z�(��,|��07B�0��X�_��1�
`ǟ�J���;A�<M�>���;���=�+u�/l*��l���	۲B�<�������S_��	|���^?66vU�� dD~����Uw:H�w�?��b$7�4�[`t|�͝P���U�7o6�`l���=@�7��*�~#'�lG �Ӏ��VO^A�3��>$A��L v�sF���YFՐ;�O�ܡS�����ɨQ�üN����Q!�y����kZI���	�i��.�/�0�ȋֹy��8\�UQq�I9�:��:�
�b3C^�#�=v��E���mca�R���m�9���[��*����c��K��JKK31�g�������t͑g��H�> uX���<h)�ؐ��d�z��aB��7{7��M��A>C�xz���f���Qбj��hx�<�W�_dh��?Y�}R6��6�{ hh�W��, q[�㗜5�To�z�� t� ��M�	��Ѧt ����3�:RpP�����}=>L��N�- �{QR�9*K�����3J1���0VOޅbD{U76�8p`2v��B�7�N��?}��2u�:4�����ZvVm��V��oA6h�w<��uv�%�N�<ٶ�T��K^Nt�q����,%�+Թ�U��3�$W�%0����!{�@]�f J�R0v��*///'Ї��8���F���6$�=0:�+\ɞ��ѐg���A>��	7W�JK��h����	����L7X��3�L�g;�O7����q@+���wyV�ú�t��@,)>�������H�򧢼��uK���`a�ϧ?��D?؜�ρ]@̛�v������c!��Y�3�<�\f��.� ��o�# Cμ��dx�����㉊��U�j7�pQ3]�\� d��u��"�XvTvȹO��H�$a��!���ܺ�7��eCrT�"cc�5Z�*�"�$F7.����ʠI��,0i:�6"��������r��B���S �::�i5/Շ���6����(�D�T�U������ZdǇqCCC��	��_��?�w�)�{�Z�J~hʁV����6z۶kjhL?LuC�PZ��`�L���)�DUP���!# ��h�>��V�wf�`@󥺄�����:�a�\s)q��dBF~����X�R=LDpx�����L�����6���o�ԑ1o�Q���6��6��S|3�B�j�?(U��1���|�#G޽���DCf�mY�o1?T��4�Y�r���g��� ��Y
�����8h�����Ti�I�x�u�!�&�e�����.�V��a)}of�8 �΄�*'	ŗƌ�s�C�iK�J����r��!g�g����,~�Niu$�r�u٫���c��-� �y##CL����i}�DYHd2��v�� �^ja���9���\ZQ�Lڷ�i;4�<F�Г �q9�����0~�e�gj���A}.�ǙZ��V��ToW��� �O&߯�~׼�1����v-%?�tN�Bۉr��f����D;#L�(�#uO�K�'��i�6��)�K��<�8�cf�;2���-̱4�1�+HQ���n`�9�Ȅ)�oZ�} 7*�qG�s(��7��&)������GR$�����������O���>���w��r���6��i���u���JB��ώ$d��ǀ�����Ԁ����PRn�In?)*�E��	��p���=�x�5	�Av� ��/h]���c(U|X�aw�r�4�O�,+q�&�wy�S�s`N�&���e� �ƺΑJz2�y)L2)[��n�6@���*kj�O�4in��=Bv�-$���F	��� Y�8��Z4�n�m@5�̡�H+���	�ԓ����n�L�t��[�i)��e�ھ{�޳�����h��t�Q=�EG��U(�ZXx�5pT�-�����m۶堺�Y�<�u�݉5��!�Є+��O��A�E�]�'����X�x�aH����^ۏ�k�;5�jd�1r��w�Z�MO@CZȚ���P<љ�y���+��h�V��. �%�[�I�5�DQC�ײd��&���z�A#�	�K.�#���3Ϟ<y�vp�;I�R�q��,����D�[�y�:it�՞d�c�b�uf߃��(�򤚢��n�Tt�#u����b�����%r�
w_X���w�2r�F�ҫ8��5Eb����ڲ!3#������70�ؘ��{I�*h��Uy�ŸzrL1���yTsȣn��>��ֽ�Ej"^���p����vD�K��a�\gcB����YWt$�ğ2���gd�l<�,��jg>�?`$u�V��c��ܒ�V���,����9S����f����h`�`��Q���ͩ��)��<0�܂�Ў�=ʱ�Y�usW�^M�+]ۊpF6�nM:�ҍI&�Y�Y-���к���u�%�Gl� v?ǎ��-}�������D�mп�������)�$�g��>k�=M�ํm���dD�Ni{,���.�;@����x ��%�u� L��
��|>a���%���@=�Gy0���ݢ��]�ϸ�)������	4��!�-��8�ˌ	M�3<�Sr$�{�,YX�j�|�Jo���(��Ͽ��4JH�|���E]�<��8;�Kt'����e�WѯH�;;��$���|(Z �8���H���r���{,G��2D��tu�v�r��e��,u��� ��0ژ*��Sv�Pt���l�2sKصI�&�;��n����$ Ey�;3��|	J�1d�����&�o�]��(t��TQ/FO�n��f���_�
�ԙq�>r�l*3��B=�Dia�|{J�$�����Pj�BKآJX����=�J�}��CY�=�Z�ZE���3��뙙q��^Z'�<�ɚ����vm&W>��	�<ˡR�Pȿ�*����ɕt���݌���a�XǌIn�W+B������ఈ7|<��4R$�I����of� N�B��vV�B;*���&w�4��uf� ̿M����RR��0����u��=h-�C��C Æ�'K�T�BB��&�j"Nn�=�N�L���T������mu�֠q`�8k ��-���)�q���8mI��`f��r�г��������u^��[L/������F��RFF�u����9T<Wj����"D�>Y�d;�����S�2�y�S��KF�
�Hw$c�b*��Nh��2�r;��gz֡�ȃ��>ة���g[�h���@B�")�0MC�����zw+`���B�!ؐ�'%O��g�#ϑ���@'�s~�k�F�`,?O�l(`'��_�R���r��ݷ�E?Q/'}*M#��慰Z��{r�q�w��^��9�c��R0}��4 o�P�:Z$�y�1a -��1����+v@RdP����xĩ�,#�C���w?��82�w	�����n�d�|�����T��S�d$EB����y�f\�+��|a�^{��Q
'�{Ӭa�jZ8b�c���3{7$�]B� �Z��]/37��d�23�gg���1��sR�@t��T�5D;�u�dNJ�ϻ^5+����u�y���.,�L�"[� ��B�<Cܨ̾�Y]�<-D\6ɼzXX��km#:�ƍ���vn�>r/~ރ�Sd��Zm�x?�s�l3���d(�6(�Q:p,ی���e�/,!��l"ET�&���϶�
{�J1d8�oñ�d�\�9Z���q����$ _ħ��w��}�����U��"���W@�Ői�0L��!�Ts�t�^���PCN��ɑ�E��A^^ֽ{�W#�Tj�Ni�����-�Gӫ: �H*,�\,
�tm|Lʭ�����H�WF�A�n|C�l �	<sn�ؘ&�d(B�K��؝��fLu�K�f!BAkԩрtD��<�����f�+���r��nZ^��R�@�n�NLYN����ت�����>��h\X�����E\���?B�JI:/P����>%�K��9��ƪ&G跼�ϴ���.���g��7��n߼J�F��ʯ�j�?���U�%��/���~o�����ħm���V��vm����k���S��Ǎ�iI��S�n�3��������} ���/Z�(�ǧM~�+��B�/YQ[ŌQm��0��r�|���Eb酐����D��4|<:{�A���62O�N��n�rwj�\�cj�+>�KKP���;�y-G�'6�z�i�D!Z��X���=���K4R�A`|��GJ�OL��:khh�U���y)��H��ce���d 5��_��@�rI��� �Ϛ�t���D��O�}����&�.�I<� B���~�H�~wn?#����������bb�ҫպ�ۑ��a�(��z�� {���5��Y /���Gs�� ��!�ai�W����w�UD+�_?ņ_Q1N���"/�MV�x4����s8�v�A����2c���rs���3�Ô��wa%s���N� ~f1_;��������)�C���b7]xE�'�S�-����M?�Iou|���[��W����]r!P&�4��$-��n\�(�����~~�߭��jL>����k��j�Sz"���X�u�4���	ݯ ����W�:/@i4��d�PB��ĉ,S�6������r���s� Ȭ ,j�i*%���d���6?S}�i3/�Y�+�\�3H�<���c�^i��V�imZ�#��	y;���t|��c���,$���uw�H��;��s�u#�K��ў�h7}�W�wHZ�6����Z�(|`M	�<h�豈�F�>%;�^��/�?a�o�9�wEj� �&n�,��~�h���q��u᧟��s�U}m�R�V�-���H�0�{�u& g�nbjz��3����d����s�a����:��X����R��/���w���v80���9�)�Ȩe?nf�����H+��X�bV�l��$W��I��Ͻ��pY��=Ym���!�.�0j\�'��f�������p٪��U�5���^=gq������T�ﾁ�����+5&�R(���0�*T���@TΘ�p[�	�=G�/�8?��j���~�=͊>�kw]��M�u�L չ50gw�4�8���C�e��j��i�̘�ͳ��y#��,�ԇ�`>W�q�9q�R_���>ρ9u03��7���wã̘���VR�>��WYW�ԕ��CG��BS��B'Z�� A\�������Qv���T�%�*i�eu	j1�b�F�Pq�@A���(� ��u�	�>p��}��ܳ|�;��{�O�X�P?��t�I�a{�Q�~?c���;�ˊ)��ɍćtV;�.��f����^���:K�t�����B����~d~ӷ8WB����ΡdH`�]����P�+C���qYwMdz@djw|0��6t�իW��c��0���R��G��FP���oM��mf �EY��$�Ō�Kc��Ż���9���ݓ�b�?|�Q
�_��V�:PRb�pH�ڧ4���2G�}*��2����g�������V�4�[ ����T"�n��F�C�36C��� ����ս��k"��-L 3H@8�/�s'S�X�]�"!���_�	Y`�_MW�,���\<�F��cnl!��ʣ;k�GD!��s'�ȑ#.�`���� ��R�=^�`l��~��P=�}߄J4v�\��y�b�Z4��D��0`��o�gI���;gŻעmR�F�;��N����JJ��ΎY!�e8I��è�ą���w��G9�V��_�ݶ���Ũ+��]�e)v������V!�=�n(<�R�#��h}��Դ��䌞�wI���$;���L�:d�<i#Sa,VnaϺm�H��=�a��T{}#�(r~��oo�| ���0;�����k�M%H:R ����GB3��Z����8��Q[�X�W�mh��%1Ke���q����;�.<y�u+ڐ���o����=x�4����.�p)�R�xW�����C6p���uO>[�Z<k�c���#G?�o�o�D��;�*��c�I��_xR��sF"Y�v�4����{�>�! �-_i ���˪�B�4�R�5�M��k�e���Q6�.���0-G._~T4v~�W!���m	R:�)�r�n���������CXMҏ2O����G�pj��V�Z��b�]��`4-����?b��]���Dtj�P�<2]��U�-���;gb�Gr��(����W�n,B�bKr5&=�y6����I��#l]q����R��Z(���-z����	��� ��{��LUe�f`kB����O�)S�*�x?���R�NEW)���^�♼N���ܯN�v�Z���S�f��.b� �j�Z�܏��<�%���r��`ΰh��yUأ��eꖑ\( �u�]q�E�@�h�kj�9��41K>	�n���Ӎ�ƣ,)[�����^�_s�j��`'"@�Wmp�]��b�
(X6z�����՞]?�A�0S�`$|���Vnܛ��8$�I�S����\]�O:1���!�C�7U��/w�+	δX ��Kt��ء
��J}$��!���B��k�bF��q1�UEEE�h 3iN����JM�Ʌ/�2l0��r���FVW�k��L���Qq��l�n<�qCG �7ۡ��?-..��r�g^�u�Ɣ|:O��HP,^����~���P�>Z˛~��JQ(6��4����>�?���zo1��O[���t���$	V̉��e�a��i:�U�� RX��J���ܻ����5�*����pLB)D3k�i��ZV�ד�COq݄nU�Q��Z�x��m�i�,�Aޑl��.��[/�r+�j�|����p-k�y� "Bݑ�a``��V7�E�;(�<|����
�jl�@N �u�Z��@�u���`��s@�by�y@Kl�b��OԿ�ܶ��r��l��'�(+��O��GM�%���9���-j1����0�������Q��2{���Y��n���3� ��Q��.����yyZmc�tҫ��wbO-�A��"�kӚ
�9�+���&�����}��a}�@����4�zTep�fT�<��ď�w�ܳiS#�9lQ�p�|3�*��#7!�n���0�s4�4Å���y�T���qu!hߔ��Lk�}���ǅ�^UՙS(���^���|�x7��U��Wr��|A��(�B������ၞSvEy�ט��S�?���ux�!�-��GW�^$A<�&�Xxy��XKol�A��T��!rFh�y�k�:N���o.�@��1E�����Y0R��H52e��S� Ъ��xҟc�qM4���-L=�%AM^<d������������l�T�hg�i��'�H�	^j�{&�^@/do�܀ :�t�Pg��2 �6#�%�+�Z�s?gDa�����y~�F}���OA���� ~�ԠǷ��J�ہ��]8��k�������u�����+�1�Y��d�����'N�]�]�7։��!������G&L.��!ЬA�b7�s�^/�x��Q�,��"�pߛ8C,�e3����>��kf��FcT�ݾQ��Zz3j��b�z��jv�J�z�)��W%P/Z�*i�iq�
N I�C��k�����7
BS�R	Pc�j�ׅ��""��8e-0�� ���)� ���)�u��eHr�g	ԣ��z{>s��t��\���H�	O`��xbe[֘��x�k��N�x����*v-뽠��n$B4�=�[|��va����y�S7b�V�&98b��%��ɏԻAU�k��m����<�p�A��}&�L�8�[ox�>'���T�]�����V���Mn;R��q�����`(!,է�B7��i�h6d.���/���ؙ\�������*k�0�߄�Q����_�
���)��Ho������Z1���Pp}8�W�ye��Oڄ�2�t�@�Bڧ�rYf�ծ��a�G��B?�8���ě�eL����?��F��#A=�m�	�B"���)�"��=�,B;NXd0���S�m�GO�K�����,o�`Z��s�w��8ԖG￨�y�5R�&Hx�-ۮH559���>����xJ��e�Uea��+�Yꢏ��-�q��������w���=�Y	L�,Њ�4�wG�n�Κ��\5KJJ�I�!d�3�� ��0�{����< %�UC��ȫj$]5�L4h��:K�'��sR!���\�@��ڙ �
�����'v�d���:ko��a5/ca����!I��X6d ��Ȟ)ɼˋ������
Y=�44����/�d��u=����v$����.�j%*�f��%��1g���Bt!��!�UOzw�Z�V^��y���'�v+-t�W�9�[�qԞ�H��~>Ϻ|��KAJ�${}K�cW$?
vt7��a��t<J◑�����Ҕ�2�=�����iҸ���~u����&8�*���yT���N�D*ډ��L���;�F��	|5}�c�!�b�8���&CL���	o�~Pc߯*��/��`�PGn@��I-�ɂr�m�]Qs3R/�n�� ��qM�k>��ء�e���%I/�L�O��iX_[�GkP������K3��Ł�Z7A'nW�Go�ɼq�ShvuԠ���Ҳ�>͏
��e������Sw��� ��|����C*l{�I�FvN[���h<�2'�Qn��-���u-P�c�����]=4�	��T�'<X�Q5a�R��D,@D��t������=_pI6�����l�"q�t�g.(Y������$e���x���p� Z�ftҲ�k{�g(��}��U��gzk֭.�kۢX�0�5}���bh-���݅�����jz�^��|/�vز�|�o���Ƒ������ PK   ���X������  ��  /   images/e758c5b4-10e9-4263-8b5b-5233ba63df2c.png�{�?�o�7RY��
��B��,3������=Y!dd��:B({��d�!;۱�v_�����p��y���xw�5^�9�s��TW�EDG���sKEY�9ε��	n�'��h�_���88ʦ���{D~��O}OmkO/3w+///^;g3W+^w��MI:fyY��)o��i5������d�����N��*�a�U7E�����؇�x$�Rtzܵ��l�)�c)���=�n{��E��N,�Q�r��M	ِǹ�S�=��nF|P�26��������8���{��bB"�{q=��#���~���e9��^H<Ձ���"qn{�����o%��魡\wq -։ov�P9���ߘ	Xz*�p�9��n,rcn_9�"�I��K���nɒG�m]���_P�2F+h�2L�������Tm|��u������Q�7�Gù�^���]�,sD D�S����L�Z)F�0d ��
yh�Q@Y퐛�\|�E��-�,���A��Ɍ��;�(|�/��}$�������"D]^��N���c%���?�V�7�+�V���fU|~��$k�/�o`c�ԭY�`�R�u�1���Ѵ�K~��c_���=`⻚�͌��l*+A�n���'BO�6�+m��;F���M匡s��~9�󭒼��6ꅛ�ˍ����C��lJ�	<p���� /pkK�M)�b�ד�V3���666^�a�B�(��B�KII�s%�-�mB;ݨ�C������*S�����O��*hM^��.ƹ��pb/��]DDٿ����Fk�7蒇.�$ח��0<�%H�yבJ<�	S7��pOe���G{ez���3���5n���@e�����'���V���p}���xU��ߖ���'PD��� nI6Y>��{v;�t	B\����R�Wk
y-���Z�C��NF$6k,>�B ���ة���ۈ��Ѝ��$g��8��s5��8��S�F!�פ�&��+'�@-w0`�C��9W�W^���-�8��<���2>�˒�P��%�f?�o����{j��_��U��-�ϷC�G`� �s�8�O;tBXp�x	�zb��8)�]\���RB #�jX(�1�6+��­!n�l=O���#�������%P4h����"(�׮>���EJ�W��{�.(ϋ����y��y"\6��<� )����������b����9�r�Lp�.n������4��|�D
�lO��8׸G��H����Y_��aO�~�%8�L�S��P�v�%\�cע̾��!]��oNf�E0!
8�U�e��6p&�?�	�X-x��>��c2�)C�_~����|�O}�~8��K��	O�~ɽ_�]E���Jf�*[��@�TN��7�V����˒�����$
˪=۬��g�,��K��{�22j��5�gwp�7�K��f����G���8�4�l�8Mh��4�z�]�[�&��T��C�I>9��t�ߪ(ˌ�:ѭiL�3Yp�F�n��]�VR*č�y�+��yQ�uY�k�iO;=��it��+�!��T��N�Z0�#NJ��>����<Q���^�~����y�BJ���lKc�Xʎ�,z^T�$L.S�R]�7m�ې����G���3����HOUԈ����#c��#��9�+��[M���������~=jڹ��V\vbe`��F���Y�|�KT&���;�X�W#t�s�v���bӋu��U����޺X�G�֐�؇����h;���i��q��B8��Hc�t*������zAu'��_�ޝ2X�#�c�`?�ԛ�kӗq"����W���Q0�9O��vy�d$�^��˘&  �՘&���"2#R�$s�<x�qu]9��t�d���Í���˽�إ���x{;�d�X
u�,���,?���&�q��4A��.�s�O�So(�a����*���3��2��v��|���3���]W\�]�m�F�ި�ݼq�%m�Օ�]o(j.�R�dV�{�&(ܓ OZI~#9J��������b�w_�Z
FZ
�>�a;�\��Ml�rc�?80��Na�&G5����<!k\s�@��m���Ro��ׯ�,i;�0u�yG�*	�vCl����B�@vL�i�Q��2����E����W��/F�a��"�kH�n���X�j7�]���Df�\v���>Q�r��wT��p�������XN?{b������bώ�<%�%}*(X֝����G�ӳ{�m/ɨ$�ٴdC/���	�j�������&cs������^L޳������2'�6'sI����൉2���?��ق��G���/�����n-��W^�d�8)g�]��9�,����U���FA�)��úR������ވvs՟��-����"�<�!�w��� 
��b�}��@�`�RH���w(v������p��9irH�%�`�K�H[��f�3�7ov�����z��+5�s�5�c������lS^w�W�&k�"A�K�71L���3H��գ*�Z�C&�[W�
���v�b@���n�%۩& t�-F�@��-��B��R����b^�3T�筭�Z�S! ������v�WS����(�g�6h+�oC�ɱY��;��t��0�����*a~Ǿ8��Z�"�dc@(ż�Vcb!�C��$45���cۭ �	K ْ�������"�[%<���,���Z�<n��C���q�i��7~r9e߫�+�!�d؈$�Frd���F���Y�ޒ������U� �Dا��J
�s9�l6_]��53C��b�ra0_-��wy�
i�g�|�W�RA��z~�z�;��OBIt}����b�.3Z��p��2��=_���-��W(��pwz	HR?I!2�\�j�������F����@Y(B���
���C�"ǌ�Z4��m>�i��G��汪[jß���3���)��.��������X������v�1Z�Y/�E	����D�-��z�#��]�hc�2���'m�j��Z�U�3��q�.��E��A���d+YnJ"Y-J�\-���|oT;t�D���h�(��v��n�ݞb�A�FZ�VV]yB�9��U\	�ھG���r/%$�\�wE�iε������k-�ZP������s_���ۑ5QJ��1��U��`��:�]�Ǆ����Ӽ|������ ^l[�����W��F��6�)�jqF���2�	GD���!
��4&��i�V���5���&������9Y���_�U�SM��O�m�⤈�'nz����ۮ�&�l0���3jw6�hʋ�+1 a1����vb\"�ix���r��:	ybs��UE.�ž���Q�3����jw�~�r�|	�xM�	`Gq������n6�N�S�S�d�!�"%,��QsF �z�;��	� F������6�2�հM��)<j�/YO����"���rK�^0��+���un�_]��t� w�Ŷ6(�I�F�e'Xvާ���cz�0�DU|���SЙ�9����e����D:LMM����O��q����"*C���\Y�FߐI_<�8y������Z���h�[3"�@��xe�su�}�d+���}�S��R�-����p&�ٳ����;�ϩ�?k.B���:ڤ�F!k��Z���sJOk���2� �"���L�I��,(�BgP�:<�ٿ�	3ш���<7d�ϳ�"
ykK���`�s��^j�V>�U�=A'��CDXt.��֛.�P*@"�	�J=`�ce�{(���rc(D�`.��x�
'�l*��..d��%!��X�.Le�6|9"ԛ:��i.�FAa�6�O�Ҽ��/:'�p�=�B���䜫~L缩�v��G��b�3R�N��j��g<�D,�ꬔD'�|���e6 �,=��x��9~K��l*ar4�[�R�N����
�����V�j���b�ho  ��f�#7b�%'�n��[Sb��Cwz��h����1Y�]�D��x����<4�1�ҙ��`�2[����b��5�ib ~�����o�]i�n
Yx�7ކ�ń���]h8�K/�L9ءD����hH�,Ԁҳ@��yL{p�56٧�Dgי����iy\'���<W$�.��7G�1o���a�N7 �x㇌��=���4p�Pٿ�bn�n�H�/+^��t�hH~�>]���pՓ�m�:�绽h�鸹9�w12��CO��iNL�S�R8�v=O,��6�&��V��_�>ϡ�r�a���^�)��L�*����5��j�2B+��'�9A&��A��w��(���.�X�.����$��G0��:���w�O�/ϒ�.Ҵ�� rF�U�-� Dx���ŋ`��:�a��nK~Q�Uv�ƶNE|.Չ�4���`p��h��Uv�'��Ug>0�
=ڜ�X�2�s}��վ��S�m��l��?�� �*��U���䥭m���B�d+3o�#�kQ��o��~4^,l�B�X�D�����h�&*�|3� 
	���*h��%�����J�Ak)h���?-�|P�LŸc*�aG��G���#@�#��W��*�?��RȰ����kjÌn��R�xe�n��ٕ(��`�l��}�J�e���=837\����4��p�$�	>�D��
莞�g!��D�>D�����	��Ӽ5S=pP?*x����Ȟ��;�`��V�jJ�U��45I�ܺg@��R�'Z�x�24�������"��aӦ���� H?yq�u�V(�R�{D�TsЖ���*��韈V�b94��.Җ,VO����TIX�$�m��&���:P�p��G.���>�bjÛ�� N��IOYH��F�t���k����+~o����<15��jo-l��V �FU9�.��ǭ�2���7�&�m�+�[ĂB�����r�4�R)�w�qPW����Jj�_���u����m ���{�U��ݘ�0��j1+F�/L�́�3���u��7[U�ɚ�f`cd�:S.��P�Z��c��#E��1UUUH�_��03�x�~@_y0ך�� m�I�L@�"������|��Hx?
���A�,Cgkw"�����k�*�e�ш��1�/��nS@�qA܄��mEU���i�b���%��#9��^7O�=G�49�����N()�	�}� dKT �U!�Tn�4�yzƤI�ۚ�'�HOKs6i������Bd���y+٪�2-��o��^���.Ƽ���G�FyO^c�4aT����B5y��TNo���g�<���5�5��e�.P�q'tH�z,�~�q �bPT��'�l�NY ���6B<�{y]5!�W#e6@'�z��5� �Tھ����.D9O�¨�]�Z����˩/����.��r��W�W���O�IY�uxn Mb����>2�Tࠎ���̮���@Y���D��Іv`C�;���4�x�ji� �Q:; ��O˂f%�2�3��޾��m�?�ܛ�"2ꇀ�P蛛dr�ߢ�����v]�{M�7�)�49�#_��߆db��NJ�����H,���PfB�° n$��?�J�쯋��ٙ��]���ۀz��ߪ������ܜqc`�	d �r��z �$ZFF�r�}+i�d���9zt�����Ȉ>,�6����<��8�T�t�뜧2L�]c����������YQ�7n���@�4`W,0�2v��k��Xs� ���4z�5Y@�K�lݪ�����?��  -ҥtSP1r�I<V�U�
��"�X|��{��>��A�Z�T�m�z�DF�*é�p�����N��t=ޞ��Ҹܩ���L�I��vt�'����'zx��&�=�tD�鳻��Nt�4
jݗ9::�R�(�g��ҳ��l�����������>��*��M��[�/tA�mo󓠶��l�N�$�������סƢS2 �ڴ� �+�C�����T�ձ�Thm���
 8�/�wR�]�~����5��(|���Q���p7-�d�P3y�a���6��i�Ej���Yeii��8h�j��?�YB���q<Ѥ��lˇ����Զ9�a0��Y����x�'Q����� j���� h�M��c��>�.�˺���hp`�ɾVo0ɱ"n`#'���v���L_����}]�2 I�2A���Za����nb3��E���#hݛf7���d�ns�	-b�d�!�Gt1������'��_b��[\\�-��p�5��)V�C���O樧��I�6zl�/ei��W���]���e��Ls�Ľ�k�vy	����<0�ft�@D�,�����@�� @���(*aܷН(���q;M���D5�z�Ks�v� �R_f4���&7�ȿ�^�f���8=�BB=�G ���&��Y%�n�-U����4FWSG�WD�vW`��>n�Y_����-��7�p����'���'	�lK��qKK�3�UN�g�����-m'`��GS���\�A���[��	������ #3-_��@w�g*
�N��R
`�T�Φ�������<aǡ�*��\L��̱�i�{"�7"��kqR=�3�U*��F��/>�� `�X�ҳ��y��5ϋ����ŕ$'Dw�-�d��f �_t��D�Kߏ�Ԣp���!6|��
��u���g��4�������κH��2@�M`sB�������9��hS2�-HL`���3�<?ib�qe�	:�p�/��t��GU�0��>	I�w^34�v��|#���u[�����F!����ы*��V&�hF��OB�H�d�����Z$�齈�j���ŊN�<����)H\"-��>IRY��:ފq�_�2��^�aeu
0[��=_].�rGU�𿻷�G�	��9A����;��k:3K �7IZr��רվ��޳��4�4�W�ì�N?�Ko���+�U\]^�.0�6#O�t��NWr�r4m�h�l� �-��&X�gŌ���,ݒ���10������m�~��WL�XP�ښ�1�]���1�4VI�����.��S|�ɒ�<��Ė�:�QG�-�b��������_ŬE0�Jx񲫦�Nd`��%��=��ܲ�bF�ީz/ uSN
�R�#srXDc�G%A͊R=:�';������h�v2�w�K_y�T@�T*i���3�O)~�?"��ٳY����t)��Y�������'���c�6dX������.�*���q0�A�/�� ��q+l�?S�9�L�J��KQD2g���X�^��$����9NT��x|��Ƃ�����nւ(�t�����&h��^�^N��Ο�@���H�)�G�k]À�)��pWw�"8��(T�V i�c��t	���ٗ)�cR�8EON�+.k���I�J�]��X|�U����rF!聩� ��꯶���H�pa__�̈І�O2�]���uvN���W?\`�J��c4�!�va��`�X;��Ecy��U0�%������׿Ňb��;Xɂ�_,x ����K����}u�4�$W�����i(�Y����ȫ���y*O@�U_���03��{l��n�{[kt��uuuM��5����������<Lx���^Ui�V�^�NL���7;�~+����j�����١�㪯vUxqjZK���?w���@���d:e�e2��Q���s	c�Ժ�����}t`�%�	�]���..�C��xwN�4�
��Z��Zo�Ue�+�B�>��`{���L�B��c1��*J��y_	^Z[{��������tv'ی��F<$S�gגǤa,��M����8���L@e�:�;�����֧��y�Kt�ޜ(LҤ��,���_x;�U�S?GT�~��v=�K�hqsu%�j:���QH����q2z��L��s�D�Hʔֈ5#==��E�e`����@�U Nl#�Q�{����q�m!ox�����ө���;��)�Fr���W��B�qR�c|���7�����Vnlj��@>R��,�P=��,��"��҂S�4�� %d��m�;:�1�)�*0C�����dq�B�34���D�H�؉ر�T�K�fK����/!�DG�k��XH�Q��K��xY�A���E��4���GRc���,u���p���e֕�q�$x���9*rM���a�"ϣ�a�SRQ|��� ��w%^}���ɖ���X}r?��a��1�,`����d�d	��C�''=T�T�2�"R`*�C��t�ê�
�����f&��6*�l�0=�v߻�9��������H��ݭ@�W`*���`觭}��9WZ f�0��v<J�y`n��3�~��f�疔�Df��vH�B`�Ą�"�,B�u8�*
,Ŝ��t�''S�C!2(����tC�	_��9P	���Ҋ
:Y���ʰ�p�#�y�.QG)d��(CZ��o@����7�Mq	��/v�b��pQ���y�YF�jy v�-n����A�S�4Y >{K;RI�<=��μ��a#q^����qf�0�RH��w�j!}��;!��zߩ�9�C="���s�l�|k�l6�k������[ɸ�;�$v�HVߏJo7�VV��:�F�0�
ĭ�ڰ���&;�9.2c <��w�m͘��i )~�1�c��,,��M��1��g���pc+��B��
A���59�숛$�}������,�x���̣�����פ�)3��#�=4�p�>�Ӡ��CI����7���XY��u��"ʁ(.����Km8�㭒009I����.j�X����%���{_ ��]t[�n��o���4bbE�>��i�`����d�P�;�Ա����R�6�'nB����#(K��w�د�N1��-6��͡>��Y���j��`gD��ɇ�W� $��Ո=�D�MM]( ��XWZ��:��c�vQ�z�����i2�3Z.���j{!�UNz�_��7뷒�,n`4UΕ���ΊA.�N@�\W���Ր�(.(X�t��i"K�HA˒[x������,�~������N`�N���%^��C�m�ni�P����3�>I�U~~���\[��}��ԯu�[ϸ����*���j��!����� _�r�[��è䢇�<%�e�Y%�����K��*�)*���ׅ�����R1#B����j�_<�)�6���=	))B����%^�,�M�`�� DQ
��>���g"���v��n�@r���vs/`��+��!�3��`����f"�S�U����;�|@E������N�况���Lc?==u�:s� ��f�L�Sy�)�\mޘx��[8<f�#�>P���Q�BM�<�U��>��˝&�*�P�\����e�J�h�>�K��n���O�-�(�����{'���ۂY�bIO(xL��_�I�(Oi%؄��`���}�����0q��B�kȃ��՚������Q)2�5�M<4�,�yo��͸S�f?�:8,Bt�(s�]D	�]w"GnQQ��L�	0DI�z�������L2�:�	~Nm2���u[��]#�t��<��8�;_-�Ckk+*�.�H0�33C��='''���^y{Ӻ4���#t{Ł=P�e��=`T1Q�!�v���-3��P�^
IƳf�5ilV��0�'i+T�|@�W�x�����;2���|��v_�&���ܪ��b\��@�<y�$��>5w��#���h�'&��%�L�H�^鮞�E�f�S�����d���/%�5�.*xK��V3�K�͌���=��M�p�m��p����3�]O�bE�RN�%, �n��	Uj\,�[��,Uc�F�~}|�=�L�mqOE�А��A����Ζ���x桿�P/!�����LWD�@b9��^�Ewĥ3�Y�bN�P��j4k%��`����;ڄ(a�>��|'䊝�%��Ũ�q�_�P\����WF�fhYb�#�x4o����q�@w=����H���V�b|[W`�	l����V�@X��eId��͟�p��G��1�l�h	-�H�d^㵢��|;o 0�*h�AN�]��f�^��̋Я��8 n��3���nP�t��pZ�
�ѝ���-))��f��*-L��J�~	윴�|�<��.�?O�p�>�������W��"��æ眔�Le2)��w�'�y����!W]À
8f�:� �|�-c4���
i_5|�/b6ز���؃	o+%�ˆ�ً�F`�0��j���0�O<<*�4�@�I��@�K�i�'5 �| ����kpxx/���yѬͿ�ϋ>̘i���ׯr�XP���*��~�Z�����^����l�O��^{��{_l�=�e��I��B����c����d�%��w�O@��q��ð����K�q�b,A�-�,�sF�"8�J l'��A�ob��%QC�����;�� ��b�����5��/ָ�$=�t���P&���ŰP9p'd�'ic<s��P}�b��{G�]�ޗ)�U�.7�%;�g����}�����˥7�8dHn�j�'Ѱx��>��g���I6�@�D}�E/��qB�>-�`�� y���?u��|X��Jx,� A�ۊ"��5[�a�������*i��{[��Kz���h�r��P��!EP��=�.K�����G�[j�Ϲ���YK�o������������Ma1�09��}�4�GB��<g[�H+i �9U_�5M��l����9
qh�F�8�;��&K}�/��p�5;l.��w��8����P�t�� O4�dBg���p)B{|hUH�#	O��̹t��uٱ/��;6Utd�]�	�l��C�={�$s���J��>��ٕ�\i%c!5��9Vu�1, �a\;��F�{�C�����ʵgDй^���GF�{QoM�r����1�����E���z[�h���y�~�E�۷=S�:���HzG(�c��	5�{��
�������wT 2:bް��+ܲߜ�Mu3�F�����h�=��2��d)�&c�(0�]�s��3L�b]�&��r��]%�q[����-���6��?:��i�5]PV=k�=g݉��
  ��pN�d+,w��v��T;g�QB��@�����񦜽Fg7�����P�"w���}Ĺ@=;3H��	.D�Z��,��$}w��.Y�P�ZH��y���/��;�n��-��N�"����D��܁���{}Fg]�p���Ғ���||"V���W�2o��@=�����ZD�V�~�K�F�*�����8� ��u�����U�����@i%7'v.��A<��V�튪o���n�� gZ�2�4X��H��;L@�M+����F{��T��xK�k�F:7��e�y��y=+H��ZP���;*�����rY�J��˞�@�����z=��hrZ*�ب�X��"�OLNVVVj� O���X㕏�R�kQ������:A;�=ޙǕ��a�c�Y'I��
��N���@F�y�y������c� �2���Dn��z6}n��7�,:�b��a]G>��:�gUZ��#�i4�]>Y	��1P��_�6�'F<oo�@j���O9�3�(~�H��k�C��?C���pӥ�]=CT഑��۶YJ�hc��ۻ����M7�$xK39�-�-�UWZ���OK�69⊍�٥y/&�}u_�Y�I�~����^P+�;��)w�	~��7.���d*���~���X1�IU���c|@Id�-(�@�[[�q�w���i����2���眬0�q�۾��1�[��К巧��R��cR����������ang�i���]�Ǧ4�������QX] QU<rVߟ-�� �`��'� �N'�����&�w����כ��|�Da[>'>�l����_�ԛ�)���<Ժ���z��׋����Ӏ0.�$��Hß�05�}˞�z ��7t�"����:�\�g�59CA����6�����������`X�E�Ӯ�� �"���pC嗁���=I\3�y�%�E989i�~Y�=�z3Ers{5Vi������ycJ�]� 86�{g.�G�1e�rE%C!�F���3���T�F/�Rj�䎻����^�E���Q�g���*'oq9������́�8r���s��ZV��2��eT@�&z��g�r�K��t뽶��pg���;�PѼ�5_�N����E��y���㮊�T�e���ǽg�c���<���~YFڵ&��Z�-W�~���ի�Ai��9�{B��{�ݼ|�(NS�e���g�]m�2v�n��5=j�D+l�8`�����}�_7_ʒf��E(]���3}�}���b��)i��Т���^�kz�������y�L^a��)h|�2�2�*�r|�:���DM��������cJ���ƾ��&���چ߁�r�v�Y�9�s�E��q~7�d�?����0{�v=ٽ�	��r[k��_oF3(wG��+eo��Y (���)�k���E+��'8�����L���}}}.'�L~&'P�5(�w3G�"�D@H�ޥ�TI���&�"BȌ(/���]z�z���4_�|j���{���r�u�M}�u�1����{ȝ�C[��ސ�F�;ƃ[Jb�A{���#p��k���"�z��Q�����N�r^��oa�og���vc(X0�%�^�2ꇲB&'Sk�����Ja�?��y<�QV�\�'�"�hb�_���g������;#���/KS]@p�\	�u��G��vK�3��h�߀�П��J~u2�Y-��E"�)`����]Q�@54\�lxxU(�Mk������:�n�"O����a���ߨ����|,���;\�0H9Y�5U�T;��Hl��.a�Dc�?T�EJ>�͹���;�|�*TIN+'''�3-��yJv�����FUi!@K�<�uJ9��%�r6��r!jĞX��s�ZaP�\D7U��w�����o��o�g�֟�}'����D �����-��^Ҍ����D�ro���K����y����Eʘa!'쉈�?ida(�]/��)$2��gL���*Ğ��.�d�%���?�se����[����a$��.�䖘��6�5շ��r:��]S[�J2>�l�L�Fs�?Sz���ʈ�x,$O�9�n��a�v�T__�u(Ɔxێ��uSJJ�����)�@귩�T�����YSjHCxZ���/M6��W&�t�����? -F�^��k$�.÷�$ǿ;�D��_g�O�f5H�*s�H�&=��^�}Iۡ'}�ٟ{�$8�8�_���j��K�֡RT[9y�uYrI�K���p6�Pj��k��/�V�K]Ц����}0A�o"JGw�
_�>��_�D�C�Ϝ��#�̒�W�S��^uϿx�B��r�~���=�m�5]��ט-Y�0m��IE��OcӿV�\I!:=y�E�l�*Ŭ���^��	�}�E^�u��U>�U��]�������՝��Xu+<�ė��\�]l���1�|�	.�� b����>��H<Aɝ��@#s�tt���j5?�ֱ�=:)� ��e�m;��aS�"u�oyS��<zhA�m�����X@�k��6���E�?Y�as=w��[2ֵƗ�K+ R1w1C�j�?�kr:f�6I���z��iȐ�z�D�PO���e�ڴ���:^_??���.�;j�k�+@�{=*:����^���(��u0U�{9a�́�������=����.-�li�]Z�&O��"ޮ�mجqgP�ޛ��Q�+&h�NxxWn#а�$��l��3���e�_�}�����ã�ɦ�w�x��}��p[��v��� *��� �xڵI_������'����Yc� )+��P�ʓ2*ۂ	�S܄ݸqc��Y�"�����t&G�J�S��DDf*��KA��\�lQA��=��$���2����i)&7B�+����f��tع�"O@���0�'�W飺|;��(@�����ޤ�il*Y^gEȺ:P\f�O����$O#�kG�bs%�ԩ�����hI����Vr���!�<%F�{ �AĆy��jXZ�<�ƣݯ��p}���2j�8��y��M�X}��U�:L?ɼ_ö�33Ȉ��W�]�L%O�B=�J����\=.��_JbF����3�A�?�f��1�(��+��C�;�_�<f��W��:tg���5�=P��y�]KWׁ�KAB��ە݄n6��P+�{1�<܂���.8��삈�T�
�ɚ2a��?=c�zdID�+�(�M��|h�x�Xp��C;A4f��Q��V���丮�Cԭq����X�����W��%�B���߽%��p��~+�U���a�����W��kQ�D��&/�%PD��;��?�����67��9�0�T�������*�@������mW5��vET�&���ͮa��8���$�ŭ�(���Z�#�D�4�&xOH%("�79�.��+v�wS�:�ڶL�Ԕ)��&E���r��5Q$��������`lW��@�����%��t{��VN4m��Ѯ'��R1Γ���;����w?�>��I}��Щ;ò���*� �<�� ��������˝��]&������H�ѝ��R�5�������N/���ߟb4f���M�H=�i2�o��Z����g��*m*)_R*j��C�?�i< ��J����0�FY��/�qJ�ﯼԆ{z���
�g�ɖ�ll���	�k:���
V��"/`���d�1�d��9�_�͌���V�a��%U�"ه������Ζ ��3SSI�,�����O�O�/;����������2�	�t'��~g���+Qk��	=򏏂U�����L�3ԥ
������|���3�y7ާ�A�}�`��G���u�o�ñ"~H��#�)�X]���y�N�ڰ?drM�� t0on}��a]iu�8/%���,�]��I���/<v�g�27��&�_�M���9ܼT�x��������NMW�ߺ����_���0�?��ի���#jM[y�8��Hޜ���|��Y�/�Wl�{�]Ҭ��YG�?�2��dj�8|�������c'o�(q�(����#ƖQ7DȠ��,��@݇�c�L��H���
`�<	��w���&nG�˱\�j����/�r�| �7T���7ǘ:r�c��_�ӓ���v	���Kٟل�,I�WJp,���a#�h�"�q��2:�4<^��i�]�Xֵ�K���VyE��Tr�1��H�o��דM5��ϧT1�������g���uW���`i�qч���<�%�F&݌[���ۧ�h�'	H�@�_ٌ!ԚBX˘��Z�`|�B�e7��VH��?�0�R�-�Z�g��|���=�������@G������`|O�r���B���/��Ŝ0���н����X�X�_�����@�<��e���C�Ԣ���/xI������!L��|�+V�ieD_����IHo���3tv|�d�9C���Z-y{B�O0i�y��+w��+MiVТd_ѡ},�����D�8��Q��&�ӓ��K��s�6�v[�q��Nq��E�����A����vb��2}O���*w*����weǼ�����67�81��f�.c����Wf5������b�-n�u}7;8�<�rG�E��u,#S��ٯ4:��@���a��Q�8�=��5����S���,:jl*r��|>���rR���T���"�@���G"y�ÍD�����N�?����+�Ա"Z��!ޑ�YK���"�F�Nu히�Tӯq%LKvȾ��iQ
X���:*�7+�H���Ew޴F~/�ы�!?�f�r���{������7���3�Qq}]]�7空��tZ���{���j�&fx����u��/��b��R��!�BBB�gU*L������J;t uImj�F� ��J3�׍�$�z�Um���ӻG�T|�t�EgdD�uڥ��V#F�� �QT�H�e8�\�<H$����	�-T8'�������*	YX��9�1��V��c�*I}0���"��R1((p(����������Z�k��;����p=K�6yN�;h�Ƶu��]�=���J[����k	 �����wB�^t����u����U,RȄ1��z&rP9g�9�55���\���!#�kMOX�X���a������g"?�ll|��%5J�T����ˌ�r4]S-KܣW�5v*�A��l�3Tŧ��v����{�O;&liж�^2����0���r��\cP���!HH��"���\]���>4�"G?��s�Fn��`�m���"{�o]����A������):�v�E5G���/��\�ȇ���������|�)j3�D/k��I�|��p�n�[s�
�y�c>�I���֗�)^��g8P� *�p�oܾ��Q�i�� �� �Ϟ,��EYj�	��=�O��y��B/��ʻ�}׾���m�܁U81d��ɨ��[�z�@�0?Dc3�4���0�㓽�Rʢ�a��7<�'��+A�v�n{��b����}��[K�2>�"ޥ�ѭ��j��%_ڝ&��?��;�-��qi[���V�JmiyOس���6�u:>���������-���t�he]�U7���Y����N&7g�S���l��:��崏�Zś�u?�U=;��@˔����
�2^��I�K�j����ae<�sX�l���AH�M��#��QjE��$��� �����~�H���n��'��#R�o��^Rj�ge+=��I�����{�z��޴Hk���$ü��6WS����)?o*���VZ@�ʍ��x��m/-6o���(Ϥ[0�Hˏ�+X����n�]�I�i�g5ߓ�>�2��F��f����?ԝ8:hH�&��1�9l�W�X_\�S�u�?�S��jl�^�і��\W1���E��n?�^Q(C��u����L���d����d[F�2��\�w����e�qM�t�v��8m�+�g�/�8Ԫ!Z둎�G+�DD8��5��y|0�νD=����K~��O��#�=̠�^k�)������><���i�n6�O}c��<ű�(˾�d&�*�1�wg�/�<�F=�S?#��Z�|ez�̆@t����ח)�Z���KCr�� ��3��E�'���������O.֗���JH��uJ��^�L�O�X	�(H2z�v�{�e��Q{29(���gA����Ƀd+�>#..�1�X���kL�����P��4H� ��0��aQn���ҍ"�4"H� %� J��tw)��tw� !-�H� �)C���<���r��9��{�Z�س�m�"���_:43n�j>�Ѽ�	I���3�J��Ʈ�;!CY�o��<���e��U� �(<C�� ?�
A�,:V���<��b6�Z��St����gm	WO����}�t9�4,����X~E��GZ�1�p�4��墙?����O�Y�}�_���3ͣ�TE����ÒED⌱�'�B`ƹ|iXA��[3��=��\� ��I�?���T�\�4%�B�ҘG�A��D��Ʌ�u�\��"�	��)#q�_Z����:]vt٬�������˒�}o�I��qۄ)��4�>�,��F���Ԏ[J6X���@d�s�+�ծ%��0$�	Шkn�`)�0ţ{������t/~��H�y5�L��2)%�|�P�J�e���A��uϓ��Id�����a�<6I�?��/H8+�=�ۍ0»�N$Q^̤ׇ@��<ߴ�4��o��w����Z=<��e$�OG&�(���jSt�;V��C��_��p.K:t����Ȟ�_A����*)f�\��*�S_�Ϗ1z�ΦԔ$%���վ�fO��Orɿ �Bo�V���l�V0���&p�MO��o#�y~V^xh8�Vu�]����V���W�+G�ۨ�7�l����+����Wl�X�E>��5�5����ˑV�T��/�g-���ի���.r�T,f�Z��lW��_pK� 	򳧔ύ鲩f��r�~�)�IѼk%k���ȁE:X�� �d9��=��N
V]�3�~{1���9���N ���V4�7p���丗�n�Ub��9�ٚ��Qr���_���sΘ��i(�d�r��?�8�z7ܘ+q����/߂B>�z����%�d_�DK���Ro��؞��ѝ-F�i?��{��3���V����I����Y9no��byp�A���s$,�y�tȘ�*��8�����M>^��A!�u���g��)��d�x'�Lg��H_�z�^�h�ߔ���#��f�r̒�)����(7��ŝ�Ni��r'��j��۾��Q��gݡ�1l�醗�w�:���ѷ3(���=��%���[���H����Q~�i���>'d���ab[2&!dw�[D�0os�$'�K���`ц�_�>ÜN�e]�_v.(0D��?^OT�����|u�'�@o�6y5��J+y�>�iw�f���G��E�����5�0�\�
7S�@_��O�vZ��&\7�b�ݜ����L��b�[�i�3�u�Y-xV��ߊUua�@�¥�0��w/��1�	�\f�ݭ����݆W	8t�/�}+�o�%1}rq�L6#((P�:��F��I�$-��8���q�O�Ӷ�H��%�m���#J�2L��%TUc�dfm��:��Yx|_���2�;h�2F�C��bcNOO��*�
0�8ѳ8Y;4[&�!��of�!I�ML!�e?�n���#��.��G~���M���`���_sM�s�'.��d�x�� D��n��w�N+ t��.��hY�)��M��L6y�=�&��օ?�K�+'
 ���f���`��JTʿ��X���=�!���IG<�I���Q�߀���MֹHr9<���-\竇�l�(���0����أŪ�u��7�����#�ZCK�JT�'&cC�{����oR�ѵUk���P���;)�HQ��:ʂD..�w&�=+�a]Xt篤����d�92�F
8H�m�����_���c��Q����	��g��P=�!Ò��%�G�V�hh��}?������6��/&n�jNI[���"ə�Tp����c�Wb��߭5gBU222`]#�s�Z�]�Ex�<�]�7���PJ
��.��)1�)��ۻ;����"�~��B��\T�S�BR��p��ֺ�'ى���
0O���#2?v������]ݝ�۠�[�P��� �b�xV}��Y���㔚�{��k�����h2AZ��tX'`�FVE�AWz�F�GjM�C �<� �X�c�Wzǽ���8��6|�%��M�Y�7�4�JY��e����j(��a�b���F'E���C�Z���?��E@)��bW��ɽ*C��d��w5���I��=Sc��ii����!XT���4�`�����r��'��*��=O��7�E/�^?a�kN��~�5���h4~��̈+�-U��:��rw�4��`N���a�-���qs��YpJ�˷�hTm��~L�׫J��)��C�54�>d�ښQ�#���p�-��qDh�v`��4�|��Zx�_�o�<(ǆ�8
3l���xS�O��)i����딗�(W�O�Z*ب��#�d����Sb�������859�T�KyX>�Q�hX���͖2��cd��=�����5��6��Sl�'A��XE<I�	jK�����|@����I�DМ��t��IJ�2�Ԉ�c��R��)q��p�������ok����E,���̱�M�?.}��k��^�bRܦ�5���>��
�^,***|��a��A~�Xt�d�R#^?�]f�$dD����O�=�pS�.�f���J�WܑI)��f�~��?�v]�����owJ�c�g�_�f���-J�D5�t��>M��F��?�NN�?Pt�B�o�R��c!|�pNBB�RK�Q�߈K�I��,3�a�4���Ԯ:JKU�?3�."�fh��twg�0MG����X
m&m4r�f���v���Ѷ��^k�|-�s.�S�y5	�7R�%����[*|��@D~|�jkޚ2 ��gR1�@���^�@H2�C+C�]�� ]TQ?�[�m�8�[2�{�`���V:�]�B�|#f����޷�F���5�5�k[��LB�J�\1aWy�<�?��-H����x��MS\D�2?Ճb��?����8����</�}ʻ�jʂ3z��G]�O���.����M*��i?����pX�hP_���_YQ����:LAa�-n"��Zu"N��{���H�
�gtm �z��gg/���V��yj2Y�[�;��~�GGG�h�\%�G�.;���e�����1�\�Cw���K��MT�܊x�x��$�����+J������.�I�h�����?Oڋ���Nn�'XX.��[>��n =ƽ�o,y...��~��6t:�;<���2�Č�����	��f�ԭr�"61<q�O�X~u<�����@Y@Z+L!�{��guNBr�fW�q��꠻l�ѳ0��8��U~El�j�v����3�������W���?�H��E�p-ޭ��N� T�-P�8f�}u#]k�f1��b��9~���ݣޙ��V ���e��]6r������Ֆ��tD��+��)%�i��r*p)))j��������u䫟�|��lG��_AJ���1�J�fߔ{Z�~�R��o�f��X٭�4���F�f��u�JR�j�%��l�o:\��x�4�F<�9﫶��� ��K�s-aF;�^��S��d��օI���T��U��I��'�O\�t��)���:����'O�P.���ٯC#e�B��?���D���YJ?����*�ݾ�$>�vD��2�)��覷�M:}ȩ�o�v7W��˟>}�]7����S��o�^����i��w��U����ha�F[�@��5c�FoG�X쓽��F;��<t�ql�Y|Y���� �f�t�7�͒�}0�~ej�}��>)k���ɟ����	$�����_���DːF�o06�7�M���J�.�`��V��[[�Yt(�#�oҬ|iF&i�1�P����S7լͶtP[\ľ+�h7�����;��t~���\���6}͎_:[*[qW��^�����$����� ��i�h���;C)oo�!]j#eڄ,=�z��,�sU�hb��~���,l�Nrp��`|���*&����uKtf�$<:���U����ـgҢ�9G���8�xy��oX�s���(Ή���6V8��S�M��W�~�5]�$�b���� ��N�a�~^;��Nb�?~�#�%����#FS/���m�,�N��$t�0�`��8PFo7m���d%v��ڎ/���7GC_�E��x��ת�I���S8��Fx�.���9�E����u+o�`YENJ	����	���l�+pl:���t��ӵ���
n�ֿ�M6�zo����!*,��������+uu
��.+�fk���!</���G�W�����Q�ј?1U��,�!4��m8�<��W7�s(t�o�Q��qs�E�
����ˮ��k�K`w�b ���j�UA�9�f��|���Ã|����M������ed��MQw[�n�Ҡ㍰Ԯl=��Бy�����9VMYX|���^
�$�d�����k2H�+M�������nC�i���1�P"�/b	k�#�~}�|+  W����M ?Ǻ�SC�̒�m�����RR"�?��0��8���\�æR#�"H���J��J�۶��3���B)�s��>�d�jL�3q5xx�lP�a@�4fz����h{�*c�e�*NM�;�� �.S�>��#a��-0�Y�lf�*����*#3���xޛ%�
[�Q�\���@{���Qd=�X	����Vj�����E���vs~��������m�Q�O"{D���_Q�0�SK�(���
ķ�����uv��H,���d����UY��B./���kf�bC�'f���aK
����P�V��p�N�͊A�!��x	3AN5����2-��¶�B�:-v�ܫ'���� E�[n�*z{�C�$�a���W�`��N;S��񼰤�E����zؒI��A�^8ml@��e�f���ܓ�����À�gg-**z����2z@�SN��kEnd/MD������@z��u��G1���nls!����\Q�>|5��}\j���
�mR�Y���2���D��%M�>K��g�c¼N9�H�W�C�_t���Րhk>&L(Jbi��(zs�\�BJ<RU�����w�n�V�S	��ɷoC�m���a���R��ׯ_#�J�#O�/[9��'Ŷ6�]C:G�f�t��M�_^�w���j48Y�r_⢣���scج��%��'�=~ƀ��&kqo��9��#��.ܾ �X<�P<�:QlLS���z�P���"����SS��4�7�4�|s��4� ώ�qo..���9Wq��ںY�7�]z��C�/��4�ٔ������S*z�|Y����g�p�b�
lO����o`gggp�����DLN���f\��<�D^�=�0#u�g�J
J���zG��/x$gj�L���ϑ�V�}s�H�O0�]�_�lLAm�й��>�\�z_�f�����6K2��)�U]e��b[aaa�p�~O�*��c�;ޮ��#U1��X�_Do�VQE������������%��X���e�1��������Zy����{dTT�"f�^K6:�4u�x<��>4���{���N]}�HEw�Qz]�$���{���""!�<� ��`�,�}I,�I�~T�5xP�"$�H��L�U�j\0�gv}���-Ϻcm7��|�~��ao�	4Q�@�}g]���p)m$/��D��bE�{} y�S�t��Ī,֢K&C����R0���)t"!Cy��c�w뚍�\��#t���G`#kf��;փ�b��H���"o�]��[��pY>�Z����*gC͖v����2--~�O�ڶƋɤV�BB������c���`$�.#'J�@�����1�pcC�S��	��3��p������@'@R��m��O������x�?'��\]��J�ĢBLQk���暧�*��G��\]���,ٵ9�6/�V��]�*��	{Ӿ��Yk_,+�X* ��ON���>_0	��7RS;�< �B/q���YV���$b�wH�\<����j���� v.\���kx�V-��i�������̗�0�:W���N������4�^����� �� ���l���2tߊZ�**�������>�ɚH�<��S<�ac�n=�44�5�V�U�A�Z~�V�4r��Ql�� ��G���_���%!�]{�����[�̆����6/4�gB.��/X�O��[�v����0�|bK�f��?O��6�i�\�	���Eb��Y `��>T����PX;]������� �l`h���w F�z�2��˃�Z��
������װ&�僳���9�gZ�lx��Ci$T�-���</m�M��>{D6y�D��n��y֛�6Ǘ�����[�"��G�N��*%��\r����k9�:�;�PUQYxhe�s��������^Bb�>VV����o�<) L�9b�y{/�$ ��)�j�/�#��_��	"��!��p�3�&j 9\N���5�G�;����O�8wxBL]�6�]�s��96��Zfr��5:K�<m(���|�#z�H��7PUW_��.�8��)^���؀h!�M��$Vc���)DhP�r7���۩Z���	q?$0����H�^!���+��)H	�ľ��*�N~�Q��y���|�ڽ?��g�(7�M�O�BD�ܩ����:Ag7��>���R}��Ģ�(R����[R����Oy�Q��	�V=B��B����B�^� �7�w����MC����X�f��*2��jT�F�_"�8B��������:��*�sD��c�l�^��|�1�Đ_�$��	����H,�2�0�ʏ�_K8�ko.��U�V���N�i҄��l:L)�bҡL9gE̹�)?
��ϽfI�x=q��W���+�?��r˟,��YQ}��ݣ^=�Y�_�zh�1�M<�����g�o��(�s{�qދ�󍝈��-S�
5���Cm�? �h�,���px�X�r�EB�62%8 L��Z켫n'�����D�Cj#4���k�YK�I�������Di��֔�,����u��!2��9��|�� .��eU��%wPS����6�����Z� �Gn�O`~{�(B��j�ԕ�|��eQ�0T�󌙱��j��H^��[ĵ��ׁd^���T���5%���h.��ȭ��i���S���]��ZGW�	���i�'9r�A=b���/4_���~��䱒<�F8�l6��k�0�K<iN�0����қ������s1�U�[mƉ���A%�ϩq�Ǆ-Q�o��X�\5�JJ:�yg���t��7�9�">I��xp�V�D��m�jj�o���/�eD��U�o�	�ec��]����1#�൵�ꆕ�������P�A܄'q$�?�c��X��::8t\^\HYL�ى"�D���r�CY���9��xNO&t����Ӟb2�����%[���-`�^�]��tٝ�Es¦��֔.�z��o�]�	��z�A�,�d�Bv�~����Χ���������� ә����E��c����=�n<�:d������%V�s������pZ�p��uT.������W����^>����c��}X�d��j���/_`�㻃��u��.n�Nx��܁?��7��o:k��L<_��紼 �'z]YbŽ��Ӟ@�z�F
��g�-w@����w(X�Ű�$9_�!�cj|w2|"mN.�ϭ�b���L��}!����Hb����76�`)|�ь
m��C�e��>���!T�h�A�x(U��DxV��L��%��c�i}�L��}�`9��ȑ%�2����r����6�����j?,D�8�|��,l��켲2떊f�`b�	��9n�N@�f�jκ��dpB������/�&CYee{4���&�<��w��2�~�����_�5[�g{��s�/�0���T�M��o�b"�Ӽ|�UW�w�?I���8��?���	k�Ph}�Ȉb�R!�.-�J�fe�^�6�fO��gDs��o}�P�sT�۬�ݵ�Sy�L,�S�$h�;'�e��=��'�gckK\Aa��[������w�
C�(*b��� #�Ǥ�mb�z�	��b�l`|��|KI��yT��9�u�{������;S�e���r��������aR4�q��ך�v�,g�mc��.O�h��bΉ+�K	��z���-0|�O�����[�����[N#����"�����?�p�%'���%��YΚ����<�'ssE]�!�\�H9�T;Nxe%I=|�9�=$:�cZ)�ѧ$��-��F쬴���spr
��++)�`#?�b��}��^o=�{��7ׯU����v��L��}Ӂ*;;{L�C��	yhfV*�����W��<��4��x�J_KJ��×c�u��P�׀4Wr�����$TL�Ꮚ����fmb����������ry���H&�5���,		+*jjY���Q��/�%_&��S�|�k���y�f��*��+R}�4�L�uxjjK���t8'?��c�`>v����k��X��eks��
6���י���>ꋄ#|N�(��պ��@E*��������w��84R���6>>�?��
�F�$��P�3l�$���_>MȈF�w%~��~}0H�R��A;��n{K�r�V��Sb乊CJ"�Ŏe[-����u�:��+c~K���8�۫�4�{@��gO��V�%�7!2H
'fg�K�Z@�5�%L���ș���vS�@���/؀��s?��}�D��܁l!y�&/z����>fە�H��B]�q�8|�PEb�}�3q������3��X	H^��1ޕ��	Z(B�p�*�x��IJ��F}8�ʺG@��h�.���P�w��Ԋ�p�鎠MpӰ�͔�V��ѳ0y�+fz�斗��K�J ��������s���*R-f'!��2l�|�����xC��S(��ӮN��o���#��ȃӅ��[ ���6�Q9���*�怂3��� '��w�F�ss��1���ԙTj����MDc����54n��dT��P�T�O�&��������g/.���P$Rl@%=�!�1T:�P�Ȅ��Ssй�^�]QF����1�" 
@>*KH���I���l�Y6����9lW��E:���U��{���� ,S��gؽ'�W)ј��c�ұ=���NS4E����6�mB�+00QI<�y�-�d�_�r~���8'����φ��{`���iN���������[��J�U�[�׊�+]TT����EZJ�����Jo�3l�}Pb~A�Iº,�4P<���w���믰�_��.����iȬ��)�qF�	L���DCC�����
}>v�>倂�C[�M{+h
ظ�ۉ��p�ՓTغ���-�33)�Ap��Ƭ,���44����HɈ\$���	]1G��գ�	�j���=�|��At�ka�1,M��M������5(h#u���)�Xe�
lf���V��ӌ�g0$��Sv�2N���G�::9e54�O!E�E��	
�c�
3��wc7�a�A�cIn#:�6f"?ƭ�Bz�$�z���rc�]Ww$n��lS���f��QQ;O��GI@}�O��?ڔ^nl��A�d��]��QJLW[��A���ڬ�y�LJE��$^��g�8!��2,tTנ�}� ��[�
t�?օ5�HERe��9؋�2/t?����0�,ə�.�^��dX~�gY}�@�v�K�7d�e]]R%���2�p�Rѩ�#�|Sɍqv�Bg�X)�O~i�g& 0��-�h��X���v��OЅz3���*�Eq6�zn��!@�/LW�X�Jf���W�-��+���T��<[��'��joS
�(|�0�Wr�՞�N�@Vz`O5���rT��{���F���]�8��~�Wy��%���v��ʅgO�;	z�	Gda�:-0���Q��V�c�~}�z��?�;�0 ���݉m�����Ԉ;��d�� ���K�:��.��2�� 2^��ڀ����F�_�#R��Q�Q�7Kˍy�(@��{4���y��+?�k%ە��,�A lBכ��KDqaa+�؍3W
�݃�y����� YU{B��)'�Y��g�t�7h& %�j����g�a*��s?ݏFgi(��� ��r���yr+��QcE���|�4��RG0�k-m����Qn��`�@��MV_�Do�C���j��a:8p[#,����h�����B�n7��mWzg#�����:=����lW��}���i�>^\\l��?�Ϣ{�������e��+[:�s�=��&7�؛�ل���f�i:�2�	y� 02��8���_~��2����a�x d�k���M�H3� e�ܲ�y=3Z4ň�T�>BA���d���l��LMMEe�b��{�3���� H��)��(+էDmL��q'�������?iaK�*��w��Bdw��W�J��ű`=��RW������$����}�	0��N�3\ �\��x�(�t��J�p�L����S�C������ �
�k�eׄ�Y3f55�Uj�X�+#�9p�.V+mki�������ָG#��l9��B�^�͍5�z������
-��a�z~Y�O�9	 �� !bA����������:{��kr36�x��]Ⱥ���^|�Ղ,&�p�e�LK�a��lYL.��X~�\��A'6�Q��m�b�`A"yBq=�F�����$�J�ь�Iy����UUU�_L�콶��=aB=�g>'fcg'��D�W
�����j$A���X~�C�kF����>������ݷ��M�u���ȧ �P@�[T�&�w�  ���+@��]_b�G���kƹ;�7�
��T�$�j��g_����1zzz��*�n�yz�u���,0�!�:_�$�2�v�ܥ� ���\:�=��`
J1f���x���qƞ�r��C	�s�q���ۮ��D�o�����S�,��Z��caaa>�+>)i�#�~�,-�!��-�|P��sR���r�ѽr�nc����̻`��W�|_c�O:$q �v�&EyxJ�&C|}}���Ĵpj�xfp�3o���|LFX���fڐ���G�O��|}�g�=�=D8`݈Qo�ۿ�E�ӡG�C�*���և�==�}�-+).F^f4��߿�/�������0��~�x8��`��H������:4k�=�l*&B���i���O~c��>l�>�vN��7����l�����?|?��,�ZB�`�Oـ�q�:%�0 J�;����\�䱽,��������S��q���u����.[�S��Vc�5y)���D~ �Y�Y���~�ŋ�cE�q�{db"0-�ö5Q� ���7uu��p�� ���r��Ͱ�ÉA�M ��LT��3;a���%HP�/t/��7A<<<�^7dy|��
h�+mm��I���Z��-������[�'�&��k�M��G�gru2���
:�~upt܄5�omo�b����s�6P3Ӄ4g�:�%4�J�o����-i�ǵ���o�S��Y�ߔ�jj��&0QQ���7�TO�y�<!���z���h�H�ժ����hu��@��m��y&��EEȭOrv-��
N�d��,gFIEe��eUԽL�������R����v	]�0f�]P��W^δO8� 'o�A�ܩ(c����*�	�j�U������ٯ�\G�r��%����փ'�q����;$��FFm�ß6� ��F�a�F�N 7��:�wk��rd�P�B&(Ct��_
o����+���q�l��v�ԂN���"vkk+F}��0��(���������j˜13#�����m���3FZ�^`:�M�Y#L���A9%pO�J'����i¡sssQ3/_It>!���f�i�4�Q�k� Ѝ0@zIF�c!�D������ P���/(-UM+h��3#)���Qm	�A#�3�ܘ_�aT�CR����N�gXJ����Ȓ�LT�+ȁ����(C�<�����O)_����AY����_lG~���+q��!6)���s���P���<~Hk�K'����j�颦���|��yf 돸�B�X�����I�~�V3C	L�J}�o��c��]`
�io�u8��� �ǈk;Uk�h(X���=��J���@/��m}�F�	7�Y�e�FM3o��"7l6`UG���"�D��2 1 �`�x��?�����CF7��vrzڽW�
��d�Ё�.�5��ӕ��)�I��k�!��^jP�"K�8Kl[0	�BA�i��>�7��`9<1���Wp�i���;v�g�p
�*�hYB�[ ����b��,��K����� .b�uD�(�fza���hC	F�f�B�yU)�uW+�����ܣ��/��'ag�}�斆t����I|oh�ͻ�	��n�"Ѫ.7�$�{@��F��q���y��f��Ó�����j2�~��*��)���&4xL����T����
�����*�j�cj���]���-�'ʢ)�`�С�@3K��;N�~�Y��A�/�O�B�d%�����񊊋���C�0�ߕ;�R$ĐD��%�m���+��vQ\��0��_L�鹇��?���E��2�CA'x0P}�-����X!I��*]�u��;�"�-#%��jp�l!*Y.elLջ"��B	0���)x~��#"�V�e�p��6{Wa����=�� ����	�Śe�?Dz�W�V�o�@�A74�-6�t�;M�`@�O��%�D���s2�c�S���ah�$eц��ƔP'%-C�b��nw���9;�/�)H(sR^92��C�r�"��v�/�u�v֎�|��5��G^�$ � 0�	�,+,�61��NI������O���]�F��*-��Oa34�ж��'��|�U��{��E
~Al��t+���ʻ�!⮸?��$�i�F����A-�?[���Bn�KK-��o��'fXOU�� �C�t��
y1PdM���87��+�xPp�uizk����cYf�MMr�/�A��pbw�+m���֮����U%��H�8��<���ǁ�fY���y7����J}�n��������$}b� mX��n��2ӳ]�!��V�D���Xb6e]��|#9�K*�˸�ƪ�K2�
�H)�ĂPysyn���A�I�׷�՛�kļh� %G���&��SL?Bo�G�\�Uy�'�E-�<��{�ϟS�q_�ܧ$ǧ��Fl�Zu����$ﺭ*7sxY�E��S鎲���EV\AG��FaS�y�w�1�ǯ7��6�9�HOOM�(�Ȉ�_;~#ppp��Ͱ~o��Bh[�R�"�p��c_\Z�{��i�����?
�d�\7����A�:�����mT�������K��:{����=���-�>���;g1�4@�G��3�a9S�<[ ns�1���V������ߺ�]���ibē��2(Omp�)R��w8s�w�˘�b9}J�R��m���ۻv��&�uƹw�'����x������!�un�[	ɏ�����p�ٶ;c����M��s���Оm'Fd}��>?S`T�\�)#>ƙ��,�������*�,Ժ9ί��{s4*4A$^�Ò`a|.U1�ں	%Q�����iF����ž Nᆲ%_�[��=�n�!��K$444�ᅇ������~g|�mil@�|�m��$�2�l��1c?4��yh�u�0?-��υRn�[�{�2���~�̒�f���iFK� �'��nZ#��$��}�2z��w�'
�����������k��/�QY�_�FFFp ��Tmu|?�����r������j����, Q$��ߚ��1-�yOD�;��Uң��-+)�5|����H���Dr���q�aA��� kBd�
�l�lI�=L��i�t��K�/�Q���W�.��e���a-��u03�.	A��s?�4{�3Ʈ�p��yUbA'�ڡ�Hz�\,;ŏ��>�~�e�=ߍU���DLUS�b8B�)���S�������l�P�v��1�rݱ���+�7�0�ÿ�a�=?
̉t�>�ZK�|[����|�ٔ�R_���;�n��i`іt~���t���8��i��jMo���qJs(���o�՜����Z�U1�4K��Vv�R��}���Q����y'b=�8T*�M'B��(������<�,Hd:��M�R[�%Avo��xP��S�G?��u&�]��̣~�����t�z��㩐�
�HmZ���->vC�g�hE�Z	�݄���y���n���� �9�����S��ەu�ϖ#�p�����/!K:C�mSSSMp� [���(Ԙ���j6��w^lO��j.�J�g�An�_Y��{��|�_�i�C(�1�FM��]�1&GF�c�袸d|;��)0D'6�?����gIv؛�E� �0����{���놾� �_���C��6��V5�/����,2�}�vs޷�?Y� i���-٫�>>�]@�7o�_ERWV�#v�����|[��{�! 넅�O��?�Eka�G�*�k�9�Њ�/����R��Y�΅����J��hQ��M,k2�k�骋×?�NW{z?�O912bK��P�n#�aogBW
x^˞��:�_l���BnsU��U����0O���T�V$e� 2�_�O�+�ׅ�� J NV���l�e��ֻP���ɉq&3�s�s]/�o#P����ĉ��!m��=^��@ux�{iݰ�Rٖz���������,/:tn˭=���:$�G���c�%9!�U��NU�( n��s�zD~̢v��r�W��~=|���I�7�Ym�=��r��uA�ybי�����%1Q�AA`:���oT!,��T��Er�0N� ��?�-�-��߲��GVWW�B�o��Yj���k=[2��n8h�w��hPQ~lm���9��tB��8U��J��>�K�ݺ�4����?����_KoH��Q�q*�pdR������d���4��4�����-��ӧ�x;����<�x ��g����vvM��/^cy���׊0���+k\1�F�ūO$̫�d�yä<�yv�j��א)G�O��֝�&���\[<���_��>Da��w͘�iud�%�i.�{=�Z��m	�=IWK�O�WFf!N`9�}��GT���P|ZQ��d�O��#��,,,Me���ӵ��-��0�
�;2�ω�m ��a�v������@��z��x�$�R�W���sx��,�t��*�V���|��� �P/�]Y��y5	�R�JLG�oⲮ�Yu�q�ej�{�����5&�%Y���:l�#����*7��9�=dM-��E~X�)	1��k�[ny� 	9�|�j,.:�2�gF!/�>���u6�L�{���gM��n�i�Z���(t���ް+P$�O��z�؏��b0^uv]f�KgM��ˉY��N��ޯzv�+.�%˕���o�!��U9˒Ѕ��03�) O�0����*Ҡ!��X�*��ϼ�"M!kؿkn�%�=.����I��'P�(�|�����@e�>������p(�i<̫VdG���D��-�OX��}Wi�g�(�����H��q����)kR�3�(�c�(Ae����3n:	�+�;��S�:b���{����޻R=�r|�ժٽ#r ��U���\�R��{���)D��7��5���� �+ �{�8�[����}�R5�u�)\+휃���q�R����c�l�B��w�;�o��Չ�B���̚dr�����{�֔O�t2�Uf��Y�r�Ui�kQSoe�&]�Q��²�fE,N*�<�]��瓅�-��o�E�O#s]�	.�c�?�'*?�����p_8�rZ*s�wlm�Y�S�26�Dn7���n������q��@��Y�5?�Y*����n����h��5Z_�ʦR���x�}���0��t�WXk�"���_�`6�0��@������6vH��x�:
����WȞ�+��t/q%c�e��E���n�BG��(�ރ�o�[�dY#�*6�Gb(V���[�g�;�s$ԉVbW}^F����Xtj�����pI,u�����,���P� B�� �k��J�R��H#���bP��8��@�d��˞{�?�C���F�NoD/u{f�T9�eI�c_�:�������{<Rf̨v�]�X��	��_�w�+m*.-}V��cL���Й���)�����q�9��(|�ԅ���D2Z���:.��Y��I*]��˰�N6p9�Y�t`�P����W����o�5�N8E���¬+?�!y���+j#h�q���691ͪ!8߲��	��]sb��T��5�.E�ݑ���b�BӽJjz�w�(�I��}��GNP�!Y���*	��a��0H �|���ъa��`�l���?��J�y��mhk��'6k�o�k�����yW��� ���9|�j�C��d>gQ=ZWf��@�q�O�������'���#�1nQ��w��{�ݚ��|b�W�驽F7Z�W���o�!M�,��+ W}�]G��|�g�_^EI��Os���+[$V��N���b�y9�YS��]����m{�UdHwh��A{gu�.��\hf�C�,����}|�<��=:S��=���J���)�i�Qf�6\Sw���gXJz&[#smOF�0�|��7�q��u��d�e/ŚB�Ӎ�O�)��h�,H��Y�[��94J�>�9$�*݋Hs6V5�NcʫA:T&"���b���<�B�+%�Q���c�>��ޑ����0x�.0 *U55�哈���gc��d�"��@��Ch��!6
`5jF�P��=��R��i�Y�=�<�OP�ɪ�v��{���zc�돗C&��&G������^1��gХ��i�"�� P��2����4�+P���Q�����HK����E(C�R�.�DK��F����v�r�®۩���t��+"�9�Z��H�.�z�VGޅ��DNL0�W">Y�L����1����᫟����U0Q YXs� �j��W��y�V�밶������X@@���tWH6��	q�(�Ql"5ڃ:�SV�!��{��#����_�7�2�q��zWű�9�*�$��Y�q P����z�,��Q�4�r���|�5̹�M%�XMuh��au�E*��U���<x���(�[���vq���ԳN/���$��k)�?ӧ����@ ��LC�P�a������]�������{�Ph:Yd+�v����e�Kˋ��m��7����
�2y�8��7�<���,k�:�W�]R�D�y�]�ؑ��'�=��7h�M��g��r���τ��!����ޗ�Cپ�ߖ"���,E�-�mdW�I�BȾ3�,m�]��K���}�RȾdF�d�����n�������{��q<�������y]�u���u���N%������f��E�a��4qk�W�-_�!b^���۰(���f�����ូk�f��Not��	ujpHjqgVxsq�>� ����?<��BI�I!s�ک�{o��<�5��me�<aS����X�v���mК�暪*�ʻ���7-�ur��/F����?zfÖ�O%��)�[��B0m�J�����8�ݍ��=��O�b5^>�g���ə���c�$;{!'&�ܾ���]?M�5��������.�٤�c ^�$�Kn(׺Sݞ6���y�Z8~z���C�}��śO�	���S�s�VA����w�D5��T�>����x`���z^�\I�3Dڨ�����Ck6��8��$Ѥ��E�t9�ڰ�,_���o��T�K���Q�γRZ�9�m^*�'���iB�n0m5�ul���$c��*%�I�ۡ�g#mr*�����~l���5{��΢��K*ö~��u_	;&��3�b�qC?T��|/K��k}c@�6m�IF��N׳<���QW��^� ������a�V�1DO�S<1�Ǘ����f�B<p0�ݠo��j�Z�<v�	�!Z3%e8*��+�∵�X����<�0%�����Ԛ)"}(�
�Ic�7�9�g������L:Z~.��yV�մ=T�J�Z�y�N.��!�f����Z^y$v1�Ԯ��a+����9��h�
H|ll�rn��Y��)��@W�W"s�h!y�S���m�-s½�/����/�n��_�қ^�!:��(,5��-ќy��YkR�9�g%�:�WOl˃��B���}w��ꐅu��Y��`�qr��8}��
h�]f��}� �'��L�j�I'�ʑ�9}lY��rq��x:ؖ�_>���]Q�E0b0 ^6ӧ�mWc|���R��
��|����{+a?G|%�f��㽁���E�A�Iei�5M|���$p��]ro���UI���vЋ��5~���Y4;;9�ORhGU���y�OҚA�+������}��9�{|ksSSS�tC'�Q I1{�y	aښ/��[e�u	4�hA`�Z�o�b���ܼ����9^��T�N�2x��ě���L�e8���G�7�.|km  B|�Ln�������m4�"?���|U}a���:��e6�������y8u�~g����c���wnBk�wץZ��8�}1�B߫a�U��ԭ�Ǖ��˓��|k�|eH�Eݍo�+6le�Ga4^�+��@�(y;/�S>L�ti`���b�f7�'�TR83�\����"�����;�I���f�:\��hSa�*69���.D�3~���n��j�7��}%H�Fr)A�Oȏ�����5�~�i_0'�����v��(��n�\��o�7��ˢ�7`�
���δѥ�}�)���AZ�������ܨ_p0D l�Z��������P;�D�ci��v��:&������G��de����/��[~��<��mT�����(`�x$bl�'�VY�]PUE1_�(�)��0m�ɴa[x��4��o��r��蜱���B͙�pY���Tߕ�^��S��W�"�����>�]P�۰ck�Y/ؙ�&�Yi�&A2�׾�:�QS��?.���Qh���ߥ���iK.�����s+U���}��=#j��rS��1��e�ɻd���<*gA3�^��?�	��~g�ڨ���r{Q��IT}�����o��.o��X�b���׹����2f���N��N���~�aj���SK�>;/���u���)Rlѧ���Ŧp�͈�*�D��˶ʅ/��*�>���2L����9�L�6}���>���%��ϥ �ȟ;M�'���������_S-�i��Ub��O�ڔM�ˊFG̸���?����0���*�R���;�<�Q<N[��^���+�&���h)1�}�%ɧF��xg�O�W�_�W�����ž:ޯ�c{!��
�_^�v��X޷���9 м��Hw]W��`�ō�^a�grC��P�J��ݐK%�@t'xrl�,��+gY��&W1�uQ�H���l�o�p	k?��U��
��ak�~�JTD�g�T?���$&}�����n��<m���_E�Q�&�e�|*��5������$�<���R`L'ڙ-}n������h�*���4ԥ�@<)%e	d�a�1U�Isx�h�#X'۰�1�"���9?�u��Z�ЪU]�ᅕ]*�R�uZx�x�ҙ*6y���;ɫ�Z=M�u��Nط?�0�т�4L}I��is���<<�<fD�Z�$�d�����}I
�e1>*�<���J��b���L2�y����d}uF�~�*����b;�oI�07	<�a���z��u
��g�������CBv/��5CY�8�3����8oC�y����Z�6+�ǖ>ΣT�S�s�W�vli� 5y������iw��,��i\�y%������H-���@���[`[���҈uZ��ħ9��-����Z^[[�!B/�J�((%�N��M�C�bT�<Q"��Z��n�"10@n~s�
���TH���F(p)N����w�9G$�;k����o �/��E7���fN�u�-�wL@��hE�:?��l�*6�\�������>�d��L[ ��F�}�H��?�R�`G}��I&J$�a�ϛ�vL#�ܛ���+�Bi�|�A����X�|]]��h�+����A��0"���y�?N�zK�묓��#��y��(ͫ[��ް�3<rM���kc/j��u�P�p��E�N9,_�n��o���`�xy���.zvp$$��%Y�/�4�"�l��1_���`�'���+�ƅC��k������}�,��KO|B��5r���.8�܇k��N1��� ����0F�b�3�Ӧ
�d���B:gs�����qW�O���V�z{Y�V�t&���S�v	O&�6�_�ˁHD�=�mH�7��\4�p����ۊ�#^�8m���.TTTɶz�N�w��Oz����,umr�p@9�w�>��qd$������Q!�:�m7��9-������π�6M	�>=Id�n�ܗ��Dh1����V��D��&M��9\`q�n��ƛ2A`s�6�0���CY��m1�25;E�pw4���5�s'�b.�N9���� �{��@s��MeS;�P%��~��I�o�z�U�-�� I��@|,{�"4�w���>5Q����T~��Ʌ�W�c��Uk�T�������^񔧟N��:M�x�;�zW"�YI�/sxʍo˩�G�gھv8��L��.�_�$�h��Z�L��i�(\��s��(���j!By:�WQ2��eE�0$A���v�Ӄ��x�HQp�Aٖ��0|6�X�o|��h�lw�Eq4Y�,����u�������I���Y��f�ZUz�,�a!~�� H�o�gn��W��uy�_��lo�Ē��G��[W���"�pn�����#�m��x"�oR(uȲ�,t<kp!�/h�^c�eᑡ����clI�'�%�_+�|������G�Bw�ϓk^F�jR�^6�w^I�H�\C)���%STZ���L�3�~R��*A��o�3��U(I���Q2�� 9Z6� ̈́\6o	>�4�o�p��Z��GXwO+\��j|!���
�8z;v^���1��0����h�h�FӪ�9v�o	����#U�z�� s�	� =�R�V}�~���i#����Z��(���SR�U� :�]�H�P<L�%�Ѫp ��+����/U����ӿ�%8��x��VD�Rcf:,�7�A��D���/�C#&�m��*w�=�^�^����B6W���9_�����X� �*;��٨Xu(�y?��E̻֫�&�����������P:+�O�t ��$H�[����P�t-�kY�8��4����Oi!�׾q2izi��T�����0�N*(�ˎޭm�����/_��������)���sp�˴��k���.@;�ҕp��m�$Y�0�F���TZ�����y[nց�H9Z'V�«B����-�}�3]��K�(> �⤤$�[�P���*;��Fir��7K���1#|KM�@ ���"�����v�@`��};�T��F�`�J����lDۓ
��b��pW(�����b�jy�7�O��k�S���}�7W�sIu��ґ�(����7D���s�����,*1���W-���2��M�/8���X�	F�Db����ȳ��<�K��.� b�f�� �����Y�g�o�Q���1�h}>] �'|�!ܚ�֕W�	�ݝ$����8��M��v~����;�V�n��w�[�L���Y�`�d�חJ�X�Q#厽��&�Q�N�ir�ip�9q�7Q�1��t��β�$�6�q��|"�L��t���g���T=1��"�����}&|N!�����d�,�S� �k�6��Hq69%ٱ�A�đV��qp,Ҵke�Ѓ$9p�vA8�v�����c]*9�����H�k�&���/����B���`2|{U6�/�z]O��p��5/B�'����6<<<-�L�::">�X�y��(�>-���y�OjZ����^���J �����`g�0㶧?LS�)��b�giii� �Y��?'��F	CV��� �(�O�^K�^&�	�|mȃ]2cp�f��0Y[�؏a��"�W
�#��Hs=�|�����{�^*I?�S9�
��ڇ襣� s{�Z�n�V'�����'�B]q���o�������75�ɶ�'��8��#&R�n2 T]M�:d���[�m�!a�s��%�b�\�@�<�I��������73`&�����P(�a@������Lx�����؇3˼��U�k�Z���`J��#����+`�y��ڟ���v���a@�]��;g��@a��i}9���4��6oU���¡��N���`�n��3#f�������� ҿ��X;��W^^.lw��(��BO#,?�A�^�z")ēW�Z�� }��d�<�-ť�J�*�?/賘LX�^b;�7���6c����(�g��Ļr�*)����<�
�G�V�P8��I�b��,��O#� �ңv��@���[FF�0�#(W��rP��g���WO%�W�����[�4�d)6m�������J�A�J�U���⩩)��z��G/���[�$c�}w�F�=��=��ś�WXlV�33�^�b�9��,���ױ2q27�=�P�s�𢬬�r�D�&�T�9���/b�U��4����Q�X�>�ꙣ sF�6m�|՟����f��������Fʿ5@��ЁE%���Ha��5�yg�\��`��.6y���1�^�1�T����%�ȪԱ7KǵrD�Z+[�Y L����`��X��&j���u�G6`�1 ���lF�9���0��uD�w&�Ԣ�z�@��j�tz����%{� q肨U�<:Ќp���{R�J1$��nO"�l��Q�a�p����μ�}�J�T�ej�z2�=�A�k�{"��B�sh�f�x0�w����ol�7kÕ�Ús�}p0rMa��أL����v;f ��"�
��|}}�oP�����?χbV-�R�ܨU�u�Ȁ�zt���"s�|��k� �~�Z3�r��n�'S�W7W�ws>'�1(+��9-i27Z��8`u���w�`r�b�@RR T\�ܙ���|;=,	�������o���i���̺�=��<"�&�l�;C�ȧ"�]A��ٰu�p����bm=��XQY.*�y�fJ����"PZʿ��a�{�����c�.{�	��~���~*r��>&���ӧ����=�^�%c�㙑�Q/��؎r��e��#s�hq;�E����WO�yӂ5n�M{+������U�
��3���Ӛ6�4�FG[{�0W g�d߽7�ܣU���|J��A��Y�5.���DO+����k~vI�×Ce$���^j6�临�^�>������h
�g��ۨ_'�(�E0t��(����ĵ�#꼳>��`�Ys��7)��H����AR1�W�{�EY�����*) ���Y���v��K�w���1��;2A������+�)r-�NW�Wt�==@ l�>���x� j�:�X��)�fQ�۷y�������fV��=��)�bmy`��p�l��7��B���� �R.�c�q��5gA��I��x��-�8
=�f�JX��E��W�DϦ�0k9��s"������R:<5D�xz��ꐟ��ڢX��T��c�֗8�Rw������jǄ�Ba���F����ԌKġ$m���]��P�����β|vp��m侩��	R��[#�C���0˯��� {���'
����'a(���Bɿ�|;�ٹѪI7s�EK G�9��\M9�X�'�_M�1�)��`����D��{�� 2�Y�\�L�PX0~�!�-qZ8�F�yR��x]j��Q��!Ҁ-RZN�k1Ț��s���ʔ?��)3h�e�%!n��K�1������3^�|���ر�ҕGj��nWŻ����*��i��Y�2�3�v�"J���.X j�Ȼ���G��{���������dU�Q�O�*���,K�����ٮ���-�r�x�u8����w�ނ������g�v��H�>J�7N���1Ɩ��Ο$��6�������j/ʀt]��<;5&爝�]�h�N�n�ۜ�ԯ�ԓ�,7�lߙ�����ÅZ`����6.Z�ꖸ�*���G�� �)m�~Y�l�����+����������՗�=��ٙ���r� X��3�-�i+�*>�
����r���d,����^s$҃-AЦ����b�e�Ww�UT2/݀?����$��p�R�E�.t���)�c��\�G��-&3��C|3JEL�N�����i���J����t%��@W8�q�D�β	�PN��tuE���=:��h�j��J%����XH��6	L[�xiEEa� a0�(����E�����2�2U����A_��������1�mil�=�ב�/�[y�h|D�����O�oV�,�H���n`�e u����*%[@�V{N�<�L����x�ߟ!�C��G˝����Ƣ���Ē�WF*I��JIF��r�;��{�
���u�R@��9XQ8ο�7����)x�T��yT�>v���I�%gi���4���`�x��Y�[d.��ZOp^TN��͝͡rW�e�	�pt��g���-��P_1Dn8���Ӝ�e�|�����.���7�c��tL�-��#�A���-ߟ����Q0zn��S#�Q��c����
	��;{V�fxg��}�Gb�}��͡Z>��U�Slo>��@$%(�׮ ʖoo��L<�×u -'��E��P|�Fь,5�{B u��5��pttĚ
Z��F�`���h'G������o$p�%b�.��/��'��L�?��$`xt��F��!�n�끮����'{
�� MҘ������? (إ�˂7\JEE��OC�B�[��n~/�;���9�P��g]8d��X��Hџk���I2��o�c�;[-	*5����6���Ey�M�6o������<<�X0)��]�R�>�����xv�)��I�h�'�����t������j��Gih�P�P�91߹S���ԈBL��4>?2�{/���G' )��a["s������׋���O�ܻ�x�BJh@:%�wx_ �_�@��"N/I?>9�V���i��+�tZ[[�em�z�y���]]W>ݠ�"��^�L�����$�7�v�yJ�*���LД�J��Y5�;;;ؒ������Rz��|	����+��E���Y����������B��<�0���H)((�V����{� ����w_�b��1�"��K���_ ��]*Ӯ�r�֭�_}	�/H�{ҵ��� w3�f,�)ia��`�E�Dz�E!�������TʱTj^L߽������߿�p�i�g��6������1� X�u��衲"�6oCТ�����Sp�j��OI�����-W�gϞ��� ���ݐ����RFz��3��K/�
�<t��c���S��%!$��W=gY�T`�6)!�9�#I?	2k�	�N��S�Ⱦ��::���5fsl�[ �.������/���sIu�85 �~��I����d������<�|�4�-���Eރ-���}��oe�{�5Q4Ȯ��y,�q��q��O���+-Fzf��a��������e7@���4m��6�3�_O%Jt���Z�����b�����U��msh�!�����%>������020 !y�\���+_+Q����N��@�5� �)��B��y���'�|| ��l��=���R7�%~�J6.�w�j7l��t�P`J]*�lUf�ł l;���&+�>���2z�g��y���/O����ZH�2����O$���_�dccK�-}a��ֱ!���,���/�ډ�>��Ă`��,^;�9�,x�ω8�ZQ0w���i���V�|U򉐛G=gG �G� s��/_:o�& 
���]_<������d�ȣK6�"��?3C!ȫ(��YY� �1 �i��WP����� bU>�?�َ���e< ���ԕk�,��qq����z&'fy�t�@���'���V[�tq%�{W�J��׼�n��_X�Mvn�L�����#���*�z�933�e9�RW�����2h��h�8t�*�l�E�c ���ڰ����R�^Т�bk̗��=�&���r�
��P\$�jh�<���-�}mR�w�Zl���� W���\���q��H�� ]����H�����zl�E�i��L���?��L�M�m��@��Y=_؆fX�՟[/(�t��DڼNlr����"��Y��7PA���^����C.~�7%�5X�$���lP�˃��o\���횽��� �ET!�1 ���S}��BBc��%��e�z�ak5`�|�̷(��<I��w0����lU�+��r�c�w��%�g�&?w���"�677�o^Hiz��	�%D0��\�h\'�n�xw2�?������cg�Y�C�b�?�N�d�3#���5��. U��珬u;�<4�*F<�	�x~#8�k������Ǐ�H�h�U(�ʻHx�2�)���ܼ0��*����ΛUnA
J$��T�Tֹ�Z9���X6fb8�X*�7�Qg��5a\lbok{��S��PsSy�����}���5��K;��}�SQh�o��@�!BU�fȧt��V��v��X�!�]BѼ���a�-�a�9�����y�sO���U�,�x|�m���>�;��Ɛi�C�W��֍��I@1����w�9Vi�)q���,I˞�;����;�~�x���.�TWrFAW;���Ms�T�|7�|s��~��ma�������ߠ��&T�Dn4bC�#?ց���6�F�W�� I��XK>�s�r�+�#IT�k/ī�J�H��SAHm2Ѥ�{(�Gk�r@�����
O�;��:�w�|f�����`c�`�2i�+��t��bqv�>N�0U�Yp�!Kbrӈ9	�m�ƨ���U)z�VL{�}b{�.Q�}Q��́���سx}��=+��.�������3��x]���7�$r�;��P�7(�+J M�p^�7��b�"��B�Eҷ.��{�~��C_���1=oj�ȳN�7�v6��6ofN�WD�{�o��,Yd��k���U�+�{N޼!Z;�vÃ_qW����_6ȷ��>{� � �.=�@]�tm��G�t."�q�틁C�H�(|���M����ϳ�1N&
�@��VN�~�]�������ԕ���r����PČ {�Bp�Q�����{P��
t��9��L��鐫SB!�ӧ��k5��q�L=�筡'i�o2�>��4�d,��m"�U��n�`�'%<��E,�M�;H����ǚ�Sk�е�d&ocW����d[w$�[&�B�s����S�+4�q�>��s��P�6bf��-�o߉M�l%b+����+2���7"���y��,eA�O^�x�pR�ٿھC	���wnv bB!Ӌ���?��4�f�-��$IIa7��ڎBfW�z�<�j����1��&U�4P[N�!�nHjG�l�s�&��!�@'�䢿S��ڮ`��f���tYg
�X�=���47̕�H����6�K������!g�Rj��Se\�Z0隷��VVw��B>jU��u�G�m���b�w�M�)~�u's�2ᭀO��uTgJ6�.�h�R�R�1����|i%���7Mb aop&������Y+�P��#�U��m�-��v.�H�5�)����c��'��!^�nº�5�v�JEHm=[$�}±���3t����"��������ϲ�AN�3�s|���4i7j^5Pq>ZO���&Z.2�;e�J&K�n�O�^��)m��b��Q|��Ӓ�=��?�^���/����$��eñ;�"�z7�\x��� P7>?%�v���^�@>&%xe��;��pJTs�
\��������ǜ_�y{a!�v{X�D>\�<���QI�~�-F(1S6��4S�%���}�h��DF�K�!@��Ȟ��k��-��[��v�����=�*5����VEA������h��[�v�O'���+9��v�aD	���h�Qea�U��*�Ͱ!���/��`z��:73���=_q���*�����M�.��x\$G��\��%)�у����V�{�V�^�˙9�W}�p��Oa[V^eɕ�)r,as�Z��+����x;t�6p%		��׶_?6��f�r�T0�r�:��o�P�Y/�V���3�sۘ�HH�9�+��Lo���M���;T(pF���E����"3n$)v�!��^m��]g��J�Ir�y#'��!T�Txy�t��sy���9���w�K����e��o�}T>���h�8z_��#B�__ʥk���+���������z�7[�*M��k�.-M�oTk�/�O+@�@k�v;���FIDN���Eƕ�����:�@;y�Qo��pv���'��M�]��Ic
�ߑ&���x�rFL<��t��8NhG|<vő�O^�ͫ��HhW����B>�$��/?�:%�K%�?�D���4���|���`�ؼ���E����3!�g�R�:Ӑ[rEhZ�͖�1�M�i����D���/LP����������~�L�o�w�,9}|_�!�Nuc�!���:jO}
��'�=rW�h�%+A3�h}������O��\�w�
��U��#��PEDQo���.��NS�,X��.,wO����ڂ�Q  ��c�[��t���V��mo�O�4�S���3�Go��0�tQ@1�9T���Kx<'����f4����'}R4B f��7��e�x^�=�X��י����?�G�{�� ��f[)b�B�y������`Kc�v�(hM��w�O�i�"P\�i��H�!�{����_q>� Z�� ��'ϨE;%
 �U�v����Xq�z�~vg�T���w1ֳ/�P����9_�Z����&m��3�>k+��$4�?a�!��rN�$����N��z:�6���9B��In�e�i�L楝�hT�Iq�������ν"�c/��2]®zZ��C��h�:?�.���t1��w�rY�-i#v�r��c��f��=\�˾ɮ�C� ��v��7?N/�IM�<�C!
���i��3-�F�0��o���v�2�Ҵ${����0��̇���R�]lL3?0�����Kv�:j�
�>
̿���.,��b��E�B��i�v^��T<��DJ跚�t�zwψ֙�9B��X���L�o}њu�.3G>�H��Z�9k�G�u�M����ؖV�����T�r�+G/ϩ�:�Ϻ��XD��T�Q��d��y�p�T ��ں���~�sx�je�}�$ў�B����`�Bu��-.�z67P�1ዩ@��&޿���6�T�&f�9\�maLr,�٫aF�4�Z<h�G��F%t~����9�L�rS�,��cK���:G9��F޼z|(i��Rח������BK�YdfLD>�ɐ�^�1�6ƛA��
���VY����CB�L��*�����u��?���_U��y�c�\���δ���i����_�O�2���ޥ�oP]��G1^o�u��>f�!�S�o��@[���ě��*�6eV�_�����.*+��Z��Mb���7ʾ~څL�0T{';���[���>�	�����h��g���f��r���:��ʙl�t����5B�<���9�t�o��l�Doɘ����,��8Q��ax�Yc�����r&�>�߶�'u�z�[x�$��#��*AD���M+���	VR�L��p�Ж��E��B��ʀ��y879���щ*,75F���L%o}��X�o��WAv����7KT��:��ݑ�Lo�3��0ŏ
��"�6�G��E*K\�=��+<l��P��1~���͜J�k��j�^�>T?l�Y������i�Կq� ���yHZ�|c�����*��{������*�]�(���Ьbe�=��,U�:��|ྴ��*�|'�o/���Z���N<������K�>K�k��gI�!,�Hd��ʫ��7M_oL���Io�(�	��S�sj���7]x���. �Jzk��Be���e8�-�^��O���ȩ8�NO�g�?�$2����6���O}�3�\����n|��]�_��G��{�i��x����KKW'BY�CN�R@㑀j��;j$v���2�<��`
�)�d�	��K�����9�_sm�pF0
�P��,	r�M�]�p�+Z`b�_��d�걦�l�7��n0_:�u������V�Gb��^,��ty{.�
J��u$�B9�l���?��Հ���7���×��F�1�O|"��k�<�p���S��o���P(�����6������&���!h퇩4�����Qh�����j?l��k���w,�������/7��p-N�Ev^� ˕�����?
����}�,A�:���=���dA��Jƾ��@+/����p�ߵx<���B����?}��}�*������o]�����g"O��"���|��@�O�N�d�TQ(��&�����Io�ǹs H���[���կe�Ћ�_򑑑.|k(���X��!��縡��*��^�Gr��D,fh���mM�D�@}����WX:�J��!��phM��)�E��'}�������[u��0���=$s���]\l��"�obuĲ"���A�k�Z��Y_m,w'X��(�A����*�q�@���.x�T��l��+�����(�tJL"� ���[��A�<T�*���g��8,_a��("��pԖ��ќL�0�R�p!)�j�*���{�^��;(��u�"Q���:��&h��mN�cZ�&�~[~1��^ú3����1�����ګ@���ˊ�1�V���_��Df�D{=(���꽆	������������w�C ��̓��Z��g�ӗ�K�h�>�;j�2��z�;�uS7�� }3x�'TD-n����ɬ��^�|
A�A|lC҅��YuG�3��>�1c�xJဗo�=l�a�b�[3&(�r�ۯ�m����SO�C�����u~M�;y|>�����c:w����DSc��_�]J�1%}E�J�z���20�$�4�ɮ���>��j���Hg.��8U$y�;:P3��H���8���i�_��J'p��dp�Ӟx�M�\���ЫY�RE(��z�m瑕e�/�M,4È$�j�{Q��"����(dV�z+`\'�=I{��Ƴ����2bWj�H������K#��7%7��=�
�W ��
���ۓx�p}ͮ9bؘ����l�&v (�������\���g�=�~�(�����:d�A�@"�=	�e��y"���n�B���N,)K���G�;���	%h?
�-�r���z�@p4�Y��H��8��v&�<�(���U���O�`�ڧɺ����,�K�oG�b@�N��g�=]w�$oGD���W�><��+2;�cͱ����F[�H:�������w���C�½f�Ǐ�7ҡ>axj������"�Z��c�7�OjF�و�>f���dgw�k|�3�ξyq&(�Z�`q��)q��'��xE����
� �ѓ��g���k�����\���{��������߃�.\�}����m���L#G���?��"4OfR�k�b�l,��������}n<&#��lN�yTy��ҵ*�ң�I}�jZ�{i�d��p2d������ǮU�D��3��-�w,��Ê�6��4DY�_�^��g>w��NV��)I�J>.�r���B���ndP�mp'�똱�0&�w� �6��uz�|o����1d���oOY�OH�m�I�����f.�C��T����	��ËJV'�='OO�3�0>�w�M2O�4�cBJ�s1�A-�r�Wl�c�}Pv�m��k�^e'�2+�/���r��seO����X�f7�?nm1Ⱥ���W�͌&2� !�PP��6������q��\m&ˉ$ ���O:�C�f�4W�z����w�j����zk���F32�� U���\�֏AY�iozf��7\7��W�L�zE���~dȇ/?���1�� n����f�L,�5O�h#���e�?=ӻ�������潻��R��USY��WL�v��+bf�7�v�TM���g'L��׆�f�����\�����k�����ݕ���R����$ܐO�½��bT�f#�{p����4%5�_��5���_��5���_��5���_��5��li����~��{��D��@Pp<�����c�Ǯ�ɷm`��&.Է?4�'3����V�4sU$�HW\�����xgg��L��~��ge���A录���nQ���_ʩA��}
e��`��l�t�������vh��f��B��V�AF��c��Z��L�!m����w�s�)dV�^�彏o&���g�~�3T�_hOJ�|9{�inߵd�k����YJ'����tj˸vv&x�iCY F^�����y��ڹ4,qe"d�''1de�RX�P=��%�]��� �F��V6#k��Ǧ��3ʭ������
{y�2�ۛ*7J��.7��x�"o������\L�j[\$����)��d&��Lh<^�k��Z\\�n�{�h���ǱZD��5���`������{P��XH��ٴ�~"���4.i0x�.v��e&qke�n�C�MZ~9{q��th׹qY����=�>�$��vNkRn��K��EH +B�򃲌��?-�W2�h�O�P��4�P�x���ij�.ݾ� PK   ���X��6�B  �  /   images/ea05fd3c-afe5-4b36-b101-0986c4cae35e.png��s���b``���p	�) ��$MR,鎾����$�����L�K@�Q]�S:PP��5�$%�$�*�(H1Z�X���X�[���[�ʞ͊�!7?%3����f�;X�<]C*漝�!�*q�����x~μ��}Ukk�Ƭ��W6���z��ɸtU|] �2U���"��y,�N�K�,��\2)��掛o��w[o~�y�M�L͊�����hom�y�̟o���3'VOן{��7�S�S&O�Y���I�i��N�~����
}��'+�?I�>���q�f��l3��4o��W,?*-o-�p���!�2Dh�S�3���O���sO���gΡ���G P�o����%�2_Ż��9�=��tiȱ?A����j{<��Y�����������g�ZT����}��ձ·�+�l��?-a�1��u}���ˮ�2a���K[��n�5[�w�3ެ��������!��4��˷L���LN���7G�=n�+��L!=�~����J�R�3m��/�r�E�5�SVs��KGj�����ҷ�O��_���8�7���@��G
E̒;���g�+�(z�{z��ݒ!^�w]�p�z��[���;W��;�c���)B��.��V����X�ua��̕72���j�?��U��U\u6Wms��Ό�:�͜皻x]꒢��+�:�v;kѦ]<WVE�k��k�.g�6a���,��ཻZ��Y�ND{���-��L�&-7�U��}���V{���[]��X�wئ�C����i�Vw����?u�=fs���I��ji뱴���9.;�u���Dq�
ߕ���:^����Ֆ%��ڋ�D{��=�r睯�褷��{��d�sL����<|�����^1��`��G�)��f���^"z���m�Ov)�]��x5�1*xꭐ.��/gO>�DGƲ�C��G锧�dL��������jx�Kc��r
m��`~�W59鉿'\V��^���yw�Xu-\t{Ҫy;�d�K%����]qv��̲u����¬�ݽI[�K�?Xx�[�4����s��]�ݹa�������ST��&�Iը���n��ޛ;�ٿ��]�m�@��@,�*m�����t���5���*���h��F�M����V��w��X<*�b��Z��5�c�~�}W��L��|�bV^5ܿ����[������,���~����X��&����|��u��+��e];������i}�1+3��,�ҥ%?Z6=��Y�J��e{<wfH���Y�@���hJS�����_���+N?{��������Y�����u=sG��W���{��6}r�.�jΏ���,w�[x�"��e�t�sY�� PK   ���X��@�/  �/  /   images/ee535837-a8e5-4cdb-98a7-fed99fa44d94.png�/pЉPNG

   IHDR   d   p   ���   	pHYs  ~  ~����   tEXtSoftware www.inkscape.org��<  /IDATx��}��u��a����� �A0�)F1HbI�H3I%��-�N%��\W���]u���I.�w�h�mӒHST��� ��`s���g���3�3�0R|�C-f���_�����=_{��%�h@�%���A.2�D��.�"�K���A.2�D��.�"�A,r�-��@U>�h�~��(P�j��B�r�%�|`�C�u��:4�h6kN�B�lv�2�I��l�XC�(����3E�9�A����,����� E��k�=����|�T9�҈��8Tܰ�:f�Hgf2B$&�ۡ������O��T��^�c{W�NL&�|6��2�� <�L^f��F��v��l��������9'�4�ᴉ�{�8E�*�amN?�)ڼҟETT���C� X��F�߉�i�x�W����bg���,��f���$���i�X��x<m�X36w����5����+�AX��Y��uȀh��.�𓇧E��H�L��[-x�`�'R8D��KƉ0՝��;H�l�@�!�rC���"��h{��s���&�5ku+�+�CX��L��B+�$�����kzUm9�FdQ_׮
����p˅A�CN��xt�Y?y�b��ʳ{8��S�z�L�맒�{p�^q"�>Ofߡv6�R�˅�� ���븅*A�(��BC�WDrҸ�9��d�~Qh�V6���q@JpQ�R5(E�YʃI*VQ�b�;��MS�8ЈXP��Psn�	�/�5�VO����ߩ]�j��o��e�ZGe�N���@p|/�_��Z(8������5t�>��S?����X�`��݁T��p���q�ߠɪ>���~����ij�>\�q�����O�mDh�m`ⵞ~���^�
4�9�6|��#?C��n:U�������w��u�7s����'E�Q��ӗ}���P
f]�qA	�����ȿB��Į�a�]�_�����[�~��p�g�Z���y0D�I4�
o���h�^9����7z��=��T:�����/�ĒB�|�Z0�n^+W�4Wp$�2R��'��#��cj�;>�LpU]�ra9�o~]�݉��%�7k�ɚ4���>��ZQs��u©k0IN��������ʂ���˥ˠ&S9��Ǟdᅢ�é��q�����Z�<o�B"G���^�0Y:c�$���/b$kU8�a�əB��C�ɳ0�>��A�a�ND�0M�w�.��	��TS�a��w޲�{���4�Y��DϺv�aŊF����K���m%9] �iۦl�҃ɩ�y�r[R�8}yj_�ӌ�_�T*�g�?�p�|I�1[�n|����/�z
�12{g��&�~�#��#���;���'l�X��Y7~��]A�85�W��j)���\���C�L�d�f�1�
`�df����4ͼ���ŏ-��PE�!���#�|,
w���X4'�$�T,�3��=�J#�������3G��1S�q�p�	b�� ��}�Fa�M��j�al����'��<�*w�dE�L�`p$$\���m ��,f�gRxkoJDV��_	��,3��I���?�<��LƒI�'+�c���}���ӄi�v;cW��􎜘�Y��%�Wy�.�R��̻e�����c�g+6�`�"X!r��OV�����e�+�&뉿ON�k�U��r�n蹸XZ�9~Q��A�V������@�Ri'���^� �ALQ��|Q�	��p�0R�Q����i��e�vN87AX4(��m�`d�.��XS��q�UU��R�d�ᾛ��yMC�e�W�%�b�vbӽ��~�467��d�6_F��h��8�̌�si'�dx�0��ay�����[���`|�}d���g���>Y�#�;��c����G�G��8Z�="�בv�m��K��S�j?��٘���!6��\�D�f2볯�AyGF�}����=�������!�|I�X�N��N�U��M�j�nZ#>D�m���q�L�Q�3|��sx篒U7R�nzZ�i\�?0��3dZ����������ƻ�>����-lߦ�i]��c��hM�JK���g�u�q�'��B����fNbl냄��ey�s��-���;���b�É��Y�h߂�RX�K�"��k���\̢-�s�Be��Vq�j�Xi/8�Q�):�h/�M}s�ь���4��SL$�}|� ��P�]b��M@�ll5�!�9���{*�͊o)N�����ng�,>q��KK,��.�E	t�f�%G�%S���C>A��s��Wl�!�3�$~�"����0�ü����hB��3:k�pfm ^,����&'�����TU��K��p��f�Z�(XRiq|*m�;p�&��d��T��S,�ҟֻS�`A�9�pi�/~�tc���qlFw����X��kV9����W�󹯂�T�Ԫ��|��u�l��6$��E9G�14��ɰ�J���>GY�}.V���"�l�T�G>����J��|�τ��L�#s�s���#ٺ3k?�恗k2�ܲ�pq�UL�eXb��}J��X�-����|�u�ZL2OC1@�V1�z��(4,��#� B���͢�8����Mɼ�{*L����I4*��HL��(��x`{�:T[��K8f�p�tX��G��c�
�F��>z'�,:p�l,�*��	��Ń�]>ɂ��s8�TR�ln���/�y�NJ4��#b���U%8>b���G��F�r�q���v8$5c�x��J��j�J\�y\�Q	f�t'v9��)����+�����vCq��gpv` ^���
mN�dt�lV862�������a�U;��穘���C�,�|�"J[7oƦ�6hV�
�s
^��6��4V��᪍k��1Ib��C1
����p�
�b[��h����k\���t�=�q��p�'���rH%3������ۜP�̉#�N������W�"��Qr�r����,%Ϙ�����#1��3å�L�,#�;g��J��¨��Y(w&Ռ��/W��r�i�=!"���7pF����B�����9~|/Bg]�IJzn5�8�`��`M;��L���p��j��c���A}�` [�Tm�¥���qt2�4'��~'R���A��k�}0;��L�%\1t�Q���fh@����H,^�^�'R�n��]_nG:�P8�`��d8_�=Ob!(�#�LW�Y��x{�p���ű|o��!����^��O���1�����܊є���"N��A>��]�D�x�~���-�e�UkH�{	8W;����w��������.��Y�K[~|<?YZ����ڊD��l�g�u2w��ֹ��?����B�&�⣠�ಮ.Wr�oV�)���u|lz&IlN򵨠*/t�H�^jϜ�(��wf��1V���AF �nϓ|._[]O˟|.�U�/�$�d���!�iJ[E$^@�h�j��K 9���USpf�N$T�C"�겹�*'kJ?�������k��3� b׮]8x� 6n�/��s�M7��������7߄��a�^�G�l�,ޓO>	]�q��w���C�����{�ASS#^|�%��n=z��������?��^ۍS�Nɵ��2Ye?�s����@���as���/��]�Tw�W���F���t:e�\.lذ?�я������̙�X�v-�{�y�����7|���
zzV�	���oࡇ�f2S��3g�!n��#8~�#K��79���k<���,���>'׮X�}d����8q�.4Hp1m��U�5�(�-U�$���)���D�;��.$�6��g$����<S�3��1��s
����������z+2_9>99���F�&!�֭[q��!8�����Crc��jii�}���p�<�\s�������!�\Pѥ|cbY���8�47�m�땳�)y��1&'�9���恗��H֭~O�Y��x�1LQ�%��=L�r�����i�G�ƦM�e��?�χ|?��32�l����d=�ײ��P�={��_Ǘ��%�\ً�۷�9�Z�
;v����>+�\(���c��@i���Mn):N������g �:�T���8�\�4��זyK;X���%�g8�Y�������"�q���K;+g��/��;�C�?��O������z$	���[�A���9x�N�>�x ]]]8y���eN�F#��j�ݻ����E��u�]x饗p!A_I��0F�ǳ�9ܹ�Y���_
��a�7�����x���YTmq%��*�7�Hz�KZZ[���g�c�=�5k�H)�����|T>y�Y�3����|�+H&S��yvk�*%n��Iᐁ�!��?."���_q��Q�dǺ�	���kYt��:������L��W���#ô��yl���� �qH�,�ߧРX"��R|g�`I�����e���cǎ�ċ&�422R������̄�{(�*Ue��ה�e>gjjJڸO����e�U�Z0�\b�+��S�h�ϡaK�O|�Hڄ�T���q�X�wWh"� H�Xs:d���x��YԹP��
��^��V�Rf�z1�!�+��LMm�O�1���$����%K�ԙp�"[��FR��r��$�%+�|G��
z+�%��:n����t����ӋgBoی��qq+ �+«o�b�z�s�zf�l%�:�E�}��>�ϐX2��*\�.]�����	��}k�y���ly*����˺a%����[���
�bt�9���ŋ�g�yY��̓��,��,���Lۡp{u�%~G`|?R�����VCYI��L��dGw�4�%���sq8G�1x��G�'N#�yF�ʗ�)t�6��˻c�n�dM544H��l/�����ߝc���p�������}�?��:���(�O�fUV�_2���C��8�Y�,?ĲE3sFٜ-Gs�;.��)%�;�9����r#e\��a�8V�?�R�^���ͭ�:5<{2L֖�_ �=�s㰬�;�h�ae���%a�Y��g�b�!�J�o�?0�3��D\�v{�q�F�'V*����p
g�m�f3b$0����~R�4�qd<�]�c"�`1��ܿ�B��c<�����tև>�,�l�$�	Xy�+V�]U�R����� ���oŉCPZ�k����N���ޝH�[�P���/|��M� ��>�7�Dxr
;��ħ�S�"*�I�ܷ��/�?~ݫ��+�}H�9*e<�O=�^��s���_�4���Y��xc�a<�'h��������C����9=2�o�ݷ�9�x�Gq�έ(���P�H��_��������я� bd���	�|��[��?� t������G�`�a���-z$c��3T�J[X�M�ch$�[��)8�V��Ki}Dqʼ��8��:p������cV#����t���[Y��<���S�f�?��w�eF����z="e@�,6b�C��y�������{�&-?��߉�߼O~���`BK�I���Q:�h�5h��-�{��i�@�Ӯ����y��<|5<��ਠ�-��d�	�O�|i�����9"p*4�W�C�o�a׹9\Dȅk�u�V�"���]�K�6���^_�/βwym`t�5�$V��5�.�|�y{���ܻ�,ӎ`��*�E�F(��,Fh�J�<�2�f��e#Psw���c���&o��vr��&��A���9�+�j����q4�ñC��@���UUx�X��bJ_��M������
	��,�b^����E>�U8j����9�KK����b��B�?W���>�:ʒ�J�r�����T��^�^��_�Z8g���ͱ���"��p\._�����w�"��9M���׫�vI����N���&��P�
��YT��@^8��W�޻F���(�^?g9A��-�bf�9�\Vߛǐ	���)�s�Q"ʢ����@KG0�Б�u�> ��5;��"�����r8�j遊C�<Y6��҃;w��d��l{x:�������̼��	���r�b��3L��V�@��$_:�H��A3�6A��xy�1\}����?j��
6߰�D��6t��8���V<2�����������(���/s�c�~HQ�m�7��$i�U���lV
<�k
��1�X�����YxS��
p���
��y���h��X� 64�#��ĒH'R�"��'7�O8u]��
d�eMŅ �FY,�u���͋�� e;z��''y�L�J�L"��P�x�'Nj8;x�'��爫I�s��0�^��3-g�,�-��z��`��\Edqe։B�FDy�G"NL�t��!�و���xah1?Z��θ;p��I��Ys�cd�x\괬Ҋ�M�6I�c8.�U'�a� ����r�jطo����s��Q\�266.�4^�;w^Q��ũ�~ٺC'���+�\2�P�C����`Ȩ���P�oC�K���v��~:^�PK]��iBs�#O�����c���x�뿋-��p���s�o��{ﭜ3A�g�?�uS7�G�з���o���+�9"ԟ��W��ǉL:�D6�G��j��7��Hq1�8v*�G��]�������	x��]с������7��)�X�d������]v#�Ȫ��s����a<⦂�F�R/��v���m�hkm���d���hBgg�~����N
��я�n?b���t>���6�Rct"7O7p��z���Ds���/jey�<��� R��?Ě���O�����;�H7��X�-d��1|��&���z��B)6uaE�>��C��b����؅��:;��	KI�ps�8b149���)�r&ڻ.�w�D"����)k�=�đAf��o���F(�>gV�B���$\D�'L�f�Q ��Ŝ�-��u�&p�=��[9�E�sf+���F��"N�!�{���J}˖-��/�N%��U���N~���ۢK8?W?����K�x�wwwϻ�C�y����q�����;?�ή������]!��Šb�2�JN�^���*{�&�)�dg#�	�r�B@�Y`)��2��Ca��8��,����5a5�B2?4����ŀ�\>���-�΄�eK+i�[�������$[*f/��ޝ_i<� ~:r��~����u�)&�5�S0zb����l���(�������ʲ�����z�Y++GF�_%�:�:]x����������>��S�XY�E@N�.�p����ys'[Q\;�,U]���u"�Ek��q���T��gɬ6;�E돋l{K�l2��Q��T����q��hJ��ld�%��_�,�X�N5�_^1+4���y�W <C�,H�_$��7F��Rxe��S-r�p�a|&��<uD��yӄ�8[�X;,��ՃV��e���oD���3E�%�dB*h4=>���)���@A���<b��=�G������_��>�������9d�MȌ^�'O��a�TH�©�Ӳ��9~�+�^1�����Ξ8lQz�&���/)�|qy\������PNG�rVf����BM�c.�s�{Up��;��UD��3�eo J����P�#�e�<"�±8:SCx�<v�\|3ߋ�bˬ��s.���������Y<4�v�zxv���
d���΍��x�r�e��P���2p��(��?A��Y�3���yø��銕���kde�2w�<n
����$��q=5�鸆�g��}q�R@zrY�wU�H�f���beI��]=��LbD���M%)��_{=�?x#���Ѹs�1O�2���u~c�!o@��G�ᣔ �?)m�(5�O��Y���3�w�jpUqv�4L���|O�0ݝ�Eܑ���ԯ��M*� �?8~5YN8��H{:pV[�p�M:*z��a�/o�"��qb:��쥋etU�+�A�J��55��ź��o��,$]��A��!{��¥z��[t�]�H��-mA2��.�]��\��j��!�~�y$rԦ���R0��F8�8�AևX�/�C!cB��D}[�2p2鮍�4;T!����RҺ\�+x'
^V���v�ݞ��7��la��H�^քM������Y�@8��u�͞F���s5�0d��r�h��:O���TJG��6�XL�%K���])�I�L�/8�V��?���o6.��ӵ�W<��ǒH�,�Z}ǲЖ1<�\=�@���"�[f��b�X�mk�82�~�o�ɗx�������8�^�{
[>~?����[�.۵�t�Zx#�����1���-�ۉ�D�E���<u~�֧�������x�,���9M*/K;�.�]x��J��5�X
Xw����_��Υ/����&��K!o�+ˣ�-đ$��VW�Bx3D~��+{N���B���TӹV�'p��UJ�Z8I�xѿ(Q��h/���+����w�%C�:���%�.wr��Q�=�z�~���\|�#��wR��ԖO��������EVͩL3������	 p:�l"��DX���f�>�
g�Rmˉ�ŀg"[W#�h� qc�rٜ�)��n�A磇dD��$��o�V�U�>�����5)ܽ��Jp�S��އ���mx>څ�^�(8�%9�^2˂��H|8�Ҏ��U�.�Y���p��~�B�>r�x	ݱP�;��O��-��'vv������o"'}�.Gu�I�49�.����w(S@�(�B��(l����5q�J����IF���ɱhp�&.�,q'�ޛ�r����1����7шhM^R^^��]nI���X���Wojö.?�t�Dƾ��я�W���o�������VЯ�l�'76�S�m7���OϤ��ި|_�(L�S�}���uuN��p*]�3��x�d���Z�BA���>/>����)�f�t������HfY�o����&��v$5�ʹd��kf���v"j)�������]M���u(���b�������7wY��8K����|u�ւ<����;��xp�K^�G����jf1������d�I���ʶ~
�49�_�m���7���օ8�u������׶��v"��"g�MoW�4`c��pqSusʒQK)/6ζCTU2�0w\�҃Mm.�S������t�~��||]�bOdA�x~�ǃ���������K�ќ7>�.����=�Yp0X��ʎ ����xʋ�\,;���q�z�a���x��][]xx{�\���/�n���]W�n_���#��f]�7|�v�b�7��q��Z� �k����r:�`����>��#�d6_Y����,o#���q�::�	2��z�ܰҋxΔ��fw����C�ua�t�V�1�ݶ�K�C�Ů2�o����h��Fn�����M�S%��m�FȲ���v���^�d@��8P���,oi^<Q�(�@]���<���]6;ۼ�������b���Ek�u����:h�����m�
�ktH_s��_9�\f� �Xk�u{4��~v�]��E�������r�"��ŧ�Kw������V����٘���-zd9�b�Xe`�G�:�Qֆ��2���<D����5�Y�sїaB_�3�AT�F��e�4S�N��^�V��˫ZC��5�#A�Ө,G�*�p�u�HE�ir�K�d�n���χF�J9gA)Y ��G����d�z���?���y���2��;Ϥ�,	�,^`Q����IZ;�46#�Ԟ��Z��&jy#K�!�ҁ���,=�}X
��ұ�-T.3��7؂L<b_ˡs�*��z�v&�J��������R3���p��jX6AX�^Ff�C;:��䚼����C�xm &��3�4�%�4PƇax�aM�b˚4��Im��t�C.5�
b���9x�l�����i@s16Q%�x,ʞ���%�xyޢ����I��Kb`/Ze���/�`O�Oα�&X*�:sy�,�01��چߺ�Ϝ�o���]�������� ��� ���(y���2(��xq�D`j��.�jw�y��8��dӉ���r9��yrx��8��G�]�َ�p�9<p���+$�$�@�,� cΎ%����i'N �
 �0�t+��Սl&��iO�8��&�����\ml�o[���T�8��a�o��� ��/(�x�_�K��wb|_>�����9���+�'�K��� ��֝A���I�x𑇼��'��Uc+J���$��!I�\�T��U└�b{�mN{�}yV���͑�f=��C^4�� ӹE�;��A��r�e�1�[8���@�����8�I$t��%�>=�]�#;E0� J]�Z]z�/_׃�=?�N�S�����N�����)����x����.�/��VLN:�M&�zB������h�9���gs����K�O�0,��so͔]
�������	�H��rq����?/�Zxq̮�a�ۙ�P��1+�^����	���a�&�=��<\XU���#�w���ډ�f�\��T~�4���������7X��F"�����W�B\�� ��パ�p�m�}����u��q�e���˪I�W�k`+/����|MsKn\� ��|�l8�Q&w���D�l|����A���6?�=-���ɭ����A	;�J�A�u9xJ���x�>�h���p��a�-��$�z�y���<!���_��K�0^�#%��޸���h<��g����{�§�hpsl�;�e�LQ�d�8�j��u0�B�>[�w�:*I�/���{��b9Սu���I4T��ZhrQ�U�'l�9-o�t���tI���Ry�OJMtQ]�\A�Ӊ��_��	I���u���2����5r���j������:������<�Ǘ�Xha��健k���-�E�..Ҭzu�@�07��K�4T��v;ۋ�K�݅Ҁ�
a���S#;Υ���T����\��o�$�i�c��R-���&�^4��|��
��3G�	y��ǥP����I���%&x����9���kw�Ɠ�C���cx�Ė�b�>oW����ˇ?{u�V�s�Q�����`{K�nEB�<��FCY'~4���CY{��9������7��o�pcwA2d�ђ"�-ɓ�φT|���T.��-V��PAp��ݒ�('�����&�����#E&풞ʠ�iǢ�p__�l�WMBc�&y��Iz��YO��םR�� L�'�_%���?����Iy%O���]���r����3�L��Uӧ�S�䠅&WmD����\�3M�f���Xa.F0��}��'���y�jP@�G��JX81�+�3}����4�|���������+�^��n��ADH�xy*��2��;?���'-��<n�.`g��v���P�x������z�n���|D;��O���gc0�[:}�(�!N��WF��g���H"���[��y[.<��w6a�B��Rf]������D��,�d��FrX1s	��`���ź�	"��S���)��������,U��G�����Y�/d��KJ��o�uų������@QBH�+��*Xv!�\��7�8��Uz�\�&H�(��}�A��>R����O�\Y�j-�r8�e>oO�;?9+��g5;�Ln��0�oտ��]��^��P[�H=���{�6z�>+�^�A�]UDt�*�8�/��W#)DW)�e�+]���%��
A�3��K)��.��Fo���Y��q	70��I�r>�����	��d������s�1�E����JDʚ_��2��ˎ'{�L�9�͡�~�YZ��"�߅��vH�x��5"�?��S��e�\cUʖ��)bnXU�.��`�R���չ����,r��;�|���%    IEND�B`�PK   ���X�T�|  �  /   images/f1ab8fe3-f826-4bea-bba4-7763291602bf.png�YyPSY����m@��\XTFа	0:bЀ
e5��	�@�D�a\�d0C"F� aT`�.a�$*;�D� YH�e���x��^��W5��ֹ��>}������.:;~�}�v��ܙ� І��{����O�h6�;�@��������s�Q ���3$��N�@�'@��� �9�7�EͥS�����π����Y�@�-����ƣ/���{��N0��	<�u�nK0Q{�8��y��-zh���g�A0/�&��{�%�V�;:�
M�/?���n�ߥ��h�4f�ݙB��N�,�B�g�}��|�}�u`Ka1:�N����7Q�g����{�-��&�}�^>(�X5ݾ9��O�1'E*��ź��i�1�2�B���ԒK��!C��>��߹K��G����>F?���شAN���B���6��K��q������_L�4��2ǲR�R�A����ii�A�m�^D����<�.�.>���Xz�$v�xZ�d�
�"l9f�ŔTڀ�$�4�⦾T:�v�,5�#��I::�� Y�GuaA��-����c�}�1��Ū��E4E��B������KR�c}�g�yzm����Ly*H�5��4��4vH}�����Χ�g���m�ߤ7�
&+ΐڒ+����H�ZwIc���T�G��L�*�P,F.��#0`���I��J%O1��&׏��٧-�΅H>�N֙lp�T="w4���s\��V,����5\z����O?�Mv���� �_^؄˂Hl��2M�T�CfG}��rN`(������uc�����f�\���.�8-�ᵒ�(p���h^���	�x4��i�5/!12^���y�n��b�\�;� Ev/��E�̹����P�~��+բH��8z�
_�ʞXD֯|�+�{��3��O�)�G1\��sԵB�X#�/��/4����<x;<�v��b���n��J���9�H���M��j����8���:<��e�*��s�K6V7'k�Ԇ�,w�;�V���N��C�Qg��h���s�_�%�Iڝ��V=�N�b#�1,��X@�Het��������]haK���S.��.�uCu:�>Z�ʳkwq=WXs� gū�hY�"�&�[�$(Қu�;Ӝf��Ē��� Fy���>��-�;���r�x�P��#��.��%qqrU��|4���N)�s-��s~����ȡ��SUvP��P�w��C�J���w/��u���wDM��`¡:}����ǀ���(ٷ%�CC��{,JL��Uʘ�<�Kl��R6�m�x�Shl����5V��.�m�O:��f��i���gPU��U����˩�匝r5��%�'=/	9R�4��:{S��]pV? �񕤃��>���,PQ����#o@����~ ��yT�Z3Ev������=3s���	�-�[�0O�7E�������~�Pƻ��7T#����o��jd���}��W�d�\^`>/ī����3}���:1�Օ�`�sQdhN�0����l�u� z�Ý��z���b'�)K�lcș{�ͻ�#ws��7l�m?0�r �ݸ�ξkC.��d���/K��M��D�ґk���ԯ��o@���Z3���:�k^��J�_TZ�D�@��C��jiE��6Qf��,�`�b�Hw��O 9LB�ă␨�y���S_XF�l�Km\�tԌE����:�r9���һzyM�N՝Pu~��<t�<=�1x:����e.V�X_�6�̖`e�g�-��do�e���J�B������<#�Id��U��ٛ�d#&Z9:��Ӭ𥧧��"!S����P�E�k�~=Gtɵ�\R��5.9F�h�˛���JGK�o�Ɣ�1?�,Qe���g����o>���ޮ�h��s��`��6d�j�d�L��=�Swt)�R%Gx1�k_S��?:#b�j��#�J/H��ٞ$�/��xtqKKc��1�s|}	���)���ɾ���*�S��[���|�.�<R��y��N_�9?�(g/J�E�
�����5��,'"f�Ci�rJ��v9N�D���b�rd���ʶ��G�twJo�$n�2�eᝧH�7�1��]�Hz��whʋ���#�ָؚ!�CQ��_�'J��.i�U���#/�b[h���c �����#KQ\����|'�6�Iy{Z�~Ь���ݝ���=�AM:dX���?�Y�����m05�����,�������M��+rI8�:���;��V��0Jxj~�i#�z0�/B��o�����#�� ﺛ �y��k�Tr8;%�����\9�;ZJ��>�P2��ޥӻ���2C�ya���rϓ�l#t�.�����I~��yt�e��E�C�ݼ+.����Ւcf��03@���NT)����R	�^��Q�в��O��)2}2_Sʊ��cb7��Oޫ
J��+�M3�}{�v^�����]9y��mK#ca�Z���]�.�W���՝��q����6?b��KgA`���&��Y�Վ
��#���>뽿X�JFey�c��!��Ex��/^��j����.���K#����E��Z:�B�������IV1�ΐ���˹���Y�3���΁c���E) `�МO[�ʿ�˺y�c�Bb���=�9H8���u*�����?�yG��Đ��O����f>�J������N�u�rGmtȧ�CE�X�:U�F��%�Z-�[O_���Io{��47 �U�Ћ�ƣ�G���m���gj.W߹r�* ��$gƃ]��k���w�^Rqvng&��4���ͩnW�C��}=1�݉�х��|������z�;n��+Y/W�^G~�˝�vu��Q#2�Aز0d�	w1ֵ\�h�h(4�V�7�k����/e�տy����G��h"j%5|�TP`���$�vg�p�3��|�~�`�!�Ym!*n����]�	����g�%�@�EV2��S��?uUc[w���@�Nf��!�n���r�ӱF�N��N�y�w֟�Sޤc��!?�0���Ȓ,P�sQ*W9:��@���&��[��U&�!��msSx�z|q�A@��yW�ٸ3�o���cБR�UtіU?/zfZ�[k��Ý�V��ci{�����ۊ�}W�~܍7\=�7k�P����C��Ĕ�;��t�%XX$�8���:T�dj=|�T��?�Q�cp���6{e�k�w9 �U��ftQI_w.Bf<`1���LU��d�r:V?ܪ*W����Q�,�42��\�������Ks���������>э �
 ��L��k���zVì��x��<�h"
�˛�	�|]\�1�&�&l������o�З[P>�:��Ѥ�_@m����߳|4�޽�����!�����p��o���Ft}��bi<@�p}�� �p�j�b��<�5�U@��kp�����k��;Ԃ�ʋu�F/6y�{����|�����V�����L�Kf=�����6*O`��w�(.6$�/�j���z5�.��ĭH2--��g�L��e���TY��T��!���ٜ�j0����ǚ�ҙ.%�s���p���c��A8�~���=��-݃���^�7��?�T�-��^��hmt5����ۉ"_S��"�ђ�v[z;�����ƗW�/2���&�pj6�'�o��7eo~++ʼp��/(P��뎦���G�diJq�	��J���Iۯ�3@�
CQ��T��SyH�&[5R��E1��'�[y���Go�q�e�Pa﫞����e�a�!L0w�~w�%����}��	֎U^�R�O����-M����u4L�'����p�ل��M4���>r�E� j�/�5|��6ދkQ--=\=�Rѹ����u�M}�G7���a� ���8�,eAll?�[���Q��͗��᝚�]QN4�n�Z���j��zտs�L/@4-�5x4/�-l�sm㾬����]��S~�Ŷ�C�`�}(�����W�M6�M^f�x����J�ie�P���8A���[oW6�E�cKg����13�tIkŅ�+��X�_q=�� �c�u�S̳W�'y�vU&��_2׷��L��8��]A��"�S8S�z�{wa�t�2��g���<F:Ȝ�" fQ�/	pM����Tb��~lK���eb����˺D���/�q"W�����=<�ԍP�Q ���3ן6�f�dR7��*��0xAQ�c��q�8�+$n�3��!T��m�{��I9�����?���t$��M ��8��:�&��n|T_���/�5G�#��#�_��������,\V��Q��ȳ�W��d,Gù�����Y���G�'4f�b_����K�uܚ?�-�3��8���0kj��{d,Ȋv\�f=��ar�ǻs�,��E�^��9h�^[���J��,��8a�򇍒1u�'��-&�RK�8m��u�U�f� !��-�eY�Q�<Kܛ�����
{�i�{��53�zܖuG�ߟ3E�P�0�[_h�W�6�LZ�l f���(�����H�!����IJh�QJ���K����
�]���+ksfR�6�ג��F4)��r��z����z���<�^6�Я���k����C��!��4Ź2˙��֯d�Z:��{�x��%̷5V3w�vb"��D�����]G��o����s��$�H�q�$�����?$J�7���µ����רy<�;O̪7T���A�w�O�'�O�z���#�{$�9�LY5!�o����g��B8�(�T[����q�bz��;}�F�!���Ĕ�C�K�7ܽtWn�)�2�n�p~�=���t�`[c6�]d�Qi�)�Gu<���v�+ec���1(��2+���yܬ6�
��{	\j���
�/�3�gV�XM}��WJ����V7Cv�o�����H����<:�������qŗ�=��i�P����ı��X��D)�����FW�ھ,z�s����_�x`�gE^�;i"��r��n�k�&>����]�Ƚ���h����@���/�7�u�v�g�R3[>D{w�k�(i��(}5>+�q��'�R���~�7���̊��[�B�PZ98.,���ɢ��/����`��qY$�/� jPT��,�͛��FJ�ࠂҬ��\䂋>"�K��5������hi��4�Į.�("�aM��^^*���ϱ��ʂ ݉�m���n��Kl�e����uHzHTx������]|`��uR�Ĝ֥y醤Tu�X%@9.F�:�+��Xs�KȜ���{��	���92!��a_��35g;Z0b�ܬ/��i���*C�6V�+<I���e�����ߜ�����1AwLfF1�?��´�$��Ձ�9��Mk�"��C oXK|>�n@��l�I5`S�����Ic���T��hꩨ��`Q��I�4)u��_�I
o��j�L�,�x��[�$c���i>���Km��\~L� :��QS�f����i��X q��'��k���	��o��n��NR��5��f���_�e��Z��n^U����ҋ$}��Z�Y�2�'�]X`�(٪튖�n�{	�c��>�"ŝ��f���(���K?*M�	���=��G6�=\�t�٘4B5����M7�{�~�F���ա�{��VG�z�n�&[���Qcl}���'�/�I�4��'���$g3QĴ��B-�u�!�i���G�~�q^�&�%��S�Su���K$Ɯj�54.��������߂a�or�����OX��8�4���?��8A�em�o�C�~1��������ȟ�ϔ�x��PK   ���XF���?� Q� /   images/f590943e-678c-44eb-a174-3243ba5f3820.pngl|	<Tk���ܴ*�})�F)�2�t�d�2�L������'�m�si,Y��kBc�Pѐe�C��4&��4���ֽ��}���u�s��[����9�~�і��!��sdS%"�^��I�J�<��}���z�߽�7���7x��BC ����V5:_6(�ex����������__�C�n(��u�C�w�Rg�d!��c�?/��}Ƥ�X�P�#�}�`bVO-NX>��)��l��T�z?Jo���c�!P����[zl����e�Kyĥ��j�������v(~9�9�D�FWo5�`�~NA�L�L�4�M���-;:�6RT��!f�Y� "��!ɱ�����?�snRr�D��n:��8���0Y�T�Ip��Ҝ�Q�A�-f.u<��}��Ha9�:�C#J?~��X��s&�D�W��t|�ljt�X�g���x<�K_�C�LV�},�2�����Yw�揹ճ�<	WF�x��C4[K�9�p��8�愝���c������4r�3�v�R����X����i`O���-��LȊ���G��	H������hhiu�r�ׯ_37lےlY���~�Z4d�6�I�革��)%�ͩ�Q�[MF�)�OV��n0��X3<S�/}K�M�8hD�2Ϟ��s������ ����~G
+���i�j�[ZZ�c�cta���{ZJ֡.�����m��cɵG?�Zpm���k�����9ׯ>q��U�X�Y�P���Y����_P5��a*���z�$LT偽��;4Hè�<H�(�?�t2��s��;f�9w�O!U7��b�+]�){1K� ��"[]�c�d�z�0Oa�[����s�>���2(�|�z��[�?�����
K�9n���&�J�����Q:���rrrF�
�^�0y���ݾ��P�8�is/3���CE\b�m�7��'���%젡A�֝��)n�;o$�)Y�?cd4�����ǲ�W���4�+���H�V8J�&55�iek��	-iӥ��PW��*��CCz~�G_7Źn�s�_w��G�m��ϋ~�U�dkih�KjC�]1� ̈W��0�펻�Mx��������$M���-L���{�����u�B>�~�Z��"T�>11�+�������В��8���B����l�C�:4���y�;�W�$#<�$�����S�z~�"2i>5v���Є����� =���h�[߄ɓQ(��	�o}��*Q�=�9�"�V���� �*�6�^�V��k����:LY�Pc31�qP,�«�gZ�����V�vЈ��$�1؂�|�]4z�`'�mB�w�F=��[vo��0�����\�����@������m�W����ю�g|S���q��f?��p��5 3C�_��+�'�R�?���Y�S����GLE�����	Ӡw��qa�d..�\�z;�m�:==m�����4)g*�*1�d�a��������'�-F\�	[����;����k����!�,l|t��b^�z�����*��+[w�ҕ��Slg����	c���or����Z�$�*
��@�����mq��jPG��5 ������K��}��v��q�X�=a7Ƀ���g���C�>k�Mi[������z���$���wk�Υ䌔�|�����Q��w���9S�z
79�8W��7�<����ٗ�fh7kM���0��X�>���3҂�<�B)��֋ZK��uF>&�<�2-hjjZ�|��T����-�2���!�xF���K4즕O8:&|Yp���S�{j�2���t�J�0�'���5�ZwX>��_�/P��3;t7��co�ȉ�Ŝ1��C#T��I��N-����k(�KR�
�:y�q��9�N!�.?���s� ��j��L�b9��&����?b���*d�C4�ew�nU`$aAE�x�n��2e�J4%!�d�.������8	�MCVBP�!���f�U��#�g)�s�]: ��������chu�u�(#X�R�h��M	�%�Ȭ��HE���J�٤<�,�#��B(Uc�̗mo�r!(��	�'�s��I���`��BBQ�K�[GS�dՍ�
(�C�ְ�n��m�n;4�JZ���|٢��i�]V"�':��-�����|K�s@��'��` ٿ�A�k
��~��^
+[RJ*���c� ks�vxpQL�� ����&��4"��Lb�%���	��w�`��i�r��
��"S����-hw�5
��B� �x��՘�b薞��;�(_8�\z��z7 �\����u];#�U#�ΊYY���Oꅄ]�������N�n�.]�!k�ϤZY3�@X��ϰ*9�	���Z9%wd-��m�C[;�Vi	��gR9��YX��1AŘr2�k����I�e�oL�c�c X�� �$��I�-Q��3��`8	YP�UsA��O/o�)hn��]����H��y�H*沠���G�F�'�b�U�<HýN��z�{y�ʕ�/kk���.U�iC��N�e���lmm�}H:L�W�jF����I��u|�OB�*�%g	\N�m��vL�e�Ӷ��I�A�4�����_L/C�I�h�9F���*56�!�UyO,Uc�P�r&MQ�e��5��s�TM�AAW����w�+=�ב�5�I�>UNva���v���������%:2ק;t�$1yX��w'�7��9dڥ������,��ij���dV��?�*Q�B���`�3~#�	�/�#I5AE=.#�}�W!f'a�9���Y����~w�"(_K���Q��
�
햘��2{ s�M-x�.X���%R�NN`Q��,�Ȭ���%�K�U�xʣ{����o�?|�y���Y���Xe��ή���a�3�P�|:)_�T�8:�<�����%VUa�����ci�������ɒ^��ީHP.��=��WJ�����,w�()��
HWu�c�&d�=Z�ܢ��V���~�
g�HR�����J�u(���5����#Y�*��V����g�����h-�4�͛7�C�x��m��w
����^����~��Et�̉�A�P𷾒�T��״��)~ޚ~�7ԃף�W΂��HU�����\`�ϸ�Z�s:��Y4]p��H���q�o			�Qw���q�� د�`u���O~d��2���hJ}�x_x��V*��xcE�O� m-����f��1��\z�[�a���5~���q��
�~���7W��i͚#?���t[�74|q�ҴO�~--U��~�t@Q�5�5J�^�Ч�%���A�Z\Π2�[l0Ӫ���d�_��ͥ[T?/{�CXy��d:>U�-	l�"[)w�#�Ȕ�4\&�Zv��GJ��>ё�Z94�7�ݯhJ3���$O���m꟡�K�$�Q_��Rą&$�R�U;�$vu*���Sæ�g\,������,G�.����ڵ1�S��T-��K��j�#\�����]-�E?�E��a8��C��N�[1�ND&k��M�R-���ʺ^1� R�\)������oʂF  �W�1Z�����Q쨿i�P N3�S8%a*��L�f_r~V�b�+��^��G�PO[ͬ�W�k^�0��:{�R�^�?�iW��,���&�ciG0h���2N%|K���h4���{>4�Җt��C  �L�u�uu{<p�@1H\�U���_7�V�������A���w #��z�Rw��T�KR,έ3s|f�!I�_ܓO	��֥D�$YY3������41�}��OCכV���I"�a8# �G@���,�~]�:�<Y�f��ے|H��R��a.�Ӽ������TA����MK�u"9i���	CD�W��~>e���_v:�v)4�4"�'%x���CG<[E��������圲�m�»K�=���#�$ǥ`n�?�P�O��K��m���Zch��m�̅}�����U1O�"����8���.�X��/s�>����&���50R���V�ڏI�pR�&�Ӯ�y�Zk|��#U��I!�^x�f�pEo��"�!��P��@�f"ml�&�v�릓"�%��"����JZfv+�AO� ���2�a5^-W�K�C	bѝ'���.����Z�r��/ՏرI�u��&��/Țī�d��s��< x�B~�����I=j��dA#0$����Ǥ���P�)�X3���Q�����i�z��?(�u�9M΀ѩ�@M���j�#!��-��G&�dD��5S!U��s��C�$t̘�i�Q��w�_�����1W2 ��\�V@�3�f鹱R����)A���;���p�L~d��(?��%�Չ����G�6���-���p���sI � IKծ��)�U�a�j�T�{�ek� ��Y�_;t�M�Z�L���i���e3	)]A/�;|��?�P��ى��{2�H����h�n�D�00QK�Lm&w�=��� 2�~N�Z������yMj� ���٢��AX��3�OcY��G��~�F�k6=��k��-E�U1��1�맽�ۀ�ݿ��OSu�A��P����U����IU����s9@y�[X`���۩�`�Iy�x�.���=.�\gu�,u�oo7�7��=H���Q9)��p�jh�XR������)	�(�j��DS�i��:� ���j�㳚��Z�Qů�+���n}{�8顰h�}o�����5�Q��3N�GL.'~=O��*�����@%iFFizfP�>�~ke조�g)�w�7������������r���C�?,��<�:~2f\ic��+fچD��#����m��H69ZQ�Hf���}��5��G���OH#G��g���%�H�U]��SIQn��C&�pg ��D��Y��{-�~�a-��䍞�'!3@N��4 '��%���_�jN�j���D�e�_���Am�z{��LBաm<A�l>��~���w��"*=�v������QU�$2�(��cƟ�u���wg�bT��ӧ�����1�9������ 0I>�����ם���������6������3��ez��G[,����ݛ�x����q�׾(�U�[�ܡg��?M),�*�7���L�q>�c|��N���j��@ ������㒒�'%?�H|VX\�:=�2)���Jm��>��=c�w���G�4Z%�w��'�(���F��6X��M�θE=��3�M�E�ȯ�=���j��e�V�1jpn����8^��a"�Ls`7M��Z�#y��?;�~ÚS��`���*�� ._+�R��PL#�yY���JJ�~�c�����csW}�6:�� �]�*���B�Aw�E?}�o�� �Z_\W��q$�w�B�˹��n�F�Q���a
]�����։�F����WQv�9�HU�������/UT�u�LN��C�9W��%��\5_��TSY��>�/�� `^��5�wSԞ-�_�W�%Ri�vĴK���7��P�=������4�J��zr��c�E�ȇ�_ذ�/,������&D|r����^U����o�t-�-�)Y���u-�w�s[�Aީ�`�㼈Gx��م\�;f�\�3��L������ٷ���?�1��ia��y禕�0��
@�pn����Yl@��&Oyvzr�ZDV�#R��f�*��1�w���j�!r�"W+q(:A���eV@Qk-�[������.�u���$�7m4���_�1݁"�P����y�a�Zdem�7I���n�³)Z��2���4_e
	�sN�m�^�.�CjjCW�nm��+�}�h5��N�j[���凢���	a���ǫ,m���K�� ��IG�y�J c�4^E�T��ӪV{_8/�H�7:�Ǡ�<��᰷�#孩\]y��4jd7f[KI^������=ԡk�g:V������s��R��{�,�D�c�����g4�n�X�k�,B��DI�[1��,h�����D�T�נZ�2%����9��*q�N띌a�
��?��j�nYP�q�h`(3SD�"`�w,,N� QX��{��1A{(��G/m��c�xUPv	MMM����}ʇ�˟J�̎�qJ�e�`w5�p�T)��~�8����[��)��I��h��
��AӮ������[bק_���į7m�d����nN��Ҏ��tƑ�4?��'(���oOÌ����$�i^�V;Zf�>?br�'o��gB�3��'� +�]����K0)+%z황*��*Uc�$�2��i��]�I��,Ѵ#����V��F�����SD`�t5�i���ԡΌ9c�#�7�幖A��QOTtƙ�5NQ�J�9si �ʀy��Th� x9����t�aGQUj�Y���/�:H��� Ĥ|W!4"�TUᥛ��z�e���?�!!�E����30{5W���Si-=n`�ۥ3F�����9QF�{���� �8�NK�>Vk�y����ㇺ0�-ӭ~�bG�$ �:dr�4'� w�m-u����G���4\wg�8����y���>k��x�3�ǃ�@�Ք��q�w�rA��T0~Vt�Qg���6G���(��O�U�����y0!�6�ݧ��e�^�^�2)o~�U��Zм5�4Z����V�����$>:��4V
(��1)� I�H�#L�`��E�Ӈ�ڀ����^�`^aVgU_�OW�*�Jޯ�D�F"��OSo�R�[�Ј�=�v��%|�|��Vh��މ�͖5���¿"o��_$��Q���o�v��!Z7�H��S�/�h�C���G���ju�s<I6;���w�|o?iv���u��T�<m^��_ ,�\�W��f����o��"0�b$g�����6�boP4^+�Zsb�W�^��_� �?�.U��W|n~]ON��?�"&�5��j���<P�����"���K
��,<j��� �(E�aFL����yj�� ��a�C�U�s��x����M���5=3nۈDv�AЖQ��|���K�9�k5��wh!i�z\lu�v:��ȕ��Y?��l,�E��rk��w�1c<�p�T%�@\�&.���J���Ʒ��!=B��^�>=	y��42H_�[���A=���������&�
�Ne�������=��M�.�at�J�+�����q�1�w ��M�� ��y(ߢ�5iJ��М,����p��.�H�	�eC#���	n���,�W����a_8#-,�?\�-�!��U^�o�(��tȄl�������6|�I:�Z�{�b~ާ�-�`���>)CA��~I@�LB��D�������g�d�;v�lK�X���l)b�Ԥ��+`h��A~��$Ŗ����ر>�H E�
��6�8hć��.���0���ݘN�d�Ii�ޥ�cV���U�F�����K�c���E���H�M�m��a�_�}3�۰0(.�C��!�m+��!��X�v����ج�}܈_?�_��$�<���(=w��漟�E�����q�n`N�.-9a��?-�/��Z� ��3����Ɇ�.����駤 �`���U�Ӊ��*Q����%�B��-|"h``�z�h��Ќ	f�x�i�\��ޭ
����ڻ�g�c3��R�L1ݖCKZ��U=.
@�ې�Z�����A��Bb��+|�C���C�KK$
G:��h7�׷x�b0����@�i�nz�v�a[��c��?(��-S �%��(�<! y�$���A�!�����),����] n�~�����?��@V��e����.$���ƨ���Q�3W8`�g����κ�)���`O�Y?T��X KF�`6^˴ ?�v���.&&��+����^��g�ysz�n��Y��E@�2A���2�^��p�>��m*�qNZ�"��k���X�����j�E��5�OYw��U���<��@�M��f�F��Jĕ�5i�f��Cp�-�N!��4Qx%h[��2��V�?@�u�܊�%Qt��_:����=���ZXD���fA\¼���ʀ{�T�T�Ϡ.ֹ�C��}�TQ��ώV専?�=�#�3z�W4��
ű2X����h\��9JkVڡ(�{�Vx�ϊB�Vx�M[�(���x�k�β���e�0��Sk�����y��Yf5���L\�q����Ќ�h����b(���T��
���}�M
��g�+��B5��h8��	�;�q���(��Ո��ۥ{$Vim��3�N7�4	���< �C�!��c����	ߎy��G�OH;Y�3皥�����vwu�� ������8�������ɾ&�ed�<<���Mݴ�@64�"%��+�p�*Q�����6v�g��z���+UcyT�P���z@0��qr������)�P�|�< ����~�a%�l�]�ݟo�:V��D(wu�DK���Q��#�G�D���ߘM�	1Ka:w6��b���٤�VӔ�^K�g�n�0��}�����f3	o R��J�	 :«W^}ά���H�N����b�/raqtŷ�T�\KG'���Kt=�s���>�(�S��h^?��G�5'����@�]�^VU-}��7�~DAf[M�kmںv�g�Ry�����s�IRn�O�a�;"Ǆ���fE��| �@��s���7�&����sQx���� �Q�&�!1������ń�����%�H��Ɩ�}� x���DFY�ҵ�K�
��%��,������ͯ�|Y���\���a~~>��G|�Լ�e`�k%����d^P�*�6!�~���A��n}� ���r���$윙D�3^�n� Y��q�~A+8��#��`9فEXD�1�Pk���p�߰0��k�V;Dn���y�]9_D��x��G[�į�_8�Y@ht�++���s��H�+��yo���k���b2e��.�H���D)9��
��g�����!x��a�-��W! �H;�N�Cn5.�^"g��v�4�A��T�R�lm,�S��ݭo&��s�;��B)+�i1��ouEM�J8�ѿ�c�# �]����p�����cW�����u�"��7%�μ?`2s)�L>�*��=�������R k��ja���� ���{XLLX:}b"����ػʄ����9����ukd6�s�Fgܩ�H����u��/.=w<������������m�H�y�<�wU�OU�>���Xw��B�d����ŽO�*�nҭJ�9[�=����d����O_�'��\O���R���|B���"���=䪄Cn�H�L:�ʈ�v��ѣ�j���B�y�o�(i��Wl���?Y욡���<G����
h�c��Z���I��֦8���@���gzC��u�q j5�Nw�����o��Vhp�O�=�
�D�0�t�hĖo��t'n5A��^�3�)ƙ�Y�[�!����F�oO�tp��@��Y���{����}�^�J��T�s�f��A�w�F>)�
��%ԩx����^�u�����-QWlzKo60x1��\�DL,���ϻ򿳃vӐ�� V�IyWgq[di�e�?�a&zyU��mbJB�)`_i����H�O��tǅ�Һ�w����2ib�X?Xj��!{��U�W�%7�<OG�p�Ϛ�e<qMo &_X^\x��5;��O>b��0����/��m��d��'6�1#'�Y�|!��	��3!�����C�f͎��@���Oޮ��D�{�{! 6+���Kx��o��oh�ZJ6���N���6��~{�L�DV2��)�b�l���tU�����9 ���e���U���.��Pl��'�*���"�'77��V�b���_����m�	��Ժ��!A�l�"���@�7��v�wU��-�?���D�|�	����uğ��f�nB3��Kz���<N��2�f=�i��p	2��B�$��)�б�k�Tp�꟝��ֈ�����s�۫�ܤ�H��,�X�����:���]�����.ܳ��
�����"Z@�9R[^� *f�!ݹYSV�����w�?yb��z�7�wr�Ԑ��>��Gn	=�q���G��o�����>ee���+�M(Ģ�	u�H�_az/�ZG�����2�0}�\�B٧<�!��-��o{���qX�*�h�#_\�q��Rz�3�n7&7���>�+�d�
���;`���W���ߒ��-Y'�|Qػ?�o��_�g�����`M������He]݊����1H<����_bQ��ɒXe�z�:1�^�dg0�V���P��<��}L^T}s��u_�3��Fd����4s:����6JO�v��[OZ1�W&Of�Y[��{���F���~M���m8� � ���f�G�[���ɣ!�aa�nn�Z��jm�1������Cۚx�:͉O�ɛ����G�wj�;���8^�B���b��6��s��f}'�3��b:�(��LU�K>���c�x��)ͻ>wvP*�O�Lh-�~�������P& ��2nFUuJ���ʽ�9�i���ʐ<��Zf6����p��^� ���Y;�h����҈A��l�r���1զ/&i�6��6�?��8Nڠ�}���˩qW�]��J�<H�间{��ɣ��N(|���>���E�ޣ~�?:��;x���o��gk�x��vŌ|��͋.�ة��h��)mFɳ蝯���B����������7^�kK��:S�֪(�2���ܪ�|9���Mi/��?����]tyE��0��2�/e�����M��[_\��{aq������I�z��/�."v�#g�|��\Z��)�+{��ߡ{f��\��q�S��+͉�x��ZS��p����Y7#�r�.���D��� C[^43��_1�ƍ0�����7��iڀ����A�<Ԑ~�r�����ϗ@�AΈF��U�ѩED�z?М0nN. w�{ﮘ��j~��d���s-�*/�H���z�ޡ��ba�_��^��G`K�T-�B����dr)�|�X%d���T��?����3��]V�m�::1팤9����P1��;V
'Q���l7.V��	E뷓0I��Nv�}�sA��ެ3ˣU�O_5N��c�m���[g��=��˷܈��p1�ysr��_��|K��桋(�� ]>{�=������{T���ZE��E�h["�P���wȴ�P�Β>�C|
���5m�=����>5��n�/����Ϊ:�q�m�ʠ��dM.5'�J;�ǧ��y��E�=��_��{��,h�����̢��<i`{R^�.ñ^���f��X\PP��ݡ�]D��Z�V���f��}���v����^56f���.o�mT|t���{m�њR.xqN����}����t(�YV4�,f�C�4���ȇWRUu/M ��| qd��o��cR���icVAL�]�O�8|B�J�6�U�ɲu���\� ����vt��{���_�}>�O�D�G��ʵ��UF���?	���ڡ��-�МwW��D!�������'�1?:�d&��hZ���l&�kw�(�@����=����"ö(�݃��J��9��n	m���G8������S�\�瞙���seu���t�p$O���;m� ��]zܑ�������v�Z��d
�ޭ���-��$�m���0ϏD!�m����	�
_KKˑ}�rO>d�>v�s��٪ sOK^5z97q8Z3�0�"Rg���m�(�x��#�z����	;��_���6�T��Y�t��c��[�&�#�O}�7_RϿ�� ����rƚGI��m]r�m�$K�8���F���N�������"��`�	���cEG��!�5g�l4����O���,D֟(��'\A�Ū��h��,��k,�J&	r�ǎ��� )�&�_��$�\�w�9��t��g���2�˷da1KV�f(�����b�)�姞�#`*���H�e(�����W�>��?�#EG���������5.g]���zR�y���{�G�vV5�7�hX/�s�(�����kH���wke='�<�-�-C�`NH��V���o��O�w�ӌ�7��Q�\.�V�1�KK�k:�!d$� ��F��E�v��[�+r��M/����r���C�{�9�v5������n���%Χ�����L�w�{�����-��l�� �H4�@e��TW.�Y˔�:n>�����t���OٗKBC�Șb���%�t��UU:CCC���Jw�]f8ѪW��η�2'��A��2�Zz^��+�Q�CHB�mY�qѵ�U�f����7#e����i��?����0����V���1��T���OF�77�q�N� #Q�������z4znPlvP���?�z�CAJ�?2�c[8��u^�w�$Eu��������$;�j�:���hek�]��A�F8)��L��&��.f0Y�O�7Lo�1�"W)��-'��+�X��n��7��W��:9��l�v�l�{7����8�ʙ��Znl_ac;������⏒����0�G����,(�	��G,��g=�w1�(�@�`_� �A��wI��������sA��P�H62
���'L>�j��1� F}�Z+��F|���4�9�\��K�3E��O�E��U6�s��yJ6v;�N�~���zl'�����?�EC�	�� T���lI����'��7����O�\:�{�;�� ��g*�Ouv#�	W�,bg+Fh��G�%j��.�~��v�	z=)�}�LN5�g�Dz���y��ӏ6��D�������/.��r&ޙp]t��p�-|JY��q�0~2���,j�m{��n2�,�CM�Q��}�H�oq�od���\�?�����5G�i�8i�+?�:ې8$�8��ԛ��I���j��]&w��0xB"�؝�]&(������{��&]_�p?�S�)K�M�KT3`$�Vf>�[3\ lB������0ޤso;��@�0��:�Lo�Ѩ���c&!�q���|jҋ�S���N}i���Ih�ܳ �T�	*Td����>�6'�Z�V��Z���+Y�/����O�ϢEA�K��"NH@6�ʍ�U��1� ��㩝w1>rM��B�11�?LE�j�Q|�8d�WU�:$��s�	����w�S1��g�3߾��_)K/j�+rv;��,#�K�r�D�Fl��=�9�\d���O8�C��������r� }�uO ߰J����5��c*�P�Ig�j�S�(:��2�����f�O��R0������|red������՘Z�>���MȖ2(�Wߴ�>�x�:Z;lja�{�^�����_���Tp5;H���V��\S���h���I~��/r���r ��y��\��m1<�z��p��!6�|XG��U7WegC o/��D��O�?y<!E~�״gn$�H�? G�������K���EE}�QI�/Z���8����:A-�m�������܃�욒P�Y�ʙ����:appǜW�@O�I3N���B�,���$q�5n���A.m�)�a�gy�U�)I>��ᣟ�CT5H�m|t�j��{ �D�� ������օO����'���I�+�|�ĦDa��j�?^H"f�"��s۱�/�[�J�:G�,lV��T����k�G��ÌH�^*�r���{h���'�^sɞ�Y����4��R���K<s�%��V����$I�O��٧���#��	��%
��؟;?[' lM��Ӧ?)��x[[3�	�Q�u#i:Nwj��]Cic(��a��$*���R��v����A*h�Z�&H�o�$��X5��
��_k�6��`b �I��q����3��؈�{Dܗ����E���=65���)Ȍ����*VY�՜�F2SS�����ݸYU�щ)�>��*��������U~;A�����x��������IV�Q	��U�~�OD�v�$��,V�3>A��KU 3k��d�9��k\�V�Ygxۀ�!����0v�
��� �q���r�OC�.@�� 	���$$)��َVkݮ��]2h��֋�<���E��0�#{4e�:���gᰟ�B��b�V���SƽtIK=���p���M��m�����o���r��a�M��	��Ah�x�Vt���U�͸��z3�,�B=��LE^}�h���^F�iq0� �}��"��0���Ji7���v�H�R���G���׌��F�/,��-3�'`�*s�U��Տ�u*>���)!e��`]��#��d�$����!�F;)}�H	`�!d�*x̠����^��	�ʲ"X����i�jR��/�x�r�����F����=������l�x�A�<uӕ���#MӮ�s�UG���� u��%/(���I��6��T�ͣ��)FF�у��c~z�X=A�>p?�����K�1vg^���N|��]�@�)Ƃ�hl w�R�{���
<���0�y��ۍ����&��n�<�����f����3\؏�����mVe?�n�#,���ī��^�pخ��,^-P���e�oW	��.*�|���T�� ؖ��t�o� 0pb�����3B�2�W!Ig�HC�����D���' ����8�7g�}f]��n�%]��{�"�@�q��� ��7��u�8�Zj������FJ�'ϢY1��*C�n�����nK��Huτ���;y��=�MOѡb����h������}]PR.x����&�GD�\u��d��P?r�Z?��7��;y�4YY��RX���K�BpbŖ��v},=���n��$-�w�A�֧����رM�-t���i"������Ǘ����n��G�)+.�p�������{?����ɵ@W`��\Z{B�{�q1��<��������`���<� R� �V�Q?Bʨm���$���=���ksH�ݬ�����Y�(�Q@�u�Ƈj��{-�tH�Ů��`̈́�E�sJ���ᴹ����h�sJ�;���ww�`W�u�]�X<�'E�r�������0�����{�pa�4�يk�O�X��!����n�PJL
����!�9Gp?1b�[/�v�G�w�n��OF�"8��e#���r�X��7���3��l�a���>�����s�AwRr��t��q??��}.�\i��ܛG8D�}��?�C�j�n���Ir�3��m�����귋�+�f��*]�D w"1d$����U�'p?��P��j�Jg�α�5��H��c��x=���"�ݞ�08�^;�p����v�}E�Z�Jt�K�V/�ra�3�s�@<�A�1�����[�%K���2�@.s%�+Պq���,$/���i�}�ȞE�?5~f!�^sa�׈�I��2�G���� IS�FW0W|1���_��NHM����6�`����)���o�����'YD����\���x�>��T��T�D��=+ۑ�i)9��^ٺ��D�p^c���e�Z�� ��9�KBl���b��l���zf��{��'@����o�}1s���a������s�:bu�<.��MB!�M��!3 �lz������"rb���Бs��ˮ�l�j�&P��_7HKNwIJ&]Zæ6�����_��L��gU��*��3�d�f�Ւ,�����W��+�.�g�	���ql'��4�����RX�3�.�z`�~�A4xk��{;�%� �{�����vB������V�{�g|j�.�����
�w+��9B��OE��/���V��!�_T�q�b�?��>#�ȉ9Yy��A_��͖�EK�Y���L�l�#H^�<I'2�Qt+=���򺺈�b�]�(GEy&0��z�ex����k�.�*`4�j��3�'�c���>����h�:(8%g$9g*�F�,�s��-����{�l�m)m"��x��M�9*5(�r�T1X�����S�{��0��8����D������g�ȭ:��� x��e��Z��0���@��>][�wh����ȴL���ؔ�c�G�	l�$�pTOD]WOk��Q�5�{�=�R�*n_/�6X�V}��"�����}��x�<�s7���_O�bg��E��+��$��	���k(TP��^%�Y�T��P�����y����e�oא;;e���(Z����~���
�8=Ӯz��P%�����Ɖ���!����N޿~Rb�<{�`j�?�k�.%b��f�����2V���7��O��"�p9��EkOo�:El��pN{�d_���G�.�'���rk�4�a�9�+�����Kb}�n���DÚ�:�C��"}��DȪ��S��O���o���>�쯥9@��ٶ�ހ������Zu��$!�m5/�ϐ��O20;���iɾ{ܣ$����G��lv�GrGeUy�6�J�P=�q�r������Hv7�<|J����n^��R��	1��K�ĖR��f�5��Y�=�e��'�x�E	��{ɷb+�o��H��I�TY����.����߈�\J���Y�b!��ҀOt4�����M́�s�ǹ��dw�r{����"�I�iչ����;>+�z��+8��eH�|�Qא�6<ᢑ�asx�����N�NuO�~�"_������)�ҧXL&��W�m&����	ϋ&5�Oq�C��j���.�w1�-��/=qX��}���6����~��e��ߟcW����' �n�sE� ���}�o?�o?�4z=�B.,��ƣ�Ӽ8c*��?-�?�B�����!F�xD{R�(EHZ8	��1�c�lz��{P�O�4�#������4���}x��т��?�s����Z�8�c�So���r/�0�wXW�Q�T��Ru��*i8n���{40Rk�x��_�*��U��_�]�K�:����LP��e�3��m2sɮ�:>
��S���8�H����͐�]#�`R@� �C���=�v��^��~��R
�>�������^
2�1�jv��Y���4�:?�XE+�/���`ȃ�מ(�����>�A�_ >9����z&$���>�%	��n:J��8dP������=��'��S]8띛{������oG8��- �D�4h����N��E�5��7��Ѝ�o��!ϙ��)�`���ڪ6�A��*��1/]�/	�
�~[�K|����N�$q�*XbG���4��C{5�)*��R�E~�W/��I��'�<� ٞ���0	ջ�m�����5P��Sg�)�Z%����o�:,�5%1�7X��9�q����/x�!��r��sw>�5� �@� ���z�Bdf R�[-A����X��ׁS0��%:�rg%]�����9���-��U������ "��Fq㈏�ذ\Ҩ��<bټ��sy= �3bI�pU���C�*]xy>�A]����?��w�15�P^��fWK��/ަ%�`tE��!r�Ԅ%?s|�t�H7�h�11�=,�H�� [m����/����L`T�"��uK����/��>�KZ.9E��Y���2�i�u��}��D�:�v�w�=2� u�p���E�\��PXY�w��}�x���v#��<�-����6~8��!��H` �EYJ��,�$�Q

��/�l�P��
)棨��<��$n��Cey1=�ZLX��V��ˇ��8�jNe}6�b�� �uO,���r'� �8�D�~�)���xT77������x�A	���t�e��4q��x�Z\��<pt���z�\�i�:���������k�#�o�U%�GN��K�7B\/��
`��?����=�8�h^O��?҄Q�9z=F�"#�g�Q���������z�x(���V��$�t�5��)��-�9H��4*5�Ց������SMm�Q-������X���z]w����������~]���z]���tZ.�M0��g�۫�� ����E"����Т�AġFպ�u��6��{��sH�]��F����+��p��L�<:r~m~>������䤢}�¬�����7#��;�e<V�>��hD���:�	r#���8Ht'�$��x��!�t������o�ʕOJH\��mE3�{{S&�ƍ��L�]҈�d����-hq�t��^��{�_�-7?,,�g�]�4$�VP(IwQS�[�+�>�]�k�nb)}���/~.&]�K& �/�l�f�~�r#c�^���@>Xr��it����g�4�3\��M'�xH��P����l�����_�1^~w����*�mF+{��\�@N.b���]5v����V@9�M����#
9�GR$����fD���a��4Ĝ��Gg�?��x�c^4r��%��@A&��a�i᠄�X]�88	�p�Lc�<Q��b	pi
��U�oe��������{y�OJw]D�C fk��zm�Z�>����A�]��}��g�:A1w��Ee����^6B��I�����8���ؿ*YZ����`����E�0Jg��L���J�'0-��ʭ
�-�n-����Ȭq�ԟm7k�cN��u�$�KQ�
W�j��|(+��*�nLw������cb���q��Qp
�3ޮ�Mӎ�ɩ��Fc����������`�S~w���m<~G�n0��,�B!/���ȔLː{\��Dt�q_�%���T7^�<�:Er�	v4����l�	eq~�ʇ�����K�D�,y�,�+[�"��YO�V>�|5�\��x���N�� Ρ�y��{�v�7�i���Ga���ܵVJ�/2��F��W��u�����&�� 
�9�����B}@J�G����!���O��Oz[�/�{���9��s��X��B#�p$�*�v�x�A(
�w֧9��I�������ޮ�Z�,H���<��]y�U!���_�ap�{��b�=�B��֞��a�aM�Z~��i��O����r��6R���E+��K/L�xkoQ{V�a�%b�k3���C���9��|�i�ŝ��Y�hX����N��W>�J���V�t���U���YQ��l��QW��vZx�˹����j�Q��D��)���6����S���vn���Lqbr��������k?��Me@��'Nm�'����R?�v}�_a�W�d��[n���:���	'=���=������U��^g��8�bU�8A�(�ȿ�0��.�WK�ޠWz�_\��v��>�YW�X"�Ѩ������L~�"�J��p-��)�d�"�!{Xc:\?s��yÐa����ǧ�6*>�5����qS-h�ڒ�B�,FW�e��������wc#.0>�<��o�W`jl,^{���%QkM?��vK�!?��H{�q����Tj�p�D�ݎ�{�M��2>��x۞f���&�ˎ����ՅNx�ۚD���$�d��IF��×|���q�R�T�Fc�{�D@cЁ��6�\�6VG��Y���q{VG�z��	s�c��h\E��r����v=�a������b?/�<t�]��-�$���g��POʝ1�ud��u\���+JGV!ҌG�O�����+��ri��z�A���&È�\he(J����Q�h8����1ΏͶ�8����W��6�!�֤�����E����im�UL��}�1Y�N�pk�~�d�ڔ�Oca3��Uh��o}��*&�ܴ��'r�Q�i{�|�ܨ���0 �G�qѕ�c���{C�Y�t���!&�Z"^k�
=�k�f����*F~*�&e3�8��D�y�d?���o��re�K���EeM;G�����,��Z�o���P�c�#h&	#�R~w4�OA� �\d��)��|ъ��+J���/uE��W�V�j�3j|I� �ױ�TL�t�i�����6��Lh��V7H�^���D�z�#a~�8O��RO�
��⅏k��],P$׭(��*ĸ�v�_Ǟe=sƑ'�\�S�>8��W�64���&�f�~�o���x�6`����~aW����o�	�r��"��p06�b��΁<6��N���Z�?�x�H ���籓tؽ�O�Kw��Vso��둗�Ak��3T�rL=h$��)����nN���m��w�����j7|�+�O��A�B���~zg�/����dJ�����BaK ��8����ӥ��	$�[_"LD��E�W!��ςcf��D�`-�i�UL���]OD���Y���9��m���\P����X�L������*�����=~�̙iCF�4�I��f���Z������:���G����Ao��U�ϫ�GMe�n"C�V7��G�_�
��PD��ƒ\�g
�pC�RqX
ڟ�hz�,��C;X8��y^��\��D��,)'YC[�Iw�����ze���S��[n政��u)��<TL?_,���2J!�z�y�� ���Ӗ.Ϻ�,�3��d�	�B��r]+.[�л/�mCB�������<���r|�L>���/��],����`=M_�.��ր������^?��ڹ�` �^2�>h&���q���P�x��g�T|�)vy>)��6$EUwU?�<8r��Ϲ��uف�����^�MYub��)Po��﷙N�o�AK����@��Ӫ�(���.l����%�/��,d���Ki��*�ǣ˙\��'�L2fY���*rҙ���T2�r���Q�t��M%5�+��H]P�Dk�'�ݽ�vJ��>���U'*WP�.����/�'�DL�Mj��)�z���w�]�d�0�X���Mqa`e�ߵ,6��w��MJ�����c����F��YW�S��E�?=��3����麌�Bk=�K�.+���wwe�UOπ�@�?��`M��Fv�4C�����^���o�����e�����6��%m)�E���d��⒔f��}L�ɍ���%	��UM�ؐ��y�y3�@ꒁoI�④r�UZ"��lAhr˔�x�]q@yD.h�@r����Яx�t�X��͏��������LL��N[W*����\he>������0�yd �!q*/9p�o`�����*ab�bBr�?V4Ϝ�M����37fZT�4̦�Ӄ�L��g�]�9��o@��)��zZ���\��R����w�y�h����v$A�x��<M%A���H�H_Wi�#<�z�n�Z��>�^ɸ�!X�'���o�jW�~}r���m��P�4-˛.͏`3��+��L��.]I��q�F��O�uІ˞]~�L�W�H�G�.&�g���Zr�zzeF�Q���ۄn�C���*�2?�<��g�Í����H�%)(�-�C�1�#��E�e8Vzd�^l�5lNo�G�J�26�h4���I԰E�
�lR�xq�Ir�^�Dnr������n�{5g/����SGn4�ZŽo[�_v÷.=8e�c��nu6�"��X���uA�A��"��f��EZze����~4yD#SoBn��wŝ#[��#�*��y�%��Hr�.A���f�\����W-Oו�`���@�9�5)@������(����~h���x�?�9<���'~�!���X�W��M��=Q~�*�=	�(�}�;)=�Y0Q!�?����~W��p�{ދ%�ֳgh�D�C�T9{��nF��Y�fZ��N�fǪX<���2��YC�=��Q̺��r�N���8�t��G�Ȫ,;�[��8�!;�QC���UO\Od�!�n��cAt5�7,���Rӂ��ZW_|�󯤴;��,l"�XiT�͝�Q��J�獮��Ωx��R�М�0"�{�F{�TŒ��qV;Y���hh��vs� ��q��N��E֔��3s�j�6��vz �٦H^�$ǆH�����W�>�X��$�����o!�W�wpQ����ug��K�ckrq��'�����zyO[��?L��r<9���7D;^�t=�5��n���d���lJ��OvͶE,���I�v�&2���U%LJK$-��I��������U��*l�/����篏k:"n ׿H�]�o�\��~e9�M�%hA
�攔��з�i�뷓b��A�qg��u	��awY���('ϔ��v�]�4��/�^C5��Yc=�ˍ��U�U��DC�5)-��B�**ý�h���O1�'�{�!c9��������,�c�)��yO@�Z�&���0�2����.�J4������NCi����Y� �-�^v��,�IvM�ӕ�c�ߐ�)�E�v�ʼ���2�'���Kʎ=�D�P6�mZ_&Z/LcK��6���vM���ZN��.�6ym��\��BV������o�}����;�ci�Ip��Y�n���+,�l��|	�z(��r��|&+������q�w�9�G>֖uس�̠�Y�)�ld��rM��Ӣ|��_��K�ݭ	#g�~�`��N�{��]������]-���{?��К�tK@�6�h�K�9O��U㲗SEO�y+!����z	J��q�R�h���O^C�d��&����c�5��M�?i�r��9�|�5?/�z6?��'�\פ(�ޏ���=�Z4�hqLJӌ;��#�Wu|<W��Co���`u!LpSy�y((u%~ԕ��Y)����" ���eM���r[\�3�B�2b��K�`��t[��`����.5����f����np�+һPD��ۧ�i+K�O�aI����!T�l�,M� h�fC�4_�S��4zWS��N�_C&a�G.o��߼$_��VwS�%��4",���0�c�LB����X�zl^Ŀ})��[�50I[���\�P���~����P&%®V|�)����;�.���;�X6Ò�n��=�����,�4n�U�O@��K�ܸf��C�h�/ٌE,�Q~l��2%��cG@����������x?�A�A�X����2��A��Wӟ����Cs�"?}���~�������H���D!��~�b���%��!u�h¬���؊�d�6�QG�v8��{��;r�d�巑��������썻�OKN^��B-���vUBv6�n���e[FD�eee��p�W���iM[aQ�-_�eQ�W�|Jb\YS���,e�?��.D��422�#��vy�$����k��^�2epy�(YƗ��-�%��\CB&�\��%�mc�;h��4�#��`2��1%���(�Df!��4tM�Y�ocW�n���|}+�U=zT��QP8����N��%,�Ϟ>�P�=Z�����ۗ��p[p���XDpx�Xz~�����΁-��>)��VU�[Uz��I:�~�GȻ�nO[1��M"c|@�"�R��疖��4vD�@�#ig����v�c�����a�E8��S'剸!�GC��MU�ZS�eK*5Ǻ�t�%��d�"0�0��3���*پ�.>]������iHK�Ӌ����u�T��!�k�!Q�j�=E��N2j�P.� 9����@�e��V�p�BL�ړ��

̚t m?�m����1Š��}>���6�.)��ǓǮ��k�y����K�R����D����0�ӛږߙښߙ[�%;VP�����7:���%���w��lVRh�ҹ��2�:qִfgZ�RYO6b�4��+���Xa[y�g��zDO׶��b���j�zudb�^("٢�����\U�;$�c�����y+�ZU���&zjs='|�𱫰K����
����;[���b�+'�������q������	Y���b�	M��??;���k����m=�+ѓ/��*�n���;n<���_�ӦD)..{��c1J��CI_P�Eq>�ۤg$]Z��l�zX�J뒉(A�7w�{Tc(����5&CH�6�m;��P.�#W�M5���/3KG��|�e�a4-���1�P�rZ��K�!���a�����'��"/@��Fr��;*e=�R%�����Ȫ�)J�sl�.�)�ƾ��h8]����k _r��8��yJӗ��W1���q�vR�Ga�5j����Au[I�yפw�q#���`�t:籆|��$�IŻ��|���sy��'���JK�:KL���ƙ��P%a��*H�=�4-�D�DJ�����ճa���5� ��5�Im�G��
�lQY�W�|Ϭ�i]����G���h<*�7����{4ȫ�,��[l��}7�0x������Y��4ׯ��p:��+~�pě��:Фc`�Ԡ�iP�������[�����z���f3~o;�V�$8Mao,��iA�D�ܦ6��Є���e4�ee�I_�%޽�pz?�磻�����K˫��m:�4���'-{)�!���1�H7Aط�R�0�LB�y�f�z7ɗ�rz�a�,$�����Y��=p�Mv��m��[58V�r9�N/_�h�ݸ�~Z�L���4ޓ/q4t����+����e��@�\�C�H>��t�w�AOJ�@� ���X�p|k���ɠ��jd���(J7��l�J.�u�y��	��F�X�� �%��ޞ��U��&O#DKx����V�m���:�O��
iق��,�mC�f�C]J�R	~��QoX�pB~l�$nxVx��Z�)ظ���j�1��c�E�-/���3L�t��q��=��j�������&RH�8�h �}�ʇZ����B5)���:#�/He��dG�&����*�H�X���g�($G���@��E��x�{u�U��8z�{�m�^�����p ������i_ٛ����A>uho�+��I�f��H�c�\Z�m/��%���c�@��~Cȋ̮Pp2�;k�����?x���8��c���
ߞ�ᆓ2ߺ��`����z3�/���+�2D?�����(.����7�=���Y�����^�L���m̶����k�z��_�,�{��g�*��9�X���Uk��޴���x+��D�l<9KJ���Ƽ� �2N^�X����՛���3���DZ)qg 棭�~��d�~V��ƻ��^�R��m�S'�Χd%�U��8�
O8V�NIk8�5]���s���W��\ݖ�I��(ga�
g�v�S<	�ϡ�\�YPꭩ�=�dΠ���r�3���+�m�P����TIҲt!����d��Ҥ�ƠKܳaY ��ǆ�ϑj�:�B�+|��]�ʲ/�F~�BW�	8�1{/-5����j�2]��`?��яyZ*�.�ń2,�_h\���������D�����[N)�lȮ��,���D�@R���ld��i'7���*�W���>��\���à�$u�	�y�#L֦��.�
��`C�L�y�\� c���ͥ�P�W?�FC>���C�"=�J�ٓ�s&�{���(�WR8#�h��O�aj�$��E�K�����`����U��y�a���涁>��8b6�n����0��fI}=��!][����VR��K`�{/ �G0����z���R?��DPg>���*���O�G8*�;��7XɠkWj����0��$s���?�[[�Υ��K�=Bw ��:����G��	�ߋn��J��(m��F���(Ě��l���.Ĥ�{��qM��nx�}$<�7m]����l��D�d<n�oT)_iڂB�cʡ>%�_0��,*���\HVZ�:�'u&��dL���2�������/k�/�p�dT�lJAQW��e��Ӟ����ot��6_��C�j`+|�P�U����C0p��,"�0����ND�P7;���Ko�7�qM:�㟽��y��fa��Jī#JQ��P�]M>b@>���S��xiR��}�t��,A����0#5�՜V�&[r��C޿׸%5��5o��� ���O��f�=��/�8�w��ۍ�Y��ġ,�
1��?�I��x� Q��&)����Ē�L�f�JE^�Fn2��l����i&��E�&?�g)����O�ڥ�|J��o�-�o��gV'Y�5�D��U������~�խP�\��t�X�.O(�G�%��u_�u��ڊ��y:���?S��{��a��Z3ra�ݍ�M��I+���8�K��˰�������� em�S�.�L�&�����,h�M ���޳�/��^���a��Ʉ;��"��[Nz^j����b/���������Di��>A�YDc�y�f��*WCSX�ZI��ɟc���5y:K������;��S�-�n6xe�	����<�%���7}�YL*��>��X�^�P�@�6�8$��t�*�D��CM������ c�HD���k2!�+)m�JW?͖����w��lM����\!�j5��=�RpI������r4��b�%���o�Fn��tZ m�5p��!��x5�e�Gd߹�E)`����=^Vm�B��pz+��5�3��Z� ��ca��O/ 09�;���I��ތ�O��z�&�W�Zq6%C�oGw��:��2YGpV֌k��F
��U�f�AM���m�(���?�^(�|z�W:�t����s�s���E.����7�#֖O�}P�wd�^Y�����,./11% ��Xv�I8���y�߷�"u��`ܘٯg���i��AI_=`�s�
&�&%6�H8�����ᑗf�V<��OOΈ�"����\Me��2�5�q�Z?�J:^�t�H���A �^�+(`��м�G(�&[���/?�ɊLj� Mbƽ�~4�mN��zs�@E8��5������66֫����_�5����( {�G��p�˕�U�U���ǡ��{77-#��u�\�r�������1	����=�~	�|:�k��PRUEg�,���|��g�^gc��Uw0�nt���:.[\��
����bCy�sZ#�\�>�^�i�!�:5A幮)��J������T��������ʲy�=�OĜ���z�"<ח3��r�JMgg1�6\v���pw%Т�=��U��S(VMn�����t��I�wњ6����1���I��Q٪�����~�^�n�Z#�jX�GD{����K��=�hO[�Yxs`�g���:����+��s�9z�	��.Ƕ"Rt%�{�C���J0��M;tEZ���P�A��թb����|e[P��ʠE(b]�i��\ýϻ���y�F�#^'g�QtT6�T��.׏+26 a{=�,ǒ�5���v�ᅵJ̺�Z�|Ü)DB��#
X�ӽ"t%��[j�#�m�G�G��q��5+O������F�:�{&`o����/�C;���Dd
::��R�A�ׯk�(Ĉ�#{��U~k�A>��T��Pdvapo�����
���x�������w���%��7���_|�����ƃ��Ë����3�L�������b5�fQWd��⡖�ɑ��//Gn�F�����_E����ª�/ő�>QڍF��"��ǯ_[,2�rUJC�/u�ӭR��ѭԼX�5��gC]ݨ���l��fm�fGz錖��ƻ^��
7�jkkg�ߡ��k�ϝ��Q�����_^lol���#����6Rh0�m�-�f��-���
1[�"#��S�;i+����9���胦��kH��x�!�-+�X�)~4|����mDͼ�(�<�-�x�J�PoA}������B��~�ʘ�ƈ�)�IvȬ��
�����Mm�I�o���E~
���?!Y��u��k�x��'��ʘ�O�b�7ҽ�j���B��i�
�٨~�IJ�VJGtכ1���EC>��� p��?�q�_��R�2�6����As�x&+d�Ӹ��W D�����k~R�뢤���2�Q�g�����'��XI��t�xv��Hjg~g�bL�a^m��T����:���������H�ېV�v��8Ո�=ţ��jE��X	81mܜ��5��]Q!�$U_I��כ��'Ȝ,�s���zZӸ��Mm�TV�[ٖ5��i�.Y�Ⲟ�∱C:�=���.���;�SD�(�j|��xz�Wh(��Z"��w��>���~��ŝcf���#V�^�h�d��qz�kZ�.����1$o����5ɱCqI����#y�L��#-w2�?��B���՚��/�^������gq���R�K��
T���t�N�z님&Oqz�ŀm(
�!�D7�C>���{�稙�����E�4A`�\�+�u����h�{&f"N~E�54��ڂ��V�ϟ@�"p�Ho(ώ��ZC^�w,�ı��^�_M��D]�^m�e=&(�b����T���q\�'4���Y�Q�ʥE/�m
����+�A@\�>��U�`��]`12�u7���y�y���/�����%Ɗ|�V�}�V���/?�Y���T�k%��`X^�U�n���v
�=��Fವ�t���w5W����D�qC]��
JY�t�Z�;�;	g��[����B
��m�?/(��K^B.���6��)��c��%�ؗ��k}mV�G�L_`�s9fL�MNcCʨ��ID�#\c���z��������6�?���,4~Z���T�,����1R�d�u�Lm�V��)���_Ojץt.T^|Z�z�W���]GQ���I��@e���gb�3�����`ڳ�]^�?o���g��,��>���'c�5� ���&P|��#��&ٛ3��Y��4�)��>����R��Y�2�#c�3Zv�S�
wӴ,�����ia��R�'�� ��5RL�5����'$(�79�c	e�1�G�Z�;jW����:T1YR�u:^S��xq�P�{,�q���Xeޟh���oG/�Vr`3�GZs	�獮9Bs7�u��\7^?��V=#0��.�R8ЇQ�xP��r��AXM��9졷R��� �\��(�C,�����E��=_q鷩ě=����ej�D�2���{oA{�-|o�}��=�|�s�_�X:��*����C1qu�[k)R�v���Hw�3����;)0�q�<��hM��K��
�5&�Ä�|��uwF��A�a	L�B�# ��Ɋ�Β[�ү��!��E�$D���� sw�w�dH.3d��x9�Yw�7�n���QY�Z�9m��= �������{�uJ�i.����e�03���)نP�� �R��|��8�H���	�iy�{�O<��0T���r�:+>��g�9��~VO�#���j2t�3�2Y�����@��Ѝ�`,Q(��d3J�v�!�L�RmTl,�bݕ�N������w��5�K��ẒR���/�إ�G�h��q�S*�H�����'X#���U>��e��0�#�"�E���}"j�G�ǅ"&���=��{�\d��l{��tZr�i�N�c�����9R(�F��m@
�L��8%j]�6RT�����|�<�莰�'��sD��\�*���{�fۻ��4������];�p��Ή�KL����x������ќݗP��t	�s��X��T�Nƭ#�hsO�^2zQ��rBf���g�6G�F��|
Lf�_����|h��ۼً��"�<������>�F�ai�|޳���i؅��8!4�2�Y�(;��y9�����ĬV���c[gC�O��uF��xG��A[�`��{|zo�L�,��h(�?�a������C��Q(\�zn_�k_؅����50�h�m�
�:F&��5_V1U����V� ���g:[�v�"�����FiYR+�{�J�~��j*a{�i���\��@X<��|̲���l��k��d�������f3P��.����%�5T���#�Ͱx�����1~�5��X��{e�_�����~Y���7�u�l� S�f�ف��8�n�CC��3��Q3�AS��5���X<�G�(5����2�]1��r �X�A?s��/���!�(O����7���]/ =�Ȩ3 �g@���&Ê/�P.�@����L'ܟq���9ձBu;�K"�����w���^�s�<U)��z�l�r��R���[������O��#�{�]�&�^V�Ǆ�����/z.��������.�I��=�+���R�+\oc�O|�3䏝�������_��Q��u{h�J`�{U�����x��rv� �տ��2?����M܋�0Z���u�y�9�����ٝ�48w-1��P!�M�?>�?�h*QsW�X.����x׳zm�`f�
g��xc]w�W��;4��uF��P��l���F���H�;0�u�R���K�*Z�8�P_�2p7����?z!k��a/��|����/�*���I[1��x�e�l&������Φ���|�<ͺ��B��5��Ƴ�E��������m$�ۗ��Q�����G�$�d���r�� ��S����נ�,8���^�IAe�eA%�Pn��maJ�<�Ƥ!��>��Jx9�ķO�L,mX�h��q����wX���=G��T�&*.h�[g���r%vR�pK���K�N^a@L��ݹx%qa���Ǧ��^�^�7rD�/ôgy����Y��NZE���I| k3C���z$:w�b�9B�-�'��l��?��d������7��~g���|i1��T�ҵA���{!o�Ǽ3���m9��Åwm����^��*��'"a���px��k���7_�-�3��a��ƫë��)��.M<�7�z6}�11����Dp[��W��aM�#�+�J�NH@N�%�&�
)=�/�Bܯ��.�r8����;�J�/�9�c����I�⿊[������[|���Y�S�<����J������A4���k=ü�O����jG�s�y�N����>��'��#PrQ��l"�pHd�2^���2T�9���{.�0��K�X��b���,^�����6�J?ieU�U�+��)�� �v_k
Ѹ���T�*��jn��C�M��g��wT�[1�IƄ�PЇYh�tMR�Wz����n�~]��,�������$aK/9�Qfsh�P�$'5�Zjs���I�����l
��<K=j�"�I��j��^4�^N�'�IK�fͥ�m^���lQ8~�]����K3�<ӧ��/Z���ܲ��0��c��
�	:�ZW�M���{�$���zmcf[|����Gr$��<)����Orz�9�|��vwَ��stZ�~E��wt �0�!%���hAi�^a���4b��O�h����m����4n�hY��W��&Oپ)T*����kX��[?d�S�����J������UdDٹ���p_�"��[�W�1�+��%��-	.*�ώ����A���0�P���n��D߫������Z�#�����GF�7<Ț�l9�'pP�t%ɜ�7��lə�����V��A�F4U#i�6`, ����]!��g�rw�B�&��^#ZGL����j�_���ׯ�f�/���f΄?�9�<>��0�5�P�ey�)"���#��#�#�m��_{����4�@��љ�Waˊ�d�Ee�pgA׸-��]�2�����N�!�7ލ7᜔�Z=�7	�nM]ITӴ,*'Be��%*���<zY��YH���_��d�P�JM,7��30"�"���"�Zq�ߠ���1XP6�_=q�zҷP`j�M���c���(��r��ğ��ii.�U���_�0�����%{�c�j������"YgA�渦�l�=���x*!6��6��1��þJ��&��!���ٰ�{4�/�������N|���$�xu.�k㛈1�Ä�5i��R����~�<^^�Ug����H�\c����9��i�U�Ec4n���i��
�41��� ����!����TY��B�׳����K����)��!��w��T�5.�)$��d����1�S6q�7Ux?�m�<]��?��,�plp�j����5����%�.ׯkKhcT�s]�	Ǉ�R�NfJ���( �6�G��5�G��U���E��ض-WQ��mꆣ�%|�H�����?�X�����#U������A���-*(�56DN�.�H�7M'����'����x ��W�C���ׯ����D��
�$���S��`I�f@=leW��7l��0�j\�|c��s�_i\�~E��M����OL��������� �©�}ʞ��H�?��u.İNP���M�n�R_�r~�7|�zŉ SxE?�蔥T�t�eZ�y$W�����>G$�J"[�(Bx'>V3JR.�C]j�;v��&����NzpJ�4H+���<n����A�Vh��4R�\�'��^o$ ��gr�ޛZ?� �[��$�l�@�)��/���s9U�$���w�뾆�[#
*�.�z���d��t�4������*�g�@$gnῒ_�g[����P�\F�f�'�fD�`J����uM��	��v��1�;<�nb�Ƈyd6o/�+Ҩ�7��.�c^.ڰ��1�h�M�py�� ��4LNk5�a��[$ܦ��P�o�a�>���Y�+���L �����&����|�3�Ug����Mp�D�Z��N�l�e��V�>��\�W\�����a����9)6�RXDy�ti{����� ���X���L8·1��~4~�:�����Ƿ����A[c�!�]A^��5y^�����f2��c8fŴ7Fy�ba�N�=��	�j�#����[�����{�T،t��32?;n�Z+�r���Z��%�A�!W� I�}�W�+9kg{�^��T����o,
K�xH�ӞaupI�cE��xS�q�mU��y��F��/	u����5�rM��5���A?/���֣8>�eʑ�P]�Z��%��#����Jw!ĸu�����5�����jROƪ��]���	�\&~ GZ����[B%A��g��a�H�J!�������U K�������E3��M��@4�����v>�K��ohÜĺ`��j�'��c�B�E�w5�1��	�7����n�i�a#v�/䰺�݀��W�a\�N=��.`�V�U�LJ�E�ͥ���m%[��g ��xU�=�U.�ʟ�?�݂�w�e��I�Y��� �`�t�9$�A�¹l���PsP:�+����'�Z��5�t�Y?7g��d�|��g&ǯ���� �?��%�=N�bC8�}H�Y�{p����$`��#I8�	��0	'����{1	����l a��iL�,���4 a���O���}�w:��1	�tW;`���>h���i�.*���o�e/MK8-"�4
@���=|����o�g��M�UAEs���tq��g�Z�
����x�ʅp|K\�L�»���&������R���Xp�f���,|���Y��h��<������x:�~�]a���#�V�� �����S�flϿ�f����&̥���Գ-F��b	�?3�����(�%㔰�}�U�<�n��G2e�~�ٵ�εm�!(x�һ�N��$,o,J�}S��=���S���|�����y�F��RCa��X�14r�f���5��*h�-���8��� �з��a���:��/<���?��OK�OS��$��Z{+A���7��(ȯ����v� �}�!;���ˢdP}��%�|�4hY�b�Q�O���)��2%غ��%c#Z!2b?����:�뚽�Q<_]�A+�G6.윶'z���t���ސ0�Ϭ�4s]�"p�t^�w��=����١�|�c{�[�omڒ���ၡI�2���'�ٍ_�H��G����ҝ���_P
Rӷ�sD^4���}dl�l�#�����8I���Q�矐�t�}��<��+�S�?w��B}P��w�d�x_sP>�>o��9�qכ��Π�XJ7X>��>]}�O�N[_q�x;�uG/�Z�k�d��x����M)i{n��wm.\NU�S�����(��)�(a�?.��l�z�o�ɾ99��<p�իz�P��P�z��Ñ�}�P��4fdLqjzB�̠k|��H�SjwQ�t1v)��1Fk�L���?|z�5�j�aC��+��
X�l6<y���C�K�\���;�G�B���캿@��um�\p�{fS�:Z-%W't�/�����S�"UI��$,�F��N�l[I���![Q���Q���Kn������Q��Ypx�F#Рʹ�!�����<r}u:�_��&�/?P@��rgc/"��������0VSK ���<��z�F�/��c��B͵����O�A�:��9 n�����b���s	��va�~h #���m��3���8��&6f�\�I��M���Io���v|��ኊ��q�v�M��� ���L�� �x��~	�c�n����П�#m�͐%����{�c,R7N��{`��p�:)1�d�v���,mp߁'��	�;� HbE">I2��`{:N������4��l�ף��-!:Q�쳓����T��2�5k8u�����j	�3��7t]&�Ґ��B�o[X����xqU�!�3��M�|��OXd)�~E{c�s���e����Y@��-� 
>�!�Ĕ�oJ別^i3j&��x�"(d'`\(�R��}��l`��7�x�? @���<��4B��<�j1
.��!�Lt�y<?;�%����W�zr��e��5�w��W�~�p6�IGR]�.q���*Չ�%��Fy#௒$�Ulۈj��7�����?��ULka)$�VB߫�?�=$�JN�c�803t>%�7���L|��i�I�͡� ����d�,�o@}8�A��� �u��.�Ô�5�i�5\_���_䡊!_�q��| �ngL���	ݾ���͠x�%���6}�f�m���G �����Ed��B�_�m4�Y�L`�{������A�HmȌ������Kg��1�2�����,��;����`C�c(>��
f�C�t��-�F��Sא[`[T�
����� ik�PT��F���̣���s�b+qf��'�������|Cv��M"�y!8d-�����#�gC�U������_ �}u-@�%5�A�����I/Ĕ�C�|9��Sߝ�c"~��qo%[��a|���Q4�o��F�+ޜvZ@���:�WVa����6�GU�l���.ᵱ1���,,/�S���?j����	�b��Z�!�T��e~��0��R	�GwNb'��r���*�I�0��M5���VQIik]��-D���p��ڎ	�!Im�~��ʝ�&��Hu.��ؘC�$j9
�2U\)�*95}���&��o$��{+Y�W�9�,�%2�`r�L㚛 $U�
p�"R>}��Q�(�ߋ&�k�����Æ�C�K������>�D��*dX�Z��s�O�q�����;���rJ��m�p]{�$���΃"a�*�z�cg��D��!��:H���t�P��M5%�D ��L
^�#\e��ѽ�R3x.LGGA���U�p�Y�[+����K����!�Ά
	H�qc58@H�sLk�h�w�,t7㾟T-k��w������%$�ZwA�/ӗNK�{�i��щÌ��$i��>���)��w�:��=oSs{,�£_)�/���Γ��*��k! �E�T� 6�����T�&r�`I���˛�# ��ըI�"�~Qw�,|���t�C
@_C��:��|(��V�`�8�f�`O��`�?�G@/�0ƥآ�X}�|F?vj=����^�t�����~xv��j��1P1"�ӱs(�C[��W��m�_�QNH>w!Gp5ӵ$D�/bB��?�!�|n�T��RF�d�+��7(v�w�6YX����{>0����7:����c=hTP8�^����F��N�m�H$�D4���܇�2���66�߯�+o�����͋�')�Je"@v�L4��p>�����:T�6s��.]=HV;ޕ��*	6��I�c'�e�$�8N&~�A'�=��u3b,D��pb�dY��O(�J��"'¥б��wv�����/��!�1!����K���`�*������BC�;;;��8�02���L��B���1Q��@.'��MMVL�i�*eHs�;e�z�oX(���w�-)V��`�oÝSq�S�^��:�p�X��Ռ��-'�e�溛��l�r�x|��=��p���G��{ͭ��I��|lCCG�0 h%�>8�K��e�]\�͏���ү([�*������7�e�w�Ĥ�öJO���%���d�*2H�Ȃ  5�Q��Фu�5��2)��c��К����Wf�1*����nA�YapJ��ئ���ɽ����&j�ͽ&dЩ��p��I;��I\VU�3r�a��J�&�3�I������w����Ӟ��Ƀ�4�E��yap�L9�m�;��A[���$�8V��˛�*��5�!,�)�X��&�VP�g��>�ӗhܛI{��;a�rP��� ���2�2�EnK��O
����/���x�d	�#P�S~ą���k�D���?���do*�|Sƛ��'�	���
iw�u&I��
�ѧ��*5��M�����a�ȷWVvkSa�"�O������2J�gk����B����˯�.�oe�h��[}��٧�.��<������ kD~)��
�����g�`�5	Xtrg��7��������?�*���6�����ԍ���>�VUA��"���K�R��r�Ip�ߛ���mѶ
�8��bqt��D3� 	���4Ữ�-�
�z�Y�%^#�v�9�sj�f���%km�P1Sˢ2K

�N�0�"�9씷.Gc�P\�-Ѹ�d��"��i͞=�i�d`~Ӂ!���e!�٤{��aw�2��� ��N��=�O
A�1h;��#LS�����\p������(ԝ���g�M�v��z���N%	�뢤 ��~"���:\�&��ը�5I�1DX��q/��%�����K0��|/hmb�~6W͹{��{���p�,�H���q�ٕR�w�K�OA�xB%g����R�>M��(pȃ�R�B�K)�g�����{���'M�ei�M�A/B�f<J�<J��m�]>b#pZ�!#����ܷ�%��"���@�4����U9����0���P^		��s|��^\���������ߥn��F���b,���� ����d+�{o��"Xl�BoQ���h@ZP����� �pff|���=�ع��5k�S�3��3�'4m�If߹�}<@"�~>ww�00�1�rO���S��>=^��9���D ������
d����Ԫ�C���3w~����|e�*r�1���9``x��mFg�\�iA�n��)��&�\�ڟ}�-���v�M�N���b�Ц�{��-Ӡ���-I]�(���y�o�1Cܵ�qy:uǤS9Jr�!��C*ŧ��.dȚ�����a_3����2�� ]��*�����h3�lS�`�`�Q��sNLB��$��z#�~�s6q�a+Z����� $ei����*3hGV	B9RNHJ�Cw8���^Ȝ�� �w�u@��j��&M��ѳ���pG"�����ϥ͚�Y4:��p�o�J�E:�rY�4<�$��ݹy?� 2�*2i�[�e�$q��J�$w��[�\dͅ2��f|%�)���H|�,��추��}�9��ս�NJy	�=��:V�9@�&chϕ�EL-Rb ��Ms$B�˙?��P&}��P|-�j� @v� �H��M��7�d!
x�Y�S&L2)�I�r���hpb���{a�I��|��Y�k�^��
��ۻ�%\��j�<�!x�ߩ��'�[P�?ޢ���9����Ѱԁ�{�4jPٿH�.�S��I�%��]t�"`�i��;�6�>��g �[���ʢ|G�fAp��ئ�u�tA�2I�:�PJ���3�,��͆��1���#0f���~��*�X��G �v��c�z(<�C9�&O`	�?ׂ��=d�ٺ����F����r(h{[��Hԃ �zx;\��)ʺ��o��n�M�k:?@�!�c%dո�
&��M��6Gʹ^�Ƕ�c�m�?�i݄&<�N��'R�_k�_�@�:~�����QA��{BeF�t�e|��̤}.m���5����ʡ���c�n��T��^�?��ѐ3���"6��7i���̃��5�?U�C3h�-5ݗs;����̆D-�r��ѭ�S�_$�aTpD�c�63��N	���WZb�zG�!�r�#����.�#�{+'�&���Ğ��A���׼9��G���'ό���T�Hh�Y�U���n����Bv�ԔJ�r�����Ԍ;g�>��3���?��jI����Aj�b�T)���,{�fr�?U�Q�0�*_i���9}?S�[��n�3�evU5�29�� {M�qH�l��F�ѩ��pn���n�=pJ�#��2���/{�ހ�ɟ�-��&�X�@�(;�C��D�&�Ѻ�nkT|����Gݧ���ly ���՛��U�
ۇ�l=
S�S�,lqm���wA�Tp��i����j���'��rP4� 9s��M�� �k|�U#J���]BB:��$��,Z�?�]r�E�JI���Ͳ1���&��>�����B�D�Af�G$ M@"ܴ��&l�b����=h3:����p�w�B����x�x��92@��� ��9~�i ��T�\E�l©��[��kιr�T����V������ߎ�;mm�eY �z����`�_��N��9,<��lتt��1�zjzň�|(��\���.;�(�*���4�d)��g��z����o�f��u8�J@(V��������{`XA��"�gz��B�&p��:�F���V�[߉e�:=�����%OO���3�>�at�ڳ���>��]Pꘈ���,E�1}�P~��5��SK
�}�p�8���v�n-􀱻�7!=V��ͶJ���VZs�6�F�kF��'J��)�@7�� ����ݦsy��ׂ3}{����n�9�������U�vg7�k�< �j���Í-�`\RӀ��;��a�u^')��NB$"�K���*]B� g��4Gd(��d�������M�4��[m�e����+4�7�-��L5)�:-O웂����p�''Ѐ�C$�M�����p'�0����r�?޷�����Z�AR�� �
H$��!���̜n�_uғ
�|�S�zO���1����n���ڂhԡF�^t���Ϧ����Up�t��g&X�� K(��zE)� ��alV�I����d�\��j��$��V� Z؎󎎏�?�x�05���fWj�#����O�_Mڋ�� Q��R��~3y[)���ځ�յ��@���ho����_<r����Dp�MS�oɝ51��xÖ�:�J�Ts�����`/���t�Ml����p������
��{��2e��R� 
�~E8�ƅ��i�v2��kh�Y�`�'��#�z]"`��$�N�n��u�M0���5J>$���� 9���0.��P%����K��Y��T5�g� x����"V��)������6m��n�X�z�\�@
%dWzŗK�m���L�k�T<�@����5U�z��:�*��+��c�Sf���k�������PdM����(�cǇ:Du�x�_ �_<"�<A��^���m��"7D�t�.��9ǭ� ��e�fQ[�^]Ȼ߫*r>U��%�d�iԣ�?P]y�Al�5����(����-#����}&t1 `/U<�1���C�|�qK�b��VX%�U��5��ѕ6ˢh3Rf�
��2��z)�zD˄�����P�<x��E2D��f��7FZ�c�Љ�#T�J��vi��f���������	���y�=��Qv�@r #�qFqS4����͜�4��$w ׸|��N��h75H���:�GI�8[Tv��p�g
�_�Ƹ�Tp x	�c��h�y�dǥ�*��L7��µ��=Оg�C[2[�~�����7`) ��Wp3�c=ɕ)��%��z�+ '�x�����8���D�.5܀�W�y�6��W����֔��O���S����R_�Kؙn�ưJ��%Ĝ�20�d���H�b8}�%gu��5b�"PD��'���O桡������w�*�qʶ?ÚV�RX��H�E��kof'�SR���<ԥ�<�[ y��&�W̝��>ʥ9]6�~�Nٞ�r?��WJ����aZcO�ng.M�F��֤�J2�RM�����qCV��F���c?��WOq�c�Z�e��<��s��]�3��ܮ�:�+Uc��1EӀ::�?&z����b!M�Y�C�$z{����̨wΙ�WZ��qu(�������l�5�]���3�c<<{��Hcy2�����sg8�~&AKъC��C?��E���ࡖ���ZL �D�R�F����C.wzY\T=雵�O�l�!u�
��e�~��伳�� {Ƿ@�O�G&ږ�V1:qfʵ�D�Oq����g��^�h�̭��f����+[�f��X�� �C��n*��ѝ�-�6�U�%��!E$g[ߧ��p�`�SC-�~�-���ț_X/_�tx��D�x��b���z�´_���3�I";q�q����R�_�tpeggP@;H����g�֫ �N�4�������(�t�D��X=����zH-��Ъ�&��~Ѓ�����2����s������1H^05rͻ��0�^
}��.�~ƌ�%v�V���EhsK߳��s�xӕ!K�I�Piϱ���E?E�AGX�#W�Ҳ������!Ẹyv��UX��'�#I�qe�ރ ��J#�$˽;�4n=B�M�f�W�xޱ��S���.���� IM󰤣Ϋޕ�wLf��+����� uȕ���r�d֭ȟ����^ P\�#���e)�mR�AySa�7t�H�A�L�-�Xي��bE��x�  �	e��=f�z R���	ߋ}��#�$�[ ݴ}�b��1�|t'$�m�W}c�uXl���>������i��j�[?�Z�X���X�������&Lac�g��Ķ��u�a���|<5m[㍼x���E�afoȱYw٠V;a� �?�]�^�8J!I�pTpa <o�+� m��do��:�P���Rt� v�E<E;q���Qх~& ��e��1�DH�y���X�!#�{+izA�u{��mk�c��#T��R&���$Y'���P�J4�k�rU����E�Z� �x+�=��5%AW!�_�q�4t�r=$�Y���t��5�(�y(n}	꭭�SfZ��6�ʚNhH��`�V^��}����`@��	<����> W?�:����J��{Yotjs����b68:��p�R��+鼖���FD�z�:�?�J�>�q`P��m�0��-ߋ�~�X��w�$^�L������$wk���$�T��y�7n�ܠ��g�Fj��s�T��`�� (U���_��4;����#3�,���Q�u	���q��3��sO~'�u؟���)�'�i-�N��a�� '�ޅAW��@ilb�>��8ٵ�T˱��t.��<����]�m�0��>�I�M|��W�5�S@t F�R�)
���Vg��y1�:enq��Q.[��Y�P0ǟ�AY�6U�i�@�J����9�
� @<�ޥm)����A$��^��5�G�K犯w�f��ʐ�@�&�H`�-�{R��ޞt�,0Y�� W �Lo�C�?�Am�i������l��+�y���JP��nj,4xZ���q\G�^j4!���H� �73�6P�UO�����
U�>@!ͱWa �JL@���q+�_6d|�x�g`!���c,#b��0F���^�d5�p��l`��̓�0��\W`1aWQi�\-E�Xc�ҟ�KΦ6��E��
��H�#nNR6	`���#4o�}�(�N��|'��ٶ�d-:B}54~\�Pn�g�V��\-	?u��˭���J��=�-������f��U�-:4�lx)$WN�&�����Rƴ^d�6�6h1�/0�p�#�r@ImB�-ԩlmD�lI�����N�����۴���`ľ�F�bW (GC�B+y&"r�����-hN�=�� ����/�u�5�2{�3n>�r��rQf�W��&���
.4Y5n/��_|��&�^�
�N�K`�ȱ��_�]�N��?�
B��s��=ɭV���� ��(�f^p2���}ǍS�
��T��ؔ�<�kX�5�;L����I�_^�.���y�ܑd~�Pc��y�11k7��7�:R��A�B�ˮ O�ݙ41���#��p.m3Y�P�R:W�[&S�>>�jS0 ��h�}�݁{~/k�%�h@�S��r�B,)�;j�ښH�� �_�N{�4�S#�R!��F�}��d�P�������vД��2�Ew滲-��.l��9���9p
jЂw>�8�E[��r�5�K��Vg�vOy�v6�J�,���X�+��:�V�����ͧB�(�A=�ߊ<�V�h{}�J�����zw&�Ԩ�-R��IS��Ky#��@m���M����C.�מ8���b8�V%� .0��]�%*4ot�K��N���p��Y�E��z��EL��yG'�ۣs����J	�͖��K�͚	�9�()����f���
����7�����潣n*�sx^�D����S�q�_���|p����������C���b�c����Zh����kZ�/������;j`�5�Τ���/́�:'���\�T�naCݨ������]���݀��Ш� ��4m!��)��J�?�q��1Xt���۝�7|�R)+N��|��.k��w���uahk}�8 ��o��H�5u  �s%���d�n��3��qe`��s�;����	g��{�'��!p��f�|2���,�F�}��ӄ"?�b/��9��u�?��xF�x|�۩�\����k]Ŕ��#�'/.tJ9���o�w�m_��:+*�Z�ڨj��w3nJ�
�����ް��>s�ӹi�Qs]#t>�֡h�V~V�Ύ����J�C3���,�P�5Vc��ۻ�B�+;�K�nwh�Z MK�+a9�ղ�Tܘ��{�~�����ߧ�T�;���-�m���&1R 1�Еo*4^�¼;!���x���-�>[K�B�#���L֢���[uO�3�?��~O+�\R��,&4�� ��ky���t�=��h}��}晊�ɞ�R�*��RE]�2�:�x���4�
ͭ�k�x����v3\����U�+�GTH��_VO%�~�-
ֱL/^^1{�d^���T%�˥�|��
�ZYh�\�<?�1^��c�E�D�C�Y�P�5��/Ȱ��(�}��TSJ�%P�=s�Ȭ�>C?���_(9D��>ܩ��#��a�Xލ-#��:��d���F���E�M�(.UѺ2�#�`�R{�t���u%����j�]	LS�B]z���-�Mp���~����k i�'�(�>�ixW��%�y߸Ew��;��X�߫������3��"a_����d �r��!��?i"�r���PA˭�$�X��4Q/4|a�n>�p�O��z( f|M	��#+z������X���z� �u��8`�!z��|ʞ:6��K��l^X���Xh�n�gi�_��I�GR�0��{u�!uCϱN���tV	Z/��-��.�o`�B�E����U���ec1r�ҞW�?_E�>7��� ��F�l�vF�=Վ�F���9�B�����	6���}fĞ�%L�򴒆�jϑP�ę���ޏ����� ����Xd�rV�404t)O��dӜ�è{��%�ʍ'_X���t����؉2[v7�o�U�F�aX/>��:n��:�2�y�9�.���5�;�<5o*�ӕ"��S�)��Дq͙D�tw��R(GS�����$��8%*�!����^G�ɾ�
��6����9�6��{�5��`��w��T�4$Ò�9��_$\�i63+�V���A�v�-K�>o�������T�\ڻI�@o��&�B�gW��V���+3�a�W�l�WQ�/�.�ڦj��X�)�%��6�����ܖ�ә�m+ʾ����xXQʣh,掊_`�KI�c��̱�Z3�~v}ʴ��O�����=�Ŭ�[ؑ���譄֌���^���SZ�������<+���	����og�����1����Jy/�^6�R�o�j���`��n�s;���{z[(ә,wzZ,G�c�(�=�YJ
�k��zph���T������N�ZD�m�\�ӱ`u�b',�����K��%�$�,F�w/𸴵�-�f>���WS��>6`+Z#\3����J��I����am7��K⼣��^�k)�pF���G��`t%���d*z՗W�!(�,��N-g�+��e�L�ٜB��9ᛸL�Vie��-�&z�����f��ѓ ��LU�N��bh�T�Y�k핲���+C�U��0?�'�!r<pW�c"P
-��Ni��Ḝ�����%`ŝzt%���H��2nhz���d��Ħ��QИbpSG����3�q��v՞�����\��.�T0+GKcb&��pw�S�N:U6���x��2V�0�^�A��h�Y(	|G�$& ��5�`ҦSH�	�#�	1��E�)�L ���X�E�������>s%��h�<,�Q�������V�>*�y[�ל��&��~4�ՠ����g�q���ϕ(o5$�Rb`�׃XЖ�4<�0�ٰ���4��@�T�I��Ř�eq�>g͝_�:?��k�9|�.-m�9����.�1�R��í\ѽD��z�L0G2z[шo1}IA�����,O�T �*�}RñFQ�M�������F�Wriʩ��ǝ��݈�P��̝�LA@k�SE��i�G{�aakj<�ê�h���S���`���)VS3}�R󰾺�1^���� '��j��7�bMx$
���c����oڰ�B[�U��Y�~�$TO���:
=��Ҝb�'�oT9g�g�Z��GD�q�7"�I%�Y���l9H$���+�]+B鲥�gjx���6ԙ�*�.����|r>�(�V'f��T��R�ĺi-d�,p��feP�wI��l�"��@��yV�m�yS�Ȱ�s?PRHܛ��kg]o� VIe�jl�)1�J]6}V|)��,<DŃ�&�h4�C�:�h
GK �:@g	<Iў���F��xj<�3���K#�7)Ӵ�	Y��O/<"�x�am�v��e��Q,�Xp���S�.�9�������%Z�Q��"B�r��sx���*�t�!�:%�)Psgx��A_�����^n������J0����7�W̣,B�W����̝[�/���/P<�+�	H��������u^�y��Jg�Ȋ�;}q%߫D�܁V(�TN$��z�\�{Lx.98���]�=|����C���2"��$�"TiI��Gj3]R����H��:)����%O���u����ѝ)�f���#Ո���\�p6r�2<!
i�d�������i�@z!����bzw��y���X�oXt�lCE�.C�Ԙ�Ĵ�t�e�w��ѝ����PTL�I�[Q��ьt 1�g�yF���ˉ�h��>/�N�2�*k��C*��Z+���C�OOȫP_m�?��B�rW�(Ժ^ײz���F�����r:�*��]��ϩ�	�'`�_������[]f�E��w��vv�U�R#ǻ,kiǰuM�
�an�D�+F�S��<)�]6�����#e{-D!5�i��Z�E���b(ӽN�����.�_�\�,w��Vr�o�� Żb�[��3m��H���`��Z������u:1?-���%�������qF;�nM��yg��2�c܁��m:	�d��__�P�^m2��4�L�2����x�]�^���+�v��^�� �@$�k��2��@U$o`��˘�	K��O�֐�s�Q�W�Va�.x��<}^6���@jG�x�N��x����A'��KM��"�VF!�e��|���f\u��.��(�K^6.��c��x�J=).6�1
�x�z��,p>�<m4�dt��9��a�&"�n�od`99*�o�ݏ�Y��[<xhN�������9<6m���)�my�NH� )���c�y���Tnus��J$r��B��3��~T����I,0M
6pwM�`�˞AM��欥��N��^�s!�)��C��pZ!ڕ��1	�M�7@9�3��k�M�Ba�+e��i��9�-&���"(�=��˨6�N�lMQT�cs���#�iXk��QQ�8I_��d9w�80��?������Y˧�3�>�3,��4^Ԡ'r��Z�WFzr��|���q�F�O��Ou��n��1Za��N����\����cf���y�;|��d����v"B�~��ؘ�>�<Hg5��ի 5x���1:.�x�S�����l�a[��|S��/��[��hH�!X�
 7����A��Ӹ�.9>i�],ם�?m:�56�V�jaA�<��n#��S&(aS����}2$����Gw�1�{��^"�Vi�!�%��������H�A�Q6(u5��>���9B�}���:��l��̼�fyrD+}�ۑ���)ݚ_Y(-R��i^��ǹJ7��h���%�H�L�?��,=��|�.��ȱ�ez�$û�T�B0M�g�V}Vh%� !��qf��%jwǥ�r�[9���
��L*�Ŵ��������]K+l4/�D��_���dN��=��Rc�\����xV��Z�Ra��ߜ�.b�+��t�����[ݚ�^"�Q�Bކ���g�e�>��[��d4]Dk�)����X8��xv��o}`��^pϹgt��G�e�!ә��NgG؊��eI�ʝ$Z�qZ���k�7$kh;��(��m`	��\���8��H7��6d��	���rw�\���/��~�����6��>��9s���1pB��j�r3BW�;�bò���^���5��9�.�3U��!�����x�|���^���?�j�4*�I�8>�k��摚F֭c�����F���-*;�����j�s����7N�	�	�@,�M��Ŝ'C��η-F {|��иEk�I��Y\~Br�l,@~e?u�]�V��ٝ��3߹���Ic�kF�FD�z×�|���O[K��Q�X���t��s���[���1տ]�N�ki(�n�ւ��o����
��Ϝb�E)Ե�i&8�|�����}יͯ�����~4W���q�eow�憌z�ޢK�3_��񧨭R��<��l��V�!#���Q���R�U_�D�����5�0&;��=�<kG������l�e���p��΁F���<E�;~�SE�i���S�z�=�f����4?H(\���\�_�o����*��좬xڞJ��������{OH���Ɉ��	�e��|��	�͜5yZ��7m�?����'�E;��d�>AR�T�uqZ%-o�����M��/>qOa��%���V��W^�ҍx�k�(J��y�qˌ$#��k��R�L1���&���,�e�ٯG��T�4^}A�f:2��
h۪0��]3��m�c�����[���a��dT�Z��y�������^5�EUfr����'�J>���	�T�ڞ7F�ǆ#]ɲ;UB�F<����b����Z�nF�巐,����F|��?�����__��aҁ�R};Ƣn軆��t1��fDl*}����֟w���)Y�����{6:�;�Ȑ���w�1����c�z�?�_d9�d_�5�H���Ύ�N!������*M/d�LA�T��<JuxF�P�r�PQ��/'z��>�m.x��4���rՁ����[�eR6w��ʛMډ��;���w�7<��S�<�\\zJ�&{ǡO�������/�z} I����}��C�zшL��5+���}�<�F��m���P,l[�{헑�O�0���.�9�$�Sp��=�k?��Yoŝ �� EÅ��S��X�̀���͆'�6���ƌ�]�������Z7�����Y��ܦq��_�}�j�s��7��3����8�>���~�h��	=�,�CcU�}�O���+#Vp��8ա�MN�AW��k`׸��{*vXؠ�Zpv*Oi�߉�O)݈����@};'-z6<d�ڴ���
�o���r���ڭn������i�j��\�/���=׌�W[.A�d^(�E������[����ڣT���~�y���T0�O gI�h��-�KN?a�	�|A�Ghwk��M���N�7���l�P?P_�����#z�\?�Zf�NR�3���{����;hh�!�3����� {�Ks4��[X;������V����<y�$�w=u:L���̇�������A����~J�ޙ��糎�c_�,wj-+ls�c�=`��L�oKsi��"�x�ݻ�v�@d���F�3sv�B���S9J|Ď�E�5���,<!pE�\H�U1̥=����2��1��ma��Z����~¥!*�Jb�2�:�e����4�����a'�N��8et�K��K�p4�c�@Z�l�����~�*����3�tF:����"Q�_����}'�������~:9�P�=��D����d�O�M��C֥�vZ,�\���|r��Mn�ڙ�!	�z��󒇁r92Ux�1n�m�8_t������ʹ�@	��d�'�;P���2/r
�/�EE��~X�Y���m�8�g�`X7�c|���_ڤ֩���$�H�aа{j�����F�4_�NG
���]g��e�wq��8^�C�]���4��i:T05)U��U��O��=��H%4��t�!����S�Cή�sU_�܈� �a�w�kc5OE�ʹ�<�%���
�����}�z���z/(u�Q�گ��^�חp�ԏ-M�p~������J���x�����]��w�'+%�U�0�?�jU3s���CQ�h�g�&��̎L�J�bS����@Ce����Ye�E��F��G��U����1L�Ѷi@�^��p��������o��3�h 8�zȓ��oވgtT+#���v��@����+��A��i��3_�@�Q(�v����Ѫ1�����W\:��Q�Uo�9��v�W�U����K��rVł���t�tW;�՞�ʝD4ML�A9��J��s)��%w�Â~p�̝�3}Y��ހ�EY����wG��~���,���3��	��v��i�D��GN��B��!��U>��od��[���	�����m���6��~����h����Te5.j�9��XP���G��U���Р.�6����5p">�� a|��-F�1���s*Ӡ�YA��АW{U(��|i���'����?�'u*�
boaI������?�/A���{q�Q� 6��*uҿ���J0���4�2�riSşm�Mʾ�?tNuL��E1x>y�/��X�3�P�|>��?��K<̸>�m�r��a�<O?���$��M�D���l%���#�[F�)k�2g&���<�7:�p��u�Va<��� �	����&�tb��m
���m6���Óuv��Jq��� ��y��c
������!B��>@��I�H�ܖ��b<EmG]�i���^`�#��Ǐ���|3�DU�G�Te��s{�g������q�O�D�����]rmr��Hㆿ[T�ȁW�cQx4�;<����&�Ᲊ�!.��O{�\����ʸ�o}R��B������g0�;?�pR��K���aD����	*ǣF�l�E�e�������#�Ӫr���dP��e���ϱ�@��z��z�K����W2u�}`{�F£�6T�ڈ�ZU��GlR���̊�0���y��XH?��m*|��x�^�7�D�_�#�/���Ar��A�_���I�k�W����S��N	�[on�����?�ϒ�c��n(U_3�3r��M��̽�S�{jw��Q,�<9K3�M��ڞ�]����F�m�ork�x����{ӔX8	Eڤ��D�����z��0MJ�~����}���̽�U拆����S���N���V����{�,�%��{��G��'����Ny3$����R?��������a����X~GP��;R��s���J���!��kg�&5ǡw�<�`���o�v�'s���5���k�P�~� �;םS�>�0\�����DL��Up�/��Q��=����%���D����������˚���}.;��w�\�	ioЭ:��v�+�"1��`�\+;��|��m�D�f�gѷ'	ܢ���Z/�[ c�"t��c.��;���S�k��4<t�$y�1>G�%���Qr�{ȢylIz�-E�?G	���k���(g���Eh�TC��/GP�l�3��P{9��9������>�e��ƿ�:�����'����O�$چs#�ی})�%���Lf�$>���03<�v��mK��>��>GU�(��Ak�ڧ��O��X8�D��!m�l���1z��:�H9�-L����0x�w�o�qG$�*:�Z_�x�7�K�J���t/\��B���wi�&]�$����pu�
���s	DHY���R��d$�[F�j˛�0�x�F<���7W$�ä|�X0�͂m�ˏ��qG̻���iE8}�����`����9o�q��3_�|(U�*�օ�(3�Mn���"��g�V�֤A�$�ݨn�v�穅�9�Z��g|ޜ�x��Vy����l�����ُ�d^�e��F�/8��J�n���l���'�0�3uv܂�Rm1eLW���>SQZO�4(9�;�ֿM���M����'�d򟐩��7��_'���+��.S����9�x�����sQ�.e橿���d�yJwI>�pXs��PC�aǫ���2����E+����$��J��㳫����Wv�Xt$ݡ������Z׮y��5<R�x�ɟC�WW�ܐ�Zƨ)İ�(k�k	Lu���Fi����p��d��ɠ������M(��]�#r�~SM��	L��E�y���
ZKi�A��9~z�}��;D! ɛ�{�����ޕ��.U�2�ԯ0ye����8\�,l^8[���1�{��"��J�/9��"��"�\'�m��&1L��9�<��
(G�q\��`E���s���P�:T�zx�W�+¬~{`6�A��4؟���qM.��5o@/E7١j-�T;[�&�q�-�Ak�͟�C����Ó91�`���c}�FP�Z�^m���4�v����d�iQI}�z���ÿ��C�!�y_��/�V]�/�=nJ�n���)=�؂�R�^��W�x�F9z��s�l?`�U_Ӡ�|��?�U:D� ��@��{����%g!<Q�A�����j2aT�!Zf̑��y1��6��25I��B|M��4Xfb��M�9�h{}J��t
}>���1X�	E�!��Ft"��Wx=����I;�U��jy�h�.�|�
���;k�;��5R׬�����.���v���������_�$�~�yf�J�^�S���5�W��Nf�S��/_/.+cNMM�4�h�����q��"�������e�k�[@��MS�Tn��I�*)*�|��,~r��+���_��si)x�Z[[+q@�U�E����wFc�C͉ol�T���ȅ/%�(r���87.))i���쌳h�o/������C�e�3K��щaFy@X�֪q;���џ�F���ˆ+Gw>�������fgei��q蠩l�pΔH&r�������B������A�v��I�A_��,&+#�aw�hq�t�y�=�9B�؂���������N��N(�{�ʘ������v���%�;���эV�u��q�<�m��4���2`;�f�x�䅠�)�[�Ȓ�J��KtOq�f�N��?:.��K�!��U?U`u��E�p�s5��Gˇ�.Ec��Ԥ�O����4��)W��(�+`Z�����i��V�U�C��vx@k��b�M#I�{L����!�A��h�l��:ʣC��5��[�=X�)&ٯ��A���1<v�����+x���Ge,w~ �F��Sf>����"�o[���jB�z�|V�|�����wHC�?�-�	.���+�����e�HђKz��?����w��d�R��zG �#mk"�v��'͛�.\GPA���#�?��v���sL���� u��թc�@//�w�!�b�n�#S�����u*��'�|�X5��+Z��;�^-�h1S��%��B`�.B�!�{�Fd7l��=�S"!. 0�1��/	�0��&ɑ�䬓+�WN���'p��|-6�+mT��WA��[����و�Έ���q�O%)�$�ڑ*&0�/�F ��h� �rLN\���U1~;b�y+M���wD�T���i��y����u��WP |���� �R�I�Nj1"��ыk���X�:SGt��{a0ó������OLZ,�iz��D_�O��'52�l���td"
x���������~����)��@���(:��#�D���B�����3�t( fF' !"핂Ҫ스Up��:5( �� ���q�v�oc�Q7'q8�T]r��	/p,q�!9J��hը����3F�w iP���D2��F��x�<D�),i�,�����՚�͎Et�M�԰0.>t�`�u��O����0�����/tP�6�o����ԩT�N�����-�.��hB��kt�вګp�7FI��ź� �����~��u�h�<�34T�B�������:�>׼���UG'�3�- �Y�F�����?N?y�D�����b�j`�V[5梌��A�K����ccJN�O�݊��mO?k��Zs�i�g�M~��v�G���DA��(T!�N�#:K>��8(�鮁�lk6{r4���#�4�J�|�=?�Z%߾]�-cZĠ	hߑLEZ�h[�AI��T��0�Ù���NM8�N&��nу�O��2Euy����uT�J�i�Sj٠�s� ��J�㥞��	�Ng�/�}K�n��)�99�W{⟓�M��ݯDl� U{��&~���Z� ��(���ǜK��?���o�e3�=1�<&r��jaKgEÜ�.�a�o����Pz�|h4r꧀���0go*ʺl'�F �ڋ8"x���k�o��*���z��� �p�9]V�f.1Ul�Q���^X�h������U�2����
vS?��U��5Y��eu(=&�o��g����TGB�T��6�_�)*!��
� �sٔ���������'y*G��Y�A���P"�@,��/�yD����J����q�$��+c�+%E�ȱ�hgr�4$R~�KS�����*��� ���Eʕ>��H�Ne�f�g}����r�ؘ��ġ�{�b���a.�վbXH^ X��)�#.�kXnL��e)@�.Fr�,��+�JɎ퓉�eA TوJ���d��	]2.����(��c>� ��1�܄�7P /xY�IT�U��=O��L�\���}���O諾�XYpUޔ��j���W��w����.B 8gg�N?9V���G�1�W7�~đ�s��	�%���b�~���OG=����V���+�h���9�<�^l�V^��1Έ0UL�x���5f��������O����5������χy�HH���7�b�X5N��<�:�YYu��i�������Y��jsǓ���}�!Y�3�.l�@xSP�?���g����9�ޕpw �,�(�Tj�V�+DSk,-@��х����D�<ԕ�lI_�$���dBJ`+��a|T�v_���t	T�_�n9OQ�5��=t�<�,x\j}
i��\����4��F`Z�Ӛ��â����x��sT�p�*��	Siv���$�]�v�G����X�Gp��^�w� e�9��q����w���Gv�ǟ���qM��|P��RR4��pJ��	y4"��s�(�2���1��	�Ikh�(�A��s���>��FH�_�g��������ѷ_42I�Dw�H��x0m�9�kK_��4�\���!���Sx�s�]\�}@�4��7W������6�����D`1|�����Q8�%�>8F�)wcr�hk����:n��M�tI�	3M�3�t{')�t�z��V�	3�[VM��̴y���)8���#a�G�i�6r'�}1Z-YhIv�4�}��a������'ێ��O�<�G�f�b�c�
�K����k��<8�����~E�����'��Ø!'/�w�4kq�Q\K{�ر�W��i��/��(=$̍W�Y��נ���1�$���?�!`޽av��w_܉�զhF�1b���O)�E�P��<^�(��͎���*�x����7C!u�c�ku}�$��_�r����
�Q�-��������2�#fk~���z��g{����^�0[}<�� �_zu��n��9&�Y�q엤�#�/l�}�4��/�G&^ׁ�4���}��vb�z�X�߿�\�l�2]I�T$��C�O�O(�����-��ᖍ�����A�-���m��=�ֽ��E��!A�W{׏G�v���)�O�����~��l�u�_<'��8�յ(5i�ْ��^��.R�Get��^;a!��p/BBs�;�9���'�>ۃ�m@�i)NDY�QwEb]^�W}�ŝ���-L�G5a�[��gy�����}Gb5����'1�x!���C�$���c�4���M.(����u��#ǗIᴮ�k�����	ۣ��C=��'�T+$@�h��l�?���DS���G�`����_�,"_�$�jձ��8&��q�%�Q��Ɲ@�H٤����ax�ջἂA��Y\�$ZL&��)����` ��Y�ɍ�V��>���^��Ͼ�>(�4���3,�
7�<vp��0v�yp��(E#��]�lBu����3�h�#	'�r��m|�}LԹ��P�ҫ����u	������+3όc�{P�� �������/�Q�$U¥�/2���|nd{'��ـ��BM��`��oI/5���^��֓6�$T
�=�r@t�Zh��tM)K�{��]�*wo�#+�@/&��I�нNu�?"dw�UP-Xhf�������;X����Ŭ3�B���q`���	��)f[���҄R-�����2D�U�-y�7�z��<����IQ-�u�rY�������|M�E���A�D�0�&Н����p!2�M�W�2��km��Z ;XK����"HC���|�n��ˤ^n��Y�n��I�jڥ�au����I�&����B`����N2�vZ�����������(��L�J���Ȭ�Z�T��{��=��G�ӄ�Õ�~��e��[@�K�0-6AU�l8s�쑪�'���:������j֎{�Bڰu%�����"�w �P�[ʅ̨�`!b����ӿ�r<�G|�;>��z��'��$��ًT�#jT�·��S�1[��k���Lf�O���\m��ғ�;��|&��5�^���l?��mA��wd�V�"�K�"���'����BY�HF#���]QW��h��z�s�bq"�Gt��h��R��z��V��IoQ�!6����Z"��|�=��Bt�y���ҁ0���������#�/��R�(���7�/{��hn�+�
�k�zB0�Bh�;�=�\<� �Y�/����Z��LJ�ƨ:%~xv[힨��]���«��8x#l?��gߘ�0N�KMr���u��_������ZԴ}-���N40R�_�`��o"�� �Z��3B��Oj��M��:�.��(:�E��]���2�>,�^�ޏ��T ��ċ?��!��Ȏk��Bc�ф./�J���r;�Q����|Gd�)���)�-l��4��xf{�)G��;H�@�9�BS��QL��� _)�?�����t�i�e��q�4<Q�Hy����?`�<<��gUP(<�NY��F�_B����|�y�J-y3�q�W�"�O2Ǔe��z
wn�B�Tgc�e�q*���u&���7��!x��'"�c?�e����ۈ9܂-����6��u�^Q:�q]cl��+�B�.�f( �hW���_��ی���O��9Pe�[)���c
�}[/�Z��ӟD�B�p-�M}﬎@>�u��3��a�&�蝔�S��mxgn�y�m�%dE�7����-�ޯF����8�s��׏��o�K�V� gs�-w�p�'C�8?}�<��o��_ș���D<rI���o~㵎��h� n�z��-w7sӨ^�{yb��9��}��$�˘O^���F�J�#�ɂ�E�4��n�6�~�_ ���5ۿՀ:��(�,�C�M��c<>���]�
"!� ��4�½"1��C�9��-��{��+��Mn��˝�}�c�ps�L�U E�h!%ቚ��qɣ]���X�+BQ_)�C�����[�`��:00N{"�O^�dB;Wq�\���q<��Ë\�EZ���w���Wi� "�0N�R�0�&��wq!���2��� '�7঑��?k<��؄��9l#�e��a$,`�A��9���PZ]9;������ �O�R�<���,h=>{ ,<7x�  ���g��A��2y��m�T�w3~�0x9�0��l����ʸ�8��ݖ~���AO���\_]ഘ>�7���I�����P�o���!���di�ʮd�ZRI�ʖ}ɾ˾���P�.���}�$E�}b0��`��`��9��<�������+Μs��}]������>G$��v�n�,>V������Vx��'�������
��~҆��)h1�'�d�w�1�Uq?
���\Q�n&�<''���2D���=K^R�<��Ot�޿�!+���k��o)����4lF9����b��@�i��H�r��T�?���\�騊�e�8NN�TI��E���������Q�x���S�~�j̑Qg�!��k�~�u�^��~��\ �;�5t)����*u��=�%�5�?!�|��z���q���dvQ�[5�撶�Q�K�E��s%S��j��dV������]�3�߱ݳ0����u+H���-I�.��h�V�"۝��&NP����DW�'���O�D���/`)����Ǡ��n'}���<�M�<8��	����?�8J��n����vD�!��� �@jlF��F�T-^-��a�T�bF0�5��x��ӿ*��~\�o��M}��|��L$6K������;��	�e�g����w��K(9Q�z� =�E��y ��`;�����a:r���&T���En���^�����)�k�P��%�
v-(}B�'F}�G~ȟ<& �j�_j��&.�R�M�2d*G�����Ɛ�6��?}��;���>�b�_ �(3�h��^�S�8�S?>���&_���/5�W�
}�sZ�8�9��/��s)��_��_���#h�HN6�PȔ��|n2P�q���&T��`��s���NOM�U��q��٫��e�.���>X��X%�&"�^�MB�� �{6��L���%�f�\���c�ŵNOB���^B�	�����{iQ����<�l��P��_�0��T���g8�O>��T3�R��a)��}�K#�m����+��#z�����4'3	�]�-��_�t-�{����M�E,��+��e`w��un������PI��������Y��u��?�n7�U��Km����?���~�-B����<���;�~�~����R�d��q��矣R��D>�$��ŐI��FȄ�I���p��}���~y�R�tt:�t�߄5������`�	ȟ訁2�wc��+�u���$�����I����������\����c;��\ur�mi����K�+����o7�w���,���c����0��^I!��n�M�����X�O8����	~�ء��.��PH��G� _���).-qLى�5ùLo�+��Q�%c#'�#ΰ��U7�Lw��s�I�L�Lղ�����7��aǯ~��r?Q�gS�5i|?�� �}y���z_��^=��F�p�)T�6��}tz+�K�)��g/@p��i�qB���8>��	P��:���	O.��ZT����2r�5���|����+�|��_��n��4h[�u�X�ϳ�n�폙�K��t�ݒ1�꾹�[2�tM��F�� $�)�jܯI�kR��Eg|Z��B#�3�o��7q#~z�}x�w.�9�ib����>�9��I��.�b����ۖ�Kx�O�RS]��Ķ}�`d�~��yV$��IP9�r��E�{/c��p��B	��Fdo% É���P�͇��y�bɄ�=2�`U*l��3���M&y��������j����NB�.g�f���ӛ٫ObH&%ނ������j�w��ÙͽD�>O^x� #Uև�5�d��V�71u��cK�����}�Xh��x���j��{�cp'u5��k��I1��ӛTG=��;�U�!��l�l���h�{s^P�L�Z��x�Ң~��I2�� �<�L��K�k�
��j�_"�!L�����-�D��	/��Ke�>gq
�l����!�l��#��g7�:�ҾT�zs�
c�u���Hmpa�4���d��o�yo���z�i���3x���?A@�x~9u�5�3�A�&�-�H'���v��8z���u�q��_e�?,c�>���R:+"���_&!��1+�bV�4�Ժl84>�l�x�~u���.+�/M����
�u�",�R��7���\���ׇk���oN�� o��p�ƠJ(M�䦠�_ek��]�bZ�#�j�Iˣ�̧���RG����q�4�7,T��ͭ-r�~\7`Pi��%8U���;�������P��Їn�#�r��<����؃kK���N����3�,�1cz�O�s^�y��4s�%[ՍKN̯�i�rHf�R��.�����jjj*�8����Y؏O���Q?�add�j������Z�U��B�~b);S�je��٘,-��Y�b����Ӯ�f-cۃ����đ������;�]�AUN��ܼ<k��b]A;��KnW��uE�n��O��o�����L=�%�94����uxտz,����O�X���c�$ hk�W}Z��[V���8�᳷���ݞˣl�o/~���_�o:s�1B��mD�Lƹ>�-����O"�Q貲��[�T����$�;����L�Y�E���l(�5pb���E�Q��@>u���-�Q�m_iAwz����̊t��Xc��	+��%�MF^��X��f���$�4�,� � ���(yR@e?/M�����c\�w?���ɢ333&�.\���.�n�@��8�([9�W�#��#�í+N��J/����'-��M�;����SC�4��a��N n./c�끦<���ۨV$��p�ȝ6���'�~��_>����{�p'��	�&C���5�������������	Q"T�0���궕�[%/�|Ge�N��P���k���t�����-���f��ne^�N{��8���r�T�T�z�h`p�zo�X�e[�͊!Fո���g��)�pR�sXC��R��SW�j�n��K������g���L���{n�6����}�qp��*E����/�El3��ҰgO�q�5��*�w��@Q6��wv��66-�����M���k� :�G��[_i*�P6�bx)y��<���\?˻���
��)	�`���j�d=Y����Ƣ�GtI�n�4�#ܝ7J%�jp��	a����w����g����:��XJ�T�ݜ!v{�B�q~<Fqo� :�+诋��9Τe^=����h ��^�'}y�%s�A�ӊ�l�����+������s������@<�b�K��L��Z�$����D�/=(F�{�e[d��PZ潅]2ɴ���477W޶|G "��݁\!8*)9���" �4�@`3�Ck�;����sK�<PDdޛ�ٛ��B�}"Yw��T�4Ҍ��3qI���d ڨxߦ���Y�#̀�xWPP�����&�_��y�Һ��A��#�x�SL��轝�Όr=�7�i��>��Oܙ�~��hi�q���DX���`�����C��·ӈ�zr�9�+�|�x6�4��]|ZN��A��5 #��/o�]��3D���_\�4`��9�G�8�h���厝c����l�!�?''%~��=4��6�n"�dм���r�-ߕ��)|-y��W�_!X5�� G���h�z/V�ge|b��;��GA�9��V�4���oye��W���c�X#�y-�tg�$v���i�ţ���o"/7��뺁�����L-�s��k�ѣr��Hn>U/p�C6xy3����mBh t�{�o)���Қ������]��5)�V(Z1���ty7�"E�fC���p33g2�O�0ۄH���8Z��B��/�(nX*zM�~Sj�۽��H�.je����oO:ל�_r0%���u,C�1u3{1\�⏌��h{����NН���L;�G�FV* wθ��I����$��;D�Us�^-�-����/�c�7'#EeX�8��:{��9�{HH�h��I�P�bS�+!!���@�x����}ܫ|SN���FA[Ӣ[!��!ؠ��� �7-�{k�X�y����� 	?a �r�"�:݇�}��K��T����RӗJ�c��H��}cz��k����}��M�b�x���E�j�3���Vf�c �|L����ݗn[K�*gW��Oȝ[#W����R|q�Rз���q+4��}�Ri���M�6ŽU�`X!���d��D+�mM'R򔁷&��	����5���o``�D����O��+����U��Upے$��h*�5�>���p"���Y�As�N�4,�n�'��;����:ޑ~$zj���kZ�1#7#K6kA��P~ Nܿ��W�UJ�"4,��Z_��꛱�_5l��7�nN}4����$��J��q@9q+�������͛d�?�Լ8�(��"��`��|����ؼ��a
e�2S�^̧�������$n���\�B���P��X�jӕ2>ՄP�uE�Υ�o��%S&z�D�qqj"[�����;�؝NӠ�HӝDI�B�h��*U��O����D�h���*���^�܀d�Vcގ:?kmU9M�a��Wy&�|���###��u�E�nI�X�4wvi��M	Zv(��,\R�`0�!Be4T���8�������lzF���%��e���s	�	Sp�%/L��-�`E�~FӾ<��� �����0c )ZH7��M�6<nɈ�rb(�id�Y�"r�/cOʷ���O*�8��醌ע~������ﱦoRR�w��c�z���B7�R8��1o�L� �w�;a��s�؇�Ur5���ߺEl%5��"����=b��V*`FJa�-sc�b-�&�����5����&>�x=_BW��C}�<���\��HB�Fp�_�D}�=I��/��Z~�:}'bё���|�wR]	�B��� ��mZ�,%�����a�Ґ'��D*�m���OE�V�'q˸���T����\�����&��QM�����кIic�rJ���M�yyn��*'�U�\_��X%�eߊi�}��m�?����[�t@8���~o3�@QG��h.��_6��7���oRӤh�����9��8Y�aո� _�A7�ͽ^1$��p<�O�W���ƌT�����څ��&͠�W�������mT7�Kn)2�4�l�ecOx�@  ��s�vm0�����I�Ҿk��o:H��5�����6��q�@�#ťi��4`Z��n����C�%EF������G�l�l']}��d���/�U}<�����cw��������U{\M�׿�~Y_�x2,�_𔋡�K񟝝VR��ԗ4m�{Ct�7 K#��uH�n�w�`4�l�]u��M�ai�޹:M/;���r��R�����D�S�:!kW@��_ɡZ^;�|��hP,&+{��	:��/��	]����ckhc�Qѽ�݁�F�.�b6�x��
q��ЯL�v1v{W�a���#���{���G �b�PV�B��]�"��A�|Ⱥ B񺾾>��⮇m��9HA@/�xi��:�L�S���ٞ/B.gl�\��[y��	�|�i�Or��7����	$ot꺝T���jd-�=��K�K��_�� 4������K�����8�h��cb������V ��"�zc��E?� �#��v�ǞͨY�UC�������W��3�/'���7T4�yx��S%���ϧ|��<�OY�'XM��J��4�,h�Eq�,ft��f��r��=E�9��82��Tb譧��M�EfT��y�z��Еc�Oݬ=v��6�rB�6�RCzZ�]k0����^��O����g�2����6`y�]��{N}��d�����I�e���76�&9��8M\<_Y��e�ș�G��70�*7��r�Y���^����;B�@2E�L�֥�G_8�)�!�u�� ����"��ȋ�ȳ�704d�le}q�p��}5��*��:��#-�U��dH���/׶x5#�m�j��ePvp�~�^������ʞ�?_�mT���FD_�Y q�=����.pv�νRǡ�k*���qh�@��7�)'� �N �ܪc҄K�Wb<J�Rxq˵�T��\uJ��\o�=Ie{��t��U��;LL�C�KK�3���;���z{��r7~�1
V	������f�쬶��M/��C��A��Ȼ;{K�y�fu�,�(����\m��x����=��24���n�W��O��L����!���ì�����BŦ�MH�� ��aŌb��|A$X�c��AD�O�J��_�7����H6��ɣ\M����Ư���-w�g��	�J��������QqqqD�Eč3:���)" �/�KcD���ئݍBO���q��yHө�dp�����c�;�|��n�y�#'��*��<Dp�2�-2�KI����b���?�^,b� �
[ow�����Z��[g����R��Ȍ�����ʢNJ����^�j�\��[Zc`�L�_]��zY`ǘ�t�p����_g��_�z����'��r!�_�{
u�LdV��7�1&�����S�S
�������������ӯ~���y$�0A��Δt4�rl1mlQ7!��co�]ZZ�f�����Zހ�^� B
�l<ѽ̭�a�P���k?
�z��ʇރd��NN�;���mY�FCą(s��exc�����h~qQ[�ˤ[�Mn�T����g栕Uυ���o���ud�($�vk l����:�N��J@Qe��.]�|99=]W$����|���DS��Qc�hzr�D�]��hO6F��	O>�U���P&�l����8�"��⁰�0���m�,�|;���/�Z�hި,���&�ȴ���I�'@�p���>:�=�#�C? G�I7�c%aWc��)V奒v
�3ҤLI�s��}K����o�d�e��3pyW"�.�Ąy��Ӟ^^���N���8�uKM��y��������7>~��MćJ D���]���f��2�kRf!�^���� 7Mز�oda�o��P������31}Ɔc#"G��ƞ���T&9��Li�A��]l��1rk�s��j$�␬tp�2t��-�r�-e�yόx]������^F��2�PE���.��k������|ۧ����~��!{){<5N�b���^"��k��m���c��U�*�b���P���Q�-p��e�n)����K]R"��6z�7�~�k�h�`c���2���Ә���̫xh.�Ю�����%F���ݲA(1�e4���wǴĥKYfb�%%%��f� 8��(.�+�V\�~ְi5�E��-M�p���z��r7T�0����q�32�w�,,��A�>�k"�팩���'8=5E��K�SwvG�t�ŮG�.�Wpx1ܯ�lV����"UN�Cr�����;Z�)~�����Tn���f
�~:�pϦ��>�@�x�"���8��A�'��,s�������_��-^��-������ew�'�O��=J�el��/�a�(g�;��7]%����1޸Rw]��E���&2��E޵¶
	=�1X�R����������e�C��#x+G��k>3�$9m� {�����ON�T[������~�S�tjj*�O������/�>l�b���|)��^sQE��Ǹ �ݑ���vz��!�[:�bb8T��������[�I!����r<�WUIzz{��.d�(��I��c�^�1��ֳɟ
�<y��qc�Tp]���Znq���1z ���O�Aؑ%DО J"�nl�w2��DӄF��@��w-Y�!*������[90��{s\Z�͆��� C���*�;=/)�D������E�5P��=h��q q�ҋ�"���~t��!�D���M)�x /doo�V�@�.r< �Y�W���!^����5����e��_�Z�O��w������{��t�ݛ�v�-�!J��!1a�����ўW��A���� gY��J�Wm\_�}�8�����`uӕ�e��l��r��j��L��.h�Z��D��f��v��t�q�6�G�*��D���؆w�l���C��/�k�.�~hȤ��"=���O�&�iԛ6���x#>�����+T����y��D��ŷ��Y&�<А��^�l������^����U��cR��|Qi���0U��� ��wd!*�Ǿp .�����:Q�L ��M�g�oVZ.,�d
�P?%m5��K�3�y����0�qؙ�V�9r�3����0�JgQ_^^~�~�X����is��n:��N��R6�PP�g	�/��Y��MNN�]_�8K�+(B�E�h���7���x����*�2m�sxe�����!��$w��mn|�uϘ�M(�;�D,W'�� �@zY[��_�wN���@�9��z�Ys��EDp�))����Q �� �Lh.�]%��.�q�
�=SPÔj�C�����}��BPCׯzC����ʰ�:�S�P�� �M4�G	���W�a� 镍��|zS�6����%E/^���˻��LMyO7�m==tTF=�&��ާ{�ӂ���^F5|�c�����4Q�.���tQQ�d��a���π��|`��ge@���t5��O��ry�;p ^D�Z �����v��6@6��2ǡ�n�:�2H$ve���uPI0���
{�1ީ �Ey�;��񩈨����T!C�Y�+)u �j���X:O��1��0�}Y�H��V[�����n��E�ʟ�t�U6�4����
s'�o~yYW����8�xc���##==nD�)ej��Y� O����@u������[��;J���Y���s�������%�&o��ء~Wf��}c<ژV��ck;���`�(D/��잞{@��׹$5��N���-r�L~��D^��f^?�i�i�A��)\=��!�]��n��qv��w `���!�sXl����s���lK�Y�Ԉv(��
{�O� �oiъ�^z�Jx�[�#�|P3o���jD�S���bccc�蛪]�s5��!�����A�4���S�yvpyY����!�ur���|t���IA����<ѐ�m�����F�����B�J�?(%��H�ಗa>�)�*��}4bz%�F`���q��rt$�27��v/).^�tn��@n��~��n���NkG ���n��?T�5+^A6QW��x���g��y�ƀs�ZG�Z�w�� ���q#;B�s���4r���� �e6�[
x�����X��M�P!����;��ixZ��7/��)^�O�vk��z^�Y��������/ ���1�+�V~D������C��ɹ�S\����c��tG�����s��/H>`aq�X``೨��7�7��w-A�q��V������ ����%�j�4���d� ����ghNQ镴.����J��8Hu�aN�� -|��@o�]�%�!JJ�ƒ/d#6�q��/��wou�^�Tx�lS����=��R'����� ���s�	H��#LL�u�l�	�'Bx�,Z3��<��f��v����I$��A�S�	1Kߡ�%��@��k؇��E�1Л{���sb|�L��� �A�o*jk?���| �ťT�c�ةO�Ү/w�L�q(ѫ{�iy���nO %�OI�� 7Ź��c��!���&Y�L[@��*�;a�tl�N��A�ɞ#���r����)�V4'�<Z�p!B)����K�f���F{''b��\�
��-/��PP��(4P�m/i�)P�P.���Ǌ󤧹SҐ5��mT�:�b��\��~I[D��~8��,���,��F3PL�%���.EX%�coŋ���W:q��0E�T#���S
4{��/䵪׼=��9(���$A
I�UO!��J�i8xx|\,<��t�(@��b���C�"����&O���}��50$3J�,op����@���ֵ�Ѧ&�<��2ẉ�Z����t�13`t�W�Hũ�����Cddd
������\�)�|9�9����1h������^���� �9�PX�xɋ*����v��vU�p�36�ܰ`��nKHHȩ�[�	t�P��K� 7�!}6~��ThEI�n޼��cz�~pFt�V���nB�h����_���(Ͻ�<IR~��8(�|����f`�������i:D�wo���䲒sq%����\ƞ��sAc���i������\D|��{���8�K�ƞ���\;����Ob|?-����i���҇]o�x�>l=��az[�B��.���xs_?ߝ�}G�e�[��Q|��w�+���w@�ކ��)���	��0�\G9�'mK9��|����~�	p0
p1�䨼�z^=�*���ɐ��K�L�Jq'�o�\�)T:Z0�F�3������Ŗ}�X����-5��=e� HUw�`��͛)MMʴ|�(�?G�~UN���D+�I��aB�<iD�8G����2 *hOEI�400�O1��Ki�L���Z-R�S_�~G�5(T��rrr�W� ��w��%̨U�`���]�.���l��˴���g���jM��g��Ѧ�����_���R+`��K�y'n���O6��4�E�X�:��x��ld`Z�!!!��Â�G.+(ht��f9S�U�d:R��������yy�v(	u��:Ͼhn��՜k�+!�QP�,Z��O&�[�>⤣�$|}�o���m0�������b�i@�-��j|�e���T��0������$��/������g~;~o	Zq����c�}JqG_<���Հް�٘&0�V�8�bu�W��G�z������V��@|ow�߀J��uB����:)���?c&���mnn��I�(#�J��ٿ���ټ�ѧ��ӓ���pd��U��S:�3f3��C��n���L��MBB❶�|_\)�Х�h�(���6�����(yo�q�	N���h�.R�&B�t�͟��?6�;{�l2 <ކ�v�@����S��WF#����JE�m�V3	�4�x69�=1a��fϕ�kL풀񯮮�V[>L����Py�2�\��:���L��{��j���V��W��o1�T����~�t��yb=����,JS:�	���M��K
�G>���?Z�`5P�s��t���i��۩���?�x��B��%T�W[���g3-h��3ʚ(e�?���ld����#��ņW�^�sE7��D��'���G�����vZ^��I�1d�8	%�Rb�B�e����2~o9���`c�&�z�R�ġ��bZG� h�{�H���g�&#�ֱ2��i|@�pf�j˶���a��]�i>r%ee�Ui��&���-��^Z��2�-�~aZ�l�c*%ݵ6Y�XU5�.XڀKv(�� �,��@h���3E
i�t�����������?���@ ��(r�g�_k@���;9�,��ө�<f�=��03�i���􅬍|��5ȣx�y�6J����G[?m�|7�l��$p�LV�Ł�)�aXxNǱ�R�4�.3Te�Sq}Z���~���Zx�,�-8�^�~�P�gRISmIG#�+/S0B��hD�̶����9� �Z��m����G�ITە־[]j��Q���{�׮��v���ԕ�ѻ�$'4b�7
W�Ҽ��$gLU܏w��\�a'�ߏ"HHJ��8#^�[b4�V��-6���Q޻�ߌ����*ǡ�H�y�;U�e��o���q4�n������ݘt�"	�yT���C�S��\��}���l�}��{t���ͅm��i=Gtw8�y��=ȴ+�Rc>��J�����x���#�wrv9�s����gU14y �ѥ���Bj��oı���Jǵ���<��� ���9w�<i��D�
'Caaa��������v��r��.���T`�ƕ73�y��i	u���o������C#,Nk�k]xg&�_�p��y:����bQR�e,�R�#R#�91��4!?w�r�|Cãq5���9uuuh�W}�^����?�����Յ/H@��F���E���uA_Hw�bc�nς�f���gH���0��/�[%ԁ�D��TM׉�HA�=%�n��`���`>*)3����e�HN�����������
x*��2w(��Rc-?Z�h ���S�黾zU�0��11F(�7!�o��)�Nd��fޅ��
���w@��,/ȣ���&ct@�m>	9���"q��h�2��_�:�	v��+Wtz�.vv���f����<�H���RM��898���J\�}[��⌡�˷�a�u� ���V� �ҩS-bo}�� �u�.s�֌�+6e|N�`��ÄW��fbZ�Fa߽r&�������b�7t��������aȵL�Y�L>����ձg�}����v�4	p'���EP���"�&S2�zG3#h{��W[J��lii����r�����}K�jM��  ��@�p�w��)�W���7lQ��v(@�4�U&��� YlG�0�����G�/7����
>o�v�Ci|e��zp���� M�r�<�z����P�����u�@���HM��v�=zSp�F�=|Í������ �@�p�T�U�_v�#A�om��ҏh_lT{?���z.g??�p�׍tٕ�:P�9 ��T��nad�U>q�C��Y�i�C������^_��m��Hˣ~a��1�=�Ҧ�B&.�Smn����oRS���3ihi#��L�*�ܡ{��������u�7�N* ���^��D/�����������֣����`(P�1�}��[�&������?z`��|��*�0���пvܤ���z��:���.%���.<gn��&�Mw.���c���z�5S�}/Χ�Ӕ�PFg�br�-Z666K�KKW��8����ϟ��o� բ�c�;`Jt�8�m/��M�>����cT0:%=}PM�񝞉��h�ʓ B
��[:48�4�!�$3��\ -j�4\yu�ݫ~0^�&��նP� ��Ÿ���~6SŧY=,w2,Y��<�6 LT%;�Z�B�R���Xy�1�=��dO����S�e���S�B=_��t@� ��Sox�X+�1@���VQ>nNQ��7��JUϧ�g�o�M�,_L��
_<��i��'�
ڈ�8>>~U�|��X\���f�����&�t�y�/6��}�c��\^� r�����{i����� ZЌ䥤��I����^KŦ�&�R=���{Z�_&���&d��� ���)�<�Ī���:w �d�Ps�s@��B�j[��I��!�	ך�*�'�����Qr+q���E�������X�Ƨ
PҠ�9M��_`7m�����y�7��MZ����K-�4#^GRu���LY�ٛ�f9ݐ�*+���xwٻ��(xK���+�:��\g���%��WvP�3�x����E�G�l����[��3� �1�k6�nᒎ�2u�tW]�2CV��+�������K��>p8��2o�C�C�95��Q�r�i\[���,���0���i��� ��C��\�1�l�9���K��ɨq��#-ҋC�cz���}AW&�����կ��&_��S�d���Ҽ�&�o���ή����6���Vɹe���[�U�{|��5��ds��v��L�e�s& S�zՀ 5����p�Cbz���&&������!JJ �O����~�q&���b����G��`�xs��!�� ��t7Wz��B��`�m<���~�$4f?�-���ɸz�N�+��K���j%��s��_��ݾTt�z���' ��EZ�,,�&l�A} ���_ s	O�1t����KR::;��O544�������Y ������ɩ��[4M���J����?@L����`l��#LH�����Ƽ|i��Yq�Óϙ���Y��$�0�+����v"���ƆL�$+�\9�S���؝)J����� O�V���J5�Q��׼�O?�C���SDw����-���*,.V���8Ӫ�_;��k{9�����vQ��N^8��� R
�O�UW�+k�鳌���?rRҖ0�9���`"�FGU;J�M�t�GLR�#Wkԕ��l��������X�y/�.����%A���[
/�,��-���+2v�j*l=҉P���14��ɩ5���{X>(ܿ���KkF9� ����wr��
�r���ݏN�(9��tߙ�`��� �{/lXe;כæ��������>mCCL�)pQ#�!��
Ͷ���:�B�o}��W��r�c�F}���ק�]��_��wtp��4Y����t��ͪ��Z�U��UVV^�b?�D�Nk+?iF���&�x'�ȑNk��㘪+���  �@��:��O[�i?(%_����ǲ]_�r:�J�ȼ9M؊��=8*�!@3�s?����nY��|g�&�JLVU�Fj�(��L�n>�B��d�X�����c��ԑ-5���� ^���[[�,оx�$��&���i䱦�b��. �wYm*������ ^�z@>�M��1)l�f�쾂p�
z�����?�۸�B�E�4$7`&���j|G�k��L)����A�gg����;�w{�$����rr�&7//�6���س�4�o'�mf@&<8��H��CgI��0/B;�.�>�'w��q�>�cXc�|~���?�T	��n������'K��(W�ِ��g�On^͈�rn���C{�`~�=ei.�rZ�C3�@O��`Y�h�#���Bx~ء��K
��웞g���)��4h��T��*�@Z(d5�������������Nȕ"�^������ni��>����j� �\�o�(��i"��7>�z����-?ڵPOY�Ӥ���� R-)9��,��cm���]�����i�hj膢"����#%�fɂ@�m[w���уX-�]��K�n�v�iT�OaKspd��+?���l(D9���ч���{�
򝾐d�Ԡ�X��;%N���q=]�2���w>5zv�������O�
���1�'~c��靉��;5΄(��h��'�����{�)u��� IZ�t�ֳ/�*1z1����_���s�%�A�GW9a��]���"�����X��о��"%4���c����Ug
�d�F�X8��ٳl�l�? _�	\�'���¶T&����M2jj2��^�Ue��S��]m����y��wX,�*V8�`q��6\����\@��+�q�s����Yޢ��?]LH;����醫�]z80�w�E�Y����1/�?&���?���¼�ؼc�"~�oO�{��Ͱ'�SSS���z��
~�ѷ"�ۃ���ll�L�ʧX�'[#;�i���́m���2�tG�/�WSy"Z����I'LՒ��]��I2e��[KE�rV�p�0SQu��d���sl��1QQv�C�Ug����z�= À�&C��ؿ�HVm<8B�@��6p��ޅ<{���y a�� �����Su\Q�Y��C��\�J��s�&u[A<
^�m��2���5������V+_D���8p�OeQ11X�.�ح�l����L������)==�Ψ���{�@$X�l�5b_: 4�ᶓ *|�N���p'!�.��Mz�OB����k�x���DQ|��\�fI�R RZ~��Y��Z���Z�l�ߘ��-�!�D[ ��L<��Km����S3��w���Rƾ*�!.�����?���F��m#��d��H���"}��,� � ���c;����v�oSn����������X��'�(��A����]�o"��?��y��ΜZ����m{g�_���^���C� (ȸ�rF�OF�b�u�����w�����ӏ=6փ��l�8��!u�7���o��4�&Vt]]H{�6%���焉�e�����g�΅����3���^�H�W�H�uj��|�<dj�!R������s�L[c �Z�,�b�X�#�ZUŵ}��R.p1���'�m��u�3��w�uI���iۏ,�g�P7e���[��z;q�ٺ�C��(�1�pzH1*å�w3MHx�s��	D�`YWA�y���ӎ�d�$�����zw�bTt����P��4t=�dp��%�l�.�DaΨ��jﮩ~0���f
�!�BBR���H�[��o-�(�o%Aqy���m��+��O�w�H�������fL��zL���20>�o��|��/Y`��|�P��0�����Z��f��{?aj!��۷��AL:n�	��4a\͌ �l�����Ù�9_�_&�O4Tч��(��q!�P�������\0>{(�������d���9)(�88/���#��'�9�%BB;E�Hh�Ǵ�:�q_0��{���nw=Oq �4���a�	�(������wҟ?.�!~v�w�|���9�]��Ib|~��:T������U�(5���3r뒞b�v�HBE�ty�^h��e��v>%^p_~��}��T�TU���C��ͥ���TWY>UMy��&�.~� B��)-��w��_B��[}��w�J� SqE��YZC=�B�J�R���*�^�� �@�y~i�f``  ��'N�|��ܽ6Ut)��ʧ�=1A����:D�k��v�>�7�hO+LD��E�|6�cpg8;=?����x�>���?t9lK�O"��6��}z#{𶔂B	�l#����Kޞ�v��� K��Ъ �ot���r´��ў���-���/�3g�m�zz�FG3?��I����������.Kоw��-\������%4��yk��\9#�uf��MP���[+eu6;����d"����Yh?����
��Ҕ7o�o�Y�'�2�&P����b�ofr�����g�ܴ��M�K'�.%Yd��B������}&�98X��m(D��B�۽�w��ʉ#�K��h�9�cP��E��%��'���w�/����y��'0���\�%ȝ;z`��ʇOq�b9&�e8����&���Ie������u�T�ZX�]���~>P��߇�� �����4�Ml��t�srptǝS-t���
hzs;��UFSUԛq��#��obl��t��7\��A7�%��1�a���='_�sv7�53r��Fi�P8�B �c�9�uu!���Sw�Hus���m�m�3�X�$c�
~���[u$dg�����q��˹ߊ�z_����S�ůƕ��b�k����A��V���,:`Z� ��GO�C'��>��V����
��M �;TU]�����Ӎ9΋,��7�I�n9~|� ڠ�騫�qm�-�'�*�����e�?��*��uC�JC�@�Ll7��(�9
`����ō��~=��(4�F>����:��Z3��HeM�cX�D˥�=��ڎ�@����?���8ύ�y(�.�R�5
&7>��j����z@e)&9p����� `\aE�b�i˄L`�6�ٳ��
�����:Ҙ?\���v ���Et$8��Kg݌�~<��"����6kQ���c�Å�bWVW���Us��)++�t�F�R3�r�������Ri�d@�@�[���E���q�w�#�4�p�r�D����!G]p �ju������c�ys~�fV����/@q��eb�ImR��.�Z�I�Xx�����D�Ϲ�c�{	P1�W2Bg'�m����l`p0���CI� KBX��KDb����n\0�
����!���&>]�5w�ǘ�
�g^tc��7��K�˲�EJ��b*�S���3���iw^�y�ҸO��g�Bش�!��d�3�Zr<�%׿��#����#u�߾s�@,����O������#�`�-Y(��ɱ�� t�~�n�ف������ 3��rޣ����i:��ՏGʁ	6�R/Q�	AVz�E�qoO��G���bޝqZ�90Wy{x��LEmFo�1q���;`LI�C��0Ţ�E��J�P:n�Sȁ�zo��O�7�b�:z�9@4n��+��E�8�Ή���쒐�)�����W;��l�B{��$��=:�L��J��Ó��l*  n'"���<S\��d���.l�n�#QOh6�c:�@UR�	G��>��3@�	���94�2�A�yǽq�o�_���2c<}M}I��d���T���5�Ǖ$�	|��r��cWii+��:�t��+��b�l��R��'����s��\�t�j'����os��M쌕�"+��^G�gώ3e����=#�\��z�(�/~tEDR	i:�[�i�$��Ar$%��C@��F��a�����|��<�y��c0��'�^{���.�+�n6,��H�&<`���ef���%�g8���e���·���U��VVy��9��٫Y�ж�$$nBi߿k ]:��i>ٟz��I������ǒ����&���"���t�_���������B�;��6��iأy�q�(��/V��N��L���`���6��2�wq%�f[���b8PVM�ke�>��qf�(#ro֛���8-�av �=���{M����Z>������AL��r����b��$b����!�΢���[��P�^6�I��0H��Q����j�eG±�:�>3?�,��3�;����h����[���D��/]�Z��Um���O�j�':�f8����߮�lo��͗x�*A�F>�Cm�BW\��p{������ P�������k�NcK1R����@�kHX��~A�9����=��� ������2�n����C�͘gG��_�˫����(�P'^�h���T��m�C�
0�8���%�Z�B[A�!"�=�D���B�x"@P�q̖����J:ٺx츂��B����X#tycV^&F�䠬֍�!�S�;��GYYY��� �ҷ�2����*'-���2I����>:4c+`�L�	AvN���i7��_�k֧�9u?�_������l��Y��W�vy��8��QOOOB�e����0�ttt��ɗ<8�o�LLȞ��
X�1Ǫ���8<~��ߥ���'t�b�z����z��� �}P����u�24��2�!� `�v�̽�<wRQ9v�7\Qp7��?Q	���R�Ӝ��'�!))�5U|��Ho��4��@cr��:�-c|
t�ҐG$]ݟ�H.�?)ᷮp�;!S���=*nmƅ�}]i�x����Ŕ��w+����%��n:P��G�ˍM��c߾E��F��Ӫ�d���r�ZҺ�Z�Z����	�U�����C�ŁT�@�%XH�/ޮ��;�M�r���y���
aT�:}�W�а�"��ma�I�2?\]�,,, !BA�P���Ȁ�	P�@�IH&�A��n"ns���F�A�I�x�ӵ1(p�9��i���W�uq�OWm��9V��!��Rjv���r��)@U�x�,@(���\�mp�8�����@����oܳ�?<�fq�@ �K�2v��'�N+��^�\Q��*oK&�Vne��ayeY\�����go���|^ʈ��y��N�-�d��Y�\诲�[��.���M��?����и�q$�v��#?I�db��c(;zF/%�gWQA�z
���L���{g�ūW����ݞ�k[[�Rd���9��ʫ�)V��~Z����;:3�������Ά�����O4�����n�"�+�m����u2���W�*�m�O�	������L4���;�[��|f�-4��p�2�صc�j�ʪ��wPG�,�ƀ�4	�C���} o�Y���^r�����L_Fu�{����.=O_?c�U���n���K{Ճv��Z��X�4�_R���U���d%�wQ��_?���s�D�QZ�3.�"��No��OΜ�<��|21S�L��Z�_/�ܝP6��XH�`ך*F�����i^�
B�A�,=�����7>&�vZ�V��*�^��h�PL�-�bmN�M���?���DEE���{�c���T���[�e]�IQ�J�zx@�1gxX�1��[�,�OAR��uA�+�,�h0�L��h�S�Q��<�Qr*�W�F�w8��<#�R?�8]�zR!�����[�)�� ��[s���v���8��qQ���O��N��#�i�ݻ��Je�����߽3�@�JP8W�!�[��M8N/:<<LP) ������L���&x���^=��^���M�̿��$"2Yu��Ą�Y��?��}z�Ҁ�l���������zӝ1��UW�H�z0���$���l���/�=Ugo��Q����ý��|֗'҂�יVq�Eݟ�3�-6���PG����1�~��Ղ$����w���mRv2���]!��)ᇐ�P��*
�!"R�ק|�uNbb������b 	��V��t�v��=�qLW����Cer�jQ��			QO�
8))�T�i�5��ڕԶ[`U��9)e���mL�@/,|8��C�n;B�B�QN��2],��Y莁�09�)AMGW`���f'��i�,{{�	�F���ޜ�Z$Hm���z;�b������J�=!�p����DHd�'�j���Ƶ�H��.�{��Z@�c�'r�ʁk�Z��: V��҂כn]t��;v�p����}��iɣ�N=r�O��_/@����S��'W1-���E	��C�e�9�dw���cE�ڀ#ϓ��ӲʃW��������d=���J���|�攼&�^�M߬A��Ȉ־�
1�B�UTp= �2Q�Se���ٍ�:�G&��+C��:*�?l`��V�Nqsuz�Ҳ�����D�o��ma\E���*��8Pr�e�	���ee�E��MMM_����A��<��QE������zӋ� �!~ʗ�[��!��RP-@�
�]�"�ݩ��V��).�����}���
$Su��;+5���y�pO�S�W/�tcj���Q%����nEe�ʏ���r'���ԣ���>��S�^o�^!��o<?s�y��f�>��?�O�PQF�L��������I�Pхnո.��}���B����F	�>Y��	��' o|߷��}{�!��٢���3n��������.;Ŝ�OԜ>/��h��Ԕ��߳�O3����y�ECb'�,��6��K����a`����ʶ5�4�nX2�su���O�\�����즋�/��9���־�l��_��݀��f���v���3#{t�ՍK��	�t�̇ք�_3�RT�'@:�F8�e�Yߖ)l�XR����V�vHVx�zS���O{�0�o� ��L�U��,hSB!z���qe��I*���:}�Y�����D����3�!�\�w��^:w���y��!�oʕ����><�Ndqe���T����Y�ʐx'�<lg�Y8�y{YӺ�~�rm��LW�Z���[�c;}D�K]2w@���"�ݫ��qA�y~�	�"ɖ5X?����B���7#�˫[�c��}�:�ThKw"yV|��&lޝ����痛P˗Zy�j�\��X��/�S?Zr[�m����8Pkk���B��T�^���ꂧ�v�~��EI&�o܍�N��K��6�
M�<T/l�������b������r��I�z2}���߽�����J-�X���ez��@��j�" �
eîk��uEÇQ�II��֯G��ĉ5�8&
�ٜ�D�o_=��s��2rSް��bu[���@�O�e(h&ȜӒ�5���Vh_D���<�=�΁U##G�ʊ�%I�����	=�b�o�7|��[��J��¹;�}��Fq�5X;���O�Uu�}>g���|��ŭS`T�`ޑ��y45�cJ�-`�C	ؓ�$��:�"���^@M�z�� )?�Ѣ7���P�-5%�����~�_�� U�y���_z��ﵜ.�PeHeJ�����A�iO^x�e��'�����]8ɶI%�,+������p,�:a�H�>nJ�zF*CC[�����k��c^h����j�'�l�f[s���u,���:�&�P�5C6w�O&�z}[x�[��?78�\����}"sOU�:�)_�8k��#�`�>�u��3ޢ��V�̃;��y{��{Uhܸ�a�a�9�I��q"\���<WP��0��w����U�U)E�S��Ӂ�����ޥ�-:X6��8��CH�c{�N?�,��:��YTG
tb}F�7d���I�Dc�9l�0�F���yx���."�;6ړ矿�j,1H���������m�H�H
m@H�i@�B��ʚp��.iC�(�,I���M/���qGVx�KdZ����W�����9@���]���+f)���U�,���DB�\�!o�Q��{�wa����t�E�"�-�<$i��1�+Tq:��]hKJURc綜V��ֈԚ�&7�G������Kx��mI'�~/	N�F+Ey��䒙���2��m��j|�����W1��
Ub�bQ4���s-Yw/��k�, Iae�r
tG�Ǝ:�I�@�h�ԛ�~�x�Y�j} 8���2��WTĕ����w�6�H��W�
�����i���['�yA�,��D��ϖFK��j~�&���Qﾫ�_�7666��׳:Yk�Gf�H��/��w�s��I���	�z/%�50�+�b����{MNy��"A��6  C���QH�i+z��a�.�b=A�Y]�Y^su@h.���BW���P=�c�Q	�N\:�Z!Fb��:v�
�1E9a~�\5�y%8����9�G7h�g�?�jb�^P�d�����Hu��5��Eِ���_�v���$�.��"Zh���gUKt��xF�j���-<+/-u?�m��^��{h�j�Ĕ��kӚ�&Z&[SB�wvv��{�����i#�5����]hߘ�>�G)��܉pz�iQ���*��%������'�
x��Ej���B�g}0tM{�ص���Z��D�]}���">h4�^YY�qq�y��L��ǣ>�89�v//����P������j�o�22
���� � HH\JB����d�����i5S4��(!���sr�*5X���7.#���/j�q�YNA�]���U�v��E�[5EyK�����)�1U74��bd��D|ŵ1���]���iճr�UPئY�[\0Xj(����%��b4m�mS���_�mm�V����YD�e��&�U�H^�- q�����yq9���J���?`�]N2e��=��u�hҼ�JA���]P����M��;>4��:� �<�M�.~rr�����4j�Zu&�ۤQ���{��h�NG�t0t �:��ODc�dC��6Q@���]/�z�����-�8�������nW���g���YKC8˘�އ��dw��� ��sN���I�g%Z5D:K䑉QF�$�e/�Ñ���W.����OA��VTac���K���g,?��9�n�^�W&�(X��KYt?��Am/�}Q11B'<�1��]p���~�T�m�t��k���$H2�^��D0�r��}��~}{��&laڤ��f�*���������Pn�xb����V�^��\[ul��qQw�����Z���뾻�"n=����Ľ?`���I���j�]er��^�Cs�eR�T�0��h����]Y�6� , ���'Y��yB�.�@���
�u��o�3���؇4�,��L���wQ=;��S2�;*�!ɭ�D�NQ�?9���(�ڪST�(��g�#õ�v�:5z{�>�t5#W�[��f}X
P�@��Bqk[[Nks ֫���q����`��1����,Ho߿�0�Dv��[�@1��b��Iܨ4�6��t���&/�\���z���K^���٩�<
��8oV�x���R��]��u�W�b[3�]aQ6��1���M{�XI	�}Ļ6�� ;����\�.&�Gj���<���@Dt\eeL�Ie��p���8-����V��A�H�,�Ȱ������=��>v�(9TRR��יn����A>�y�u����W�V
� ������6o�ԅ4Xr�٬$tb���y��Z0��t��i�����������زM��,���.�/��6�D���������|��Ne�2����B����*p%�ׄ����8O*svͦ�/HKl)�5w V���Bނ���uuM[��޽�P��+(�+�&��C[�����֞�t�Φ�����
,�E�ք�L�R>j�Z?�?>����:�������K�Z�P��J1جƅ́���m���M��3H�q����I�?���8WP�h�����C*�clzxɘ*��1��u���� ��XVV�7o���5��)�1��/��?K�x4ϖ���<��V����9� �~�Z���mv���|g4}���~"���u?_ߗ�^��K2< �J�T���d⿂6�그�^�
�!�i��

Ớ���ͭB� m!h��~}�.�u"��yt��%�B�Nx\����&@M�O.]�cf�l��	!(h�� !%�k�C�$�XAɺ�y�9'Y�TM�_.�5�7iHf���f=-a�Z_޽?׌�\���W�kH!.TF�F�1�F�j�(:p�m��xuZ���q������
�����2��%���I�WP� \�v|�C�M����3.���		9���|%V��)�*B@@^h��M�m~^�G�<�Y������[,��C0�+@n"��MY�$�Ϭ��G�9�����s�L�F=_uޥu/.yP��-�����z>:��!$z]�ׅj�^ > K�%�>�F��
��S�|��kɃ��M���ad��K/1�:�âDu�n�on�0F{���F��&%K�^i��a�J�Ir� ,����l�S���(Z�|z�IiO���$�F[��p-*Y^~P��m7{~^���f)��X�����oNr���Ub�N�YJ�V���l(�����]8$3Į�� � bݽ��f���񡦥�7�RLQ멱h��{�
�.�qP���l[�ˀ���_�Hޏ����{,0�X6(G=�Ŵ���l�ymLTcv�6��,��˙���y�`�º��u ��Y��S��iZN..�Z:Z`�D3
+**^�[^y)�?a�Z9�	��������`%��$�6}	�)��h�M92-����^��ʴ��4�d_%f�>�Ara�е�#w~�F�	��B�
��v1;l��rH���1�s�^0��D��+�-��F��8�J��h�ài�~�����.��#��ad�~�Q6��O��:��4�Ǥ�k�]� ��>�;S�֓#Vih��9t t��A3�vl�ׅܥ$xx~���9��(ǝ��O�M��I����IfUn�R�� �Ϊ���(r�#��H��v����d{PP�2���M�}��0�~�@c���,9���R�;��	�}"�!��2mS�|���_�'�&�sn��^g0�Q�i���h���e�}*tA��N�u�`ܟ�^Z��7c�S��va/W��T	Ph ��,��v�0ښ	��F)��eb�J�~|_/�e5�.v�{Jd�u:Ql<�"��i�RZ:t��Aɣ�%��\�02�B%�BJllp|:��@=���67�V(���k=\+�&��r�a���$�k���#�G7N� �#%%rZ@�٫1/I>>W��G�ߛ)�\���6X,�ڙ��g��,Y�EMC�����%���.���c�KK�o�}�z�y	���	���a!���T�B^����M��D�m�eNj*�0N��c*q�k�	Mxy�U&�^]����@�T�se��K(�1���1�x���T�7h=1Ԕ��=�Y*��+&[;������v��%" ��h��l I�F=�C`t���D!�]�!�����}������K/��L��b��� � �eJ����ވ�@u��w���-~����l)��&a`�6��i$�ͻ����,ߗ��r��RA�I.Ԙb��eZ���Gm�4�L���
z�0�� -�j� �
wQ�ʶÇ�W���#�[�݉���Z���4��7�qֶ�����8�\�b]m���i����@%eݝ��(�UF��A5fm����Oݍ�ٽu���-�l.�hj+-���\a���ѫ��}(^Zj�'������A�b��?	u�)�s�d����6Pe��g����Iq�"¯_�m��<=� ����:����x���CΈ��V�����(�m�P���&F���*4U ��Ҿ��TUUE��v�hd��CݍXU���
�f�I�8�����M���4ť*���Y�܄\��B:Y@���G�� ?s���L�?�X��RHhi�@ĕ���TyF\�/��Z�I� �Qf���7���47��t77#��~΁�>�~b���D�������Ww��"��!��ʉ���Nʾ~%�*n�{>�0;��C� ����YZaA.����8��E~=/�����GFF�Jzaf,�h[�נ݆W�MG@'�+�R6޺i��Ky�6v%ͩG"5���_��!��z�l�ڽ'���a��q34s��o�������qT�P���TFM�����M7V����W��׼,-uǎ<h�ݳ�=�(P�Z����eB���$\�7`m)K��tO-��`�Od��X��$
�] :�W�-n��c�c��ݫ�,RS0��F(B�qtl�GN�.Du��LB^S)q��`.+%3)���c�hT��P������ge�|��J��L RԚ�EKlS��3tSSSs����U�5.AA�C9���0;>��bԥ.�E��!�S3T�%2z�D��;=��<Ř������܏v��3��H}\x3"֤��m�n�n����7�J�_]�����0��d��c�s2������,�F�PK�8���2)����?���Y�3�萳t�L�f�"Ham1�P��7,�ۥ6ܺQ7���9mR�����bS�a�����-�ȟ�#���Hº���N�WOrKQ��w�: �j�ųȯ�{��<��Mש����״&.�5z�l��K�׏���Q�H��G)��)��f�d&_����\]�[�t�X+���R��Ȓ��2�_Q���PC�ǚ�F����{;nz��G�J�Ê���u�_�4AU*1iyq�a�@��Ta�`����`r�sx���A��R[���T��tvz��x�%Њ��v���9��!"�F���8���>��&���}���h÷n��iO��P<����A�����@"��!ƴ��>;QȒ;�%�/���;g{�ݸH�!Rw�>J�N�<�FPsN���*|�H������(�L�M���	υS��.� 9�,ҽ%5��ͥ�i���)(0�YE���ݻ����]�Nk�*�L������FW����Pd��b�-V	��bsxD�0�~N#�)e��i/�jI���P��^I!#;����8wsn�fgg3}��_A9��N-��S�l��u������	P� į���������4�  �PK�&��jU]M-y��.���ܨ�T��]��3w��ͱ�&eCcJ^��������^A�Iu�al���!���� S�N��s �Rr�'9���hպ�u�v�r�n���Oܴ��[��¸ğ�@	�<��q&�҃��e)�k����(t���y_�]W�t^���{�n�r��U-.斜��6ض�z�d<N����e+�."]]�U��Ҁ��ZyEP���Fxz1ꨋ�9C��5'/A:�`�gr$��^m;�k���Rlw����*d�ЦA3�u^?�ym�o6L+��:�*���;�6�clq�֯_<�I$~d
�C5k�.1���$ �5\"��X���Jz�	�JJz���'A����:G/	;Uy�<h��Xp*����x���z]�sYu���]r����	�,Dq�^6�9���0���u�4�w��*X_>O9�&|L$/� ���Qh]r��bm���\E���|0v)_[[{t�/~�v������w��������K�*�DgM��M[�Dt������Xþ��Љ��3�7FM�SS����ᦏ���\}ɫ�D�sۛ����4ৈ�s^��6jp&����o�5�4���)u��X]2H���(��0�����i�����w|)j�.�@ˣ�z^V�Z@�[�s٩"o��<�_/ ���3���wJ�}��{���p����[NT	�c�
�g� �>�֟�����޷�dR�!9��غ�9\.��1��)|,I)���c ߁���h�I�`�|��<����n�,"Wi���}�q�Ag�X�0&��O����RG)���졹������ɶj�5�����әp+�_V�@B�m�&I��'a.T�ot���'�������(^ �k>|x�5��ȯ_��΀��Z�6�����*��T�%;?*wu;?6�5X����+�公*�.�w/�NMM������PGQ:���K)�n�w�o��D��@�<Z]��8GÅn�4����{���u^�@<�$k��xDLY��H�ˤ�W��76.HII)��D��)t�Lm+(00ӱq��z�Cc��#����▨{�)v��>�IQ�XG�O� �W w���za=]����l���� `B�,XNN�ፍ3�+�^[�mm����� 5���4��q]���V��;L�|(l)�Z�$C��=tyR�c虂��Uxn?~♜ @@ñ��]�&x�R��>Z�\�����Gu��WK��k��s�G��OM=���ݱH賴��}Ʋ$��y�w�T�1�K}_1:9p��2ь�R�G|��ܾ>��z��f9�G���,�׮]��#{2�!���+,\٬$�����bbzO�����f��ʄ���o�j��Z]��)]�c��y��*���[��5u�⫚���&2iJJJj���� jH)���)�Cx��t�A}J|�S�ĨB�5�*�&�.�,ӞR�i��M)-�<;�6Ԁ�p��� w�N�#�yR�a��v(�P�L��`/Lgڼ�����т�6�b=tNY��߫/��^�kx��;i���^C���.�����O�'|)��54����� Gq���X�0��T�� ^(,�F�w�:���[60>�����Z�#��L�Lt|~~>~�b��:t恺٩+q����oz:��	֝N�9{�U;�)@~cO�k"��5P(�@�tSp9W�	�E$tU̢��������R;Urguh���w��=.�� �~H�N���RF��*�L���V����=#����\1/�m`��	��{X��Z�'�M�3gM�bm7�*�+�x�F_w����{����J�����#�=M�Xr�s�R]�b���烙MY���Dt�p��E����c3N�
� h��I���-�^���&�ĩ��V�INd��-�Ւ�L���p�;!!����B<ِc\%+]�X�!T�F�d�����/]ʶ�G�N�>�Ú�*c&��#(Gs������ǧ�v--31l��L<ij��A&�Œpk��uВ����aR��5A5�2��ؐ��2l�!� �VX/�@VVV ����H,Ɉ7�w��_�y�e�4h'mnp:���KHT!��3��ط0ڢ E�sv���[gS�~�@���n��~t��*�=zM�����	"Ү�A�!�����E�ZZ���("
j�?��
|n�|u���&���U�c��+ Km�`�_5�����L�~(���+J�vo9��oY�O�4W�.IP��T�0�ң�d[|����P�V���`Ogܤ�aoб�J���4�. L�	��E���}UFB}�7�C,_R�yg�w�����anWyE���sss���RA���K� %���Kt44GF�'O6^��*:H
������7��\ �<�$�3�#�ohtTg ������T���`����d�;�7<�_p�k�*��Y���<��
'�u d�	�<�8�U���C�o��;8��nw`V��͌P`�B�{��7�P|P�ӵ�(W����m�>kR���<����]�&:�p�( ��Q2´�o޼%B�zy��!��H���湭"��ḏu��;��F�PSv~�66��z�Ӌ������(L���{��G'�Jq:u|½�Wo��mV�\)��O�����upp��z蜴UԵ�kdd���ll@(P\�k�R� a���p�}�JP�~��|P�k�fTL��mU�LV Y�,�&GӞ���c	<5C�i�g7��@'�|]Ԋ���J�"��h{e��h{��_��c-�3@pLR����~�_��5�"��B"�`}k�>�/m�r�W/BA�����u�X���2wƛ�2�7�B='�c��4�>��������f��������bu��D�䉛�k�"����RR�w������}ܔ��
nm������w���4�y�뷿�OH���}�
��(�0-�!^�Ͼ��,rt�qe  L���:��T�ϓt���Y�����W�s�	����O�-nu��YW��㗉�'�Uno�k��BS+�ٱ�������n�H�C�Mhr�s�)aD�$����	:{�y�T����ח����r��H����jWWW�C��^$/TI�]dR�V�0^���ݔA��.�C.�^��#�����(�����OO���R�Z7�Xv� 햟��j�FFP�Hʬ�tQx���������B�ί��<��0�#'��N�����R���A�<a��ˈ_� ����̌z�R��ޟ�����m����_��ʭ\ֺ�IK���[[rY��;�����w+�]h	��0�sm/�_$t�:IOCÞ�Ӗ��֐݃F�4`�D���9�xm'8'��t:�����u�R���,�ǉ0(?��ŏѵ&�#5���ם�����yM?ҫ4��?i��S��UUU�DDD$������qݾ|����S\X�S��E���	4hƜww轹	��N����˘4�s�=[y9晿.Z�UR���YI~C'��D���IY�����z�<�W{]�Q}���.3�'��#P��R��X���>��[pY���kh���&W[Z�q��?�Pow�}��f��H���u�89��ۘ'��c��Qr��С��sH�)��X@o;<S堼:>ɒ��x���N�#�O�X#%.�vrr�4}�[J�Iy&]SS#��Ύ4��p���]c;<rT������-&�ئ@��H��:�s੮9^c��)ո�,��к+A�MrvVN	��杒A���ec�r\��A��0Iӫ16�4�`���K|8]��o��X�5�V��RG)�=��	����4:1�oqu��G�� c"55��C��O�%�~�Ee�<4����J�����g�w�	JLk&~d���Dia��@�F:L�I<��6D{|�r+�N��+[̕�:��@A�y(��xz�ǵ��ǯ`0l�J:���ccV�sdR�<��|��#��of��_xh��&�1�Q>�k5!	�U\��〓P��N�v����-=����3�E�Q5�?k$X_�Ծ{�f�&�-P#�����ӎ;rT�z�� S��f��:Q���}��?�����y o'z����]bbbi�,
%�"qWB@@��t������q��ڵ?���]�����t�z�f^���o�7u~�#�![-pX�����>��0[Vb�鈨����|�6I^�g}ZF����^3�X�'%���%?���@;�Z&��%%�<�y"V��!���F -�-���'�#Y&���q�t5�=_֠��̌��k�tb�ٌF�r��K�p���8��Fbq�kpڲkc�KO2��n�����;��1WR^�b�s����s~~~�,4Q��6�k�@%�IB9�Gջ����e��:�΃ާ�&HO.���
ї��,�O�Qq}�Q�磞��n���k�o�v-�Wb�4���鎂���5c��Ҭf���Sw3 ڮ�9 �	�r8���+J�t����������?���51����<.��T�hc�25��w����rp*kR(� _��	�L�;R3�k�ɫ�u��g��22U߳���*)�L �����a+F��~Cߦ�\c�D�~�5CC�?j�!5'�>��@背�{�Ne������_�:�;����jIQQQJ۞!�^�1�`P����?yʡ�!��C���ˤ�66f(�������'���75�A���Rj���k��>ibk
���%�3SO�:���X�dni�	���K�=@�n4ʃ8���M��}ZM��t�}[)�Qک���:��"�V�S (��q&x�h����<�Ǳa�u�\������m��lQ ��}�!e�*�+�5U�$�Ӳeee�5d�IE��RW_J��1��F�`�y�_p؊U�o���T�o�I��S �-���� MM�>-�%��gQ&
^7  �6 N�Q�m�l���?���hdoFS��la����|m�&(����h�\$�'\!O~
��gąν_�<\kG�4�f˲ǣ8A�cc��~�G�\��֊YF���7�Ʉw4��΋���?���w+��r��;��=RXmI��ygP���n�PJ�uyttoM�/��[��Nw��z͸:<:.3�@�f'�� ,���\��?g��0݂�Knok� 0 ��(���D��(/�Bל""��G�0|o�S&�L��n H�x��6�]�]�D��K��O6��/	���d�bT���j�~���B�&�`dIP7�yID^������8��B"��)��|!�!�6�Z���E�����	?�y�ڹ����殮��3bOZ�x%�O'�܄�4dW����8��N�MMM&ו��2�,7�����׍��/�O�6�!�?{�U�Ӎ����13���������Q���D���PJ��:4jbi���N:�9��w�9��$Y5n$�{ʱ2�r @�4����g�zmx�[r���iA��y��fb+�
��)��[�Qr����c�o�j_Ix�ɐ�� ��t)���ߘ�� ���q�k���
X&b�V(�q<(xUQ��H+\�����\{Й�;+�󕦤����,���]��}�|иA~���
9���dJv��lbb�����j>5����d�mP����󌗉�|M%8�9[5U��������M�O�c��P������mh��  ����w��TѺ�������7�/���3Õdߩ)�X3��\K������+���S�h�g�H�������}v�=�:,���i�{Ӣ=��VewR����E�'�V����P��t��t�r�Ó�!��c�۝A�e����#S�- ���쉃z��kSR��īL��# &�a�&�I=����G��$�1YA�U��X�Z1	�R��y��JN��[���p�-�C�����Q
S濉w�D�٦�{.�C��o�q��P3Oyߴ�|����L�uF4����ޕdB�9:���b�8����"�%۵�����03{*?�vm�@�ę���2^s��D���p�LBs{�qZ�Գ��񍍍����[��|o�/�lw��M�5]_q���O�U�cjr]V�F_�x��2�SL���oZЛ9`�<$�BE�^�z�y��ʄ7�F�Z�'U�S\�*l���9�J��R�s��6ڒ0�����c�F"n=�"��;2����_��i$ҡl���k�-<���tAP����R���Iܽ
C?F"�9����A���snnn�?,b��%܀I��1N?@
���@z��E"d��ii���LPt��{��3V��>㓚�\��Y<��^�U q����.0�:���$��	���r�|�ݹZS8
�P�3c���_���Ȥc/{xxԮ��Uk��r����py6����U~�@2���]�ƌz�W:(,��TO6��sۻ�T�a��>�z�y< ULl���*�3��0\ɢ�����-��@"`�-�y`cRkp�1�Y�4la[ZeÜ�IhS���'_ښ�R�+t� h�S!n���#',f��߸�MGn��>Z�YY��k	�t(rd�q~]��A;\�=\�_��<�%��-`��KD��)s�Y}���8F������������;���?xˍ�O���j�C�R"����R߼�:�H���`��w�}�p�X��%�s�m~�h �h[U(aǳ���V�U8���L	?��$^��C�[�a�J�V�'*�~�͓��0b3��&Cr�m�ڐ=T#St?� v�^����#�0)YY�*D��ڀ=�?go7ra�Їԅ/p�����ek�ExH2hMڸ}���{�Y���R�d3o���OC�sG\>o8ס�Tt���6@)#
�j��"x:�pd�t�Y����V�L�J�!�O��}�Mf2m,��U�%:�II�8�7m��Њ
������[{{��=CjU�Ȃ��e>��t��j�y�{������_ԢG�5yZ��жR��IIA@dTR�7 &;�9�Y�1�� �¸�o炤��������)�s�M_)�B��M�p_#2rq$����ȗ�f�_%�b���#�����dq����s�!�B�_A���&���-_v���;J����s�
��r�?��6E��?nA�|xf��U$5+���$��Z����W�o�B	��[,<b��ҙ#F_u��"dX�F�Lu�&L�UiSE�-���хF���V�li����7r���_4���B� N�����z��A�����W��a8u�-4�3��30M{ذQ%�b�J��p�"H1?0��9��r\��k-x��	S�yo��=E�}��_X���Mq�A�ia�ez��%+�/a.%m�W���({���0�[ܤnf���w�I�W����I�����f  v6�e��o-�I�S�g����^H�HBw�j�?)v�l޼G����$DN��7�}�p��K囬����sk��u�H�"�| ��?�|���U�PD"�ޤxi�ono��$a���N��E�	������C7�Xqi�.��0���>A3��y���B��_MNR?�WV=���{�F}�N���9�~"�+@���<}Dw�iz����܇
�9���>ZT�ԓ�8`I�~�d�8ڨ?���I��MMq��#X6�R��K�3+<(W�I<�a���#��o�!a��X�Jbŗ��h�ݚ�3�֨��6j��TZ�ӡ`v��eE�_I��N(��"yA@��*�}��G�h��~��E���D4"
`��m�FN�C�Fׂb��ֶs��ε��ʞ�.J^`WN���9M�+�eC�j޽< տ]"�i�:->Z�r�끪�����d��vs���5"""1�u1��ML{����.��K�c9M�Щ�EG��Jы��P=65��z��AAo�ϥ�D.����w�R�q�# �C��]�����V«o`���;�(�8w�
~b��K6�$(�%.ҧ�n8�,r�y�F����b�)oVX]�e��wO9��J[_K�|�U�u����Y8;0/E�X0�I� '���X���������V�g;_�^"!����c����E��[�~~��֡�m��M㘦���tY�|z?9P,ֱ�tK�="2��K�0Ƞ���U=��1+�9^9�w)q����p!�����VhP���%�B�r�Ҡ���P�vT{ �P"/����o^���R�l�ɮ��:[������t�Ö�'(ׯuE([C��'�Sь±��*���Fq���X�ߝV�P����N���\I���MJ�G�݋MIs�q�L�Z�+Ѫ�Y���?��Ȅ�]D,"��M��[����Ƞ��� ����Ѷ���#��:�s������z�?V!�����FA�(l��u"]�z]���id�:��BC�\~/7�J|V-Њ�1+��p���������Ty����|��Ifb����4����X� � ����Ŝis����`Ͻ�-N�T�\V��l���~�lH��b�$5�����B�0~�L��+x���>��|�	hc����ٿ�0�����?L]w �o�?H�"e�
e���������u�Z$��"��ޛ�	�{�co�w?F������<�}_���>�纟�y�������B N ��0?�2A��:�A[j2I)E��c��!	y�䅬OJ�r݅�9+#eA����x�bI�[�ۇZE��V]\L�����!y��ȱ����/�0Cq�n��ϿZa��sS�V���i� ��(�����D�Z���T�I2H������J���ӊԩ�7�XZEj�O�N���%9�"�i(>�Y�>�&}w�Vc��c���ʫ����G��lm=qq)I=����F�J�X�?�7
�Zpl�U�����8?�U_�{W��'�D� ��.�h�4�A��[rW�v�"�<��R�55池��ۂ9��`z76uy������pb��Q�?������f=ͥ�t��Fp2U�E�������ra�ΠW5�z�����cV���W���"n��%I�A�G��-�N۾���%���|��g���ĒB���\���u�P��l.�Vc$=�
�3�� 2尨H��d�u���Vdi�w��9^�!����p�nYW��g�a�c�E��E����N�o�y���>6����aOq�Q�U���S�p�����R�K�&Z���K�N��rw��ݛ�6�/��ι�}@�r wKd�SU�����	�ˡs�{s�%���V����\����}��⢓0�mq�� �;��4bill�3*�%��/�];]d̹�z��_�6��;h���ϱF�����kV��:l��:�^b���1�'m��INX��3;>��}���'���N�f,(�P�������ߠ��|���oJ���k��e#N�.�����#�����>p�����F�)���:Ar���:�B7QL���g���)@%���N*~�����#f�����Z�&���Z�����S!EMi_���V:��#��Ag�*��l�*m�Qz:��Rݲ��?ǀ��Q�>��KE;��ay�S����_�����W��R��iR�}�?2�o,)��xa��Q~�������+z���,��	��U����f_<ߝ��J]��+X�.i���BEĤi��<�d�ykng�;�2��ZGV8A?ft���p/5��oo��ǲ�U'������s��q�n%�wwu�v�׌C�)��wZ�1��H��E1Sc˿L���"G�1,.,����mF�?�{Z\X0�X3��9\�p�W7a�Լ@/Ƕ��M'��.�|ys<��<F:�>sx�$���0��W��l�1��|Q��#���0�$m����u�X�ګ�)K���-���M�>�Yl��"�����m49{9�^�s��-�r�t��s���R�o_<ӊ��D���a�G����Z��>��S�����$��%a�����K�
4�Y ��~���hG���=� �Dٳ=�'����7n܉e�*-5�{c��I1���|����)ނw��5u�Eh�-/{u���� 3��{��9�H]/��Hmm����Oyo|0�ߤx/u|�rxq���UQX�h@c��������[m�:�_TI�>����l���H�s9V��0J��vN��J��3��O�U�Dd�]�u>��c� �Cq��b�{y�����+R@�8�oY�`&�٫� <��b ;�:�U���=�'�k�}��`ɱF�PS/2/�ݺ�<�����aX:���Q��vdU��z��p�CܡG�ŝ?sx��㎖��Mu�Ń�� ���(����z+7_����(��v5[[�����3��K�Ci���1�_XAO�R�������j�^�[��8�!i#h�*��A͒:[�����������\�e�ɷ�̈́�u��|�߽#�d=Y~��Q��q�m�퍌 :d�����&�ci��lb7�U��V�A���%l�$�-�����q����z|���:6��y�<�H�'C���m�l��=d�ª�D�c��KQ�����4r,m��	Y�@�t"+���h�2�����.�0:����~~8-�^�`�Q7�'z�_srڱ.>h�#X��"m�q�;ֲ~K�Z��t�,� �ǹ&2,�����\=�U����L���i����R�.����ݴs,�2��K�lw�˕ɽwܫK�71�&����n�O��$��	��)?�*�L4��HU�a@�P�Ő�8�u����?�}o���[���I4FA��
���z���d�uCܼ���H,�hr_#�����m��bF�o֓}i+7��st0�;��kk%&׳�C��х��J׊� #��S�{�[�=�RI:)����ʊ��5�FS�\�e����q縀�{`���>�Y��U��vS���){izs�,[��~����Um.o���~>;�T[���۷ɉ��w��ߗIWN,�����h��9�Gb���O�E]x翕�(݉H6K��'w�wF�k�����.E�|�0t޳?���>v:�'�f��?0j��o��7��f�z>�=ꖧ bk<09����AN�x|�&,���Nd����'�����<��K���-�4��)�	�W�g��'آ���쿲/�͞O����c���\J��9��B�Ky_1����H�����������:��@� �l�<Z���P�@��qA�`T��"���Ԍ�dVUv����P��Uzn�9�UzN��ÿ��\E�0�v9��D.�,
����Ӡֻx�w|ܠpHG<1]���8l�35s���x��������h2�O6e3�خW�p��'|�{��tll�k��B�w�7���[3�w:K�u,p��|������>TV&�;�����:w��j��Zwi�)�*x�X�\x~8L+E֐���MP
֜����ݫ�\=<�������?��A~���@o}}�F�G��(���D���
R�\���9�+֞p�+i�T!C��I�N�<U-]ɫxM�+������i	6y����Z�N���:��G���_�:¥W.�V����:Q{��1�@%w��%ӾC��o�|[x�0U�p��]�P#���l�bDDD[�ws��X�\*�*P���FFFzg��
�j�x�zOq�b/8|]������t�.�CK�b�VI<�&��0�G���<0_�T��έOn}�����B���V��3��EΔ/x�b����bxr����ҿ�<�ĒȮ������Ci��l�˰'w�B)�GG��]��������[�3w��wv�k�R��'�lj �yf�K��dp=�W
~n��ZhYCS�*E2�j��C��M7Й�M|]ǀ��WB\�7"J���}�)�]VJ�ӣo�xq@�G�d��`}�����N���I���iV`�ul�K�r�޶׺ �j�vi��o�ָ�o���2^|����[ZE��������3���Z���� ��0��r�"��LR�<�	�^u��ષpj�-Y���lfث�� �9��ڎ��`��>�ۮ��ԶuU��^�����$��:9�U�>t��ڏVn��%���Q^w��#��!.�(��z���	%�(f��ş�v�g6�P��x%T��v���kZX�}+�P��M�NP��M[b���'�(Ӿ%*�ϿJDd��ibec��]#���Tg8���n~�=�v\���x�{@�W����
��o A�3�(�_��g�ݫ�B���LbJd|�-��vt��距�<��xb]~|����e�����\���TogѦ3��Ȇ�x�Ig����dC��ً����姃�>�6��Jk2��� H�և?��9��.o��]C���"�鿭؄x��*�7\i�w^R��AG+�p>U!��̱������D�!���X^�P���._�?�2��V�-x�%2;��5}������ݓ��5���b�E+�E���hb�Ϛ^NKKВ���f\0}��6�g��2:��2)_ZMu�5�� �)�QG(A�ŧ�(k��P��H
���o)�*�Q'�����U?���������|�׆v����CX-�
<ݎ�^��3{S<:�R��ȳW]s�U�u�5U�^���=���ݜJ��3$q{ 7�*�,,�ο���&�7����<��Yu[��gG��2\��~�vU����Y��ӻ_ϳ����(������+%�G�[����e�fj�\�{i�+�E����{��wm�����~jjj3=��pq3�_E^����M�G�>ۢ` jW���U��Z�sasw� �u�lP��B���	�RW�;��΀����`�:	�����M�3�X)R��%�	$�Q}4�e�_�-�*ɫ��,f��w?���ԋ99�^�.���b�	`�Kߦ�B�Q?ֽOI�u�ڿT5s#|���}�{�O��G	`�v�: ���;y&ѶU�xcF����vwJj�]+t�� � l��v��hy���Q M�<j���*
q�]��F�Ѹ�,���=���WVV�:�˟���Dp�ͥZm�8P��5>ma����>3�A���#S�����^��h��D-��2�<0�C�^a��C�{�JF��`P��X�M�:)�&!�D��pM�q��_kk�Q̰˕�!K��˜��m�x|t@��'��(�$^�ځu��ۇ��Ź-1�����1U+�$�!�����6lP��g�l.�=vY��}�k2ds�=�حX�J�{��L�ׇ%>�
��>�BoSnpͶ���)1"���YT��<$J#�z��bуy��px�s�j`1Dm(U3.��rP�"��ݔ�nj#G�aI���e���/�c���z&C��C_҆
�-uL@ُ��\{K�~:|�C��-�X�N�S��˓�ޏm]V:�9l�=#OAI����+
���谪�����x��&�D\��ѭ,���V�a���C�Zk3 ���r���s�xǖ*XF%r&Dʎ��S��@r߇>�[���	<g|�]���r�A�QB�k&ѷ������WRM޽P�w��=��}w����>mGk#�k|�}��S:��؋u(�T���;���P�f	N
����orM]���Cx4وE�Wk�7l�1�yz��~��p5|i)�E�O\�CiX�OO������#�,#ܓm�U��I��A��,�? n�^+[Ά%�����,�����($1ٶqП ';{�z�(g4��,�Y���F���"mA�RHnF��񍍍2PB��+�xG-��㞈P�@�>L��P�:Q��I�7�_����W�,��s��ӍԶ>פ��'��<���iޑ��ɘr���lk�bֹ�f�9uy�kS�{���xMM_v{��ѝxt�kH�m�*�o�����p��?��2�lŐ��9���bKw�Wd�~Q�-r�x7{w[�n"�����\��vY��5{�Cȑ#�����~�_豰��1�h�@[�%����'�ƍ�^%���5T�Γ~��Y���E)�T�G��qJ����8�\)���'��d%<��dO�Z��ѡ�hh��������_���
?�8� �/M�&���23��*=ѻ|�~	�R	}~�άC�����{�6��p��s��U_��� ,�8��	 �,m�[XنN� C�xJ%�x�cϤC�xarR
8D��?��YZY4	���-�]�BYl-���k�$^<~:�M/�0�5�PDإ��e"t��s�Pz��S��&\��@���~�WYIC�̂�a�]eP3���?��{7�<Ѻ����). �>�#���+A65|ɜ�
L�[���7��Ɨ��3s�|�ʼ"Bl�X��:��Ӆ��,�A������������oҾ�UX15�H�"��uOO&���J󤨴�*3���و_U�Ề��� .����=�6�@-�Jш{�&��R��|ؔxД@ {�ǒg�#�9j3.���p;|IP���R�eS�+��p�4`���{�����0IC�V�N�D���H�>(�����iR*�9,��n����H8Ȓzp��n8��$��[�Y"�/^y?h��)�D����k$(7҇����$`�W=f�͎�k�x;���NΠ(t�3�Ƞ���;�8f�{3Q�������_�<��NW��zU1,w2C�f��������swM���~NX�?ܔ� �u���؎�\;Z]�f� Un9+;{L[�@P�"�P�m ��G�|ŗ�ķ��Fp2k�3]ݑ��-�ƂvqL�����n}6|�ݚ���~��IJ
��DӮMY��N��ϟF<7[��8 �j^m��:��n�ƌ�ݾ�bm�h&H�����W�b��d���1t5��
�u���._I�Y|4��A(vC"����ȥ.8�q|��[�HӐϾ26������Q��\��th�2^ޛ�>����W]{r�2�=u�Tv?'<��XJ4���`~�H`
�����<$�`�,�iJW�W���b��3*?D\ځ>{Se\1����� x��G �gq�'W}S8Kx�哙�4��&$q�����<��J���a@�cl �	0��8�������W zEQ��Hu*%x�fs����VJ8��r�9�;�S�,שO��7��o�#�4 �cO:{�^a!��r�KF�m1�?1�5y*|(0Z����9��n���.*��r�̠�A������:���qT	)�'�<����0K g+�s�p�|��3���`dPE����i�.���(١J�u�1	�:`jf�hQY�u %@�	�V�y��r���}� �m�B�abr�9���K���Wj�)�����*^b֢X���W�6U�,����
��"�=�T��m�!�<�KI� 5 ��98n]�)}T���d�W�2^�KxA�|ff��	d��X����bdz;��T�����k�~U��b83��F����V��)�]$#{"�QE�)�����h��'�\iDف�i�:@`�T]�u͇b�{�˰�������{{MLR�7#�A'���m`d$�,ыpw�EƵ�p��fO���o�%�&�� \�\E���s!��bO�3eX��0�*�p��s2A.|�|u����I�G+,�!:!��R���D�D�t���v�\ms��RG�Ē��б��`1��	�o�h��w��g��v�
?Nb���@~C�	>h�3��җ����K���v��=`%�F�@������/����NáYy���^`9:��WhC9�*W���~AL��'+\$ Ё�>Y�9=$��㸪7�e�JK��>\t�:�6�/��p�7!_������<����s@A�$
Wr ��Q]��)��I����u�.�����@�����s
�o���_Ck⁍�х����ʿĢ����vkpW�W����V�߈v�<[9���_/��U�K�5)�q%̊|�Q�{��R��ng�7 G�Ұ�ڟ`;����d|��ĹuH�umT�y�Eؙ";V~��(?�^p���[�����R<����%������'c��C��s�=�K��~K붠���&�TU��~�X)v2`>�T�Ar�6�Ü��>k�����Ү���]�ȓ1;L!W��yزǾtF�O���V$��5���	��Ȩ(J��J�1��Owܫ�={��:�\9������8�k�Ve��h�rG3s���N}������0�jm43�oT&�A��Bo���r�Z8���^۽=�U���G��߿}[*�.����8�ZR+��=�@5��x�z#� 	\����M���b����L٫H��oJ��Ûz������A_�J�R��0\��S9q���tzg1W�~��Suri�o!8�ψ	`2R�$.^��^3���XQ��Sݏ��69'�ݓvE�7f1��4�_ݪ1�xȯ���>pU�=IXa'Ш�z�0���5��`T� �^L���!ШDԫLp@nQKW���(����(��a]U�দV�v
�П�Ӏ�C�˟O��}��Jx@C/)T���Z�����Uw�Z��0��É�� �؃��[j�%�ԟ��l��&�¸ve[L�g�c�_�prq�c[�K&���989�B��j�@�����t	߅���}�~��1G�N@�g� �gz������[�h��!��x!VN|�m����ޔ�u��hPTgT=҄B>��Ʃ��8	AA�����&���w5�H2ivv�zH1���M���555U ���pm���9��W�������S1�	q�`��ga��l��,�uw��
8�@��d6dh�ki?[�h����f�9GM2g�SF#�^�r�}FF��Q���E�_\x454Ƣ	��A����Uq����,���H���쀸����I���,�z���Zw69nv���
�9DY�זA�3�ڟ���a|��X��Ӝ�@���?��S�Cz��|���4z�i�(<����WݍVe����p��Bn\:��m��p7�2L��Te��f.���5j��i�$�h�u�I�ߠ=�������9e�!ڼ���X
k�p"��쏬�W�I0ŨnL���hd�)�?����ax��юL����z��:nB����o<�l��Ms��j57�(�0ɒ^ʅG=f���R�]]]�S�p%P�*�W_��^c�h��<aUfUz���$�� ���<�W��|q��yN�eQPPD���:��YD�U@`��	� v)�8&�N�$E�h���~eZ#y�&�qos��{����2J�t�*}[�7���3O��,�]���g/�	e?彉��)G-Zǈn��
�Ņ���Wɬ��K ����qm�2Rͮk�����յ�r#�E�|1�!@{��@�U�$��ܱ�/�@Qr"�<���]+R��hx������
���Ӥ����4P�}N �4JNՎ���h����D���8q����l��Wн��剛��8�G�HIӕ�Ӟ�솲�CZ�~v�t�*^%҄��s�4���c3��l��K[�`����I�����afgLQ�ҍ����5l+p�����B%��V�4�V��F�4�q�6M�t�+��O�6Oy^Vu����H6Y�D��������9ˤt>�y���b�A�i����2��|ד��m�{��o��ȼ�F&-%�u�9���:y�����h�o�ø���G�$�[V�ҲR��!&�Sh�\P��Bֹ���pB��3m/?�b��j����v�T�t��E��Dt}��5�7��i��}'�y�J����G��p<�'�<����QL�i�cn#���������[��FF!L�	\�>snv"��=5J^�L���&-�.��d��	"BP\�J����X���={i�+�Gl���M��)x@��Fw\w�#��;�
�Ea��nޠ4�Mki[S;�����vGa��ۏ�.�N<W~��_��o�N��@
���,�Q�3أ[�{ȳ~�S/{m��K�b�A��r���N�)�-T���~��b���Ch^�;��;gyo\��祃�%�Q�#��'t����?�Ot���5��~�8b��,S>.���h�K���A�!�a�{��B�-����8�Q���-���K���u����a�vE*�9�8�69=T�YX�M��$���(�MT�K����⶚�/Q���k�ϒ3�Vmn�6L,����V ��G�}·|FtmZ��V�ڋ?����aS��l��3�ڟ���0����*_�_-�r������ae-{�@*�mj���َ;�6�`!�ޛ�w�9a�Z�
���5+��Kf����yh�~����x	�	�L�FI�l>tt�?u���#?�lv�>2@B5��X�d%������Ѕ/�4� ��ɺ�{��:�	dD�W����~�9l��Iz�\���RqS�݇%���Yc,?;<�G ~Ч�:7yU�?_: _b���cM�^���M�!}~�='4���9��o�U��3G�W�C��T$Da<G�˰�z�:E�<^䨬����K��'��#�.pE{$.%�m1	�6��K3x�i��{�$ܡ��)f�o����GzH0>���.��xm��p2f�"� %�ڑ��`�CI���w���˟�I{���1�J��aP�K��m�+LA���l�ڠ�:��}��Ԙ�����ɬ�V�7�r�d#_Q1�I��E���(~�91�AS�u���[����#L��A��-�%�f�������{�-,؜N+����[L�1v���O_���|/��W��.=�ڡ�#�m���@U���Fm�o�d�*��\�UV~�������،�j�n�?W�K����59E�/�6�tt�iQ�1���'��<��`-}���Kb#y&Y�k�b��oY|����#s�_�k�	iVI?u//�ne�4M�
h���SCp
�ĩ�Jl�0��j|'1� ��E��B����U��!��S�B$Z��&�v�w�a��i�.�Mpt�%M>�w��bW���Td �d#���Ϣ��mc�%�	$#G�go)��}��1hm����Ԟ������YvŽ�8M��6�RY�� ��9��&<WsK��d�Y8&|G��5脋���_�/���:Zr,�f�&���y|�$��1@�O��ɤ?	7�[v�i���]%��)�-=�})�U�_ޣ�on~�H%y�Q
��l���ʅ��&uM�����������wRq�bZM3�ts�����ł�[�(p�Kucec��O�+$fg,K.�)���,�b�7���Q��7��t*�ו�s.'��zj�9����s��|���_��r��h�G�E����=/���qN�P�*���!'��!KY=k.N�����>im�+������<q�̇��@7�O����b����@ ���-���FP��![Gk>2���G�+Qf���p;}����ڋ�z�_y\�37�e-��+/��A�)Ӣ�������~8��|�m�{@�츑���`��p��hEv����µ9�SP�6^ar��q�}t�C]^^�n���QLD��_W��^���:*ʬ��<'WO/.f�(�N���� ��ك˩�_��vFG?�2N���y~ �K��ؔV�7���x߶$W��b<W�����:Z�Z�ڔ�9����:�>���3- N�'�W�E�)@������*X -f,`*�����4I\1�%�F�*D�Z)޽+���/��7mJ�͙;��Ԯ����QߚHLk��2B�����jW-o���x���)ۆv|�9C�e"���D��[ 9��y�<r�>��y�FP���}~Ӛ�_���Y�M��/u�f"�ڮ��	�����"MR�����t�D�SS�! \���N���h<q���n8sd.��(��Q�M��g1)_���]��r��!�\�
�]h����h����+�usKK��!��������Q����v��ŭ�Y�b�L���@���%έ��v�X-_z	�ӥ����Zwnu3��+ �N_?*�2[��Bu\��Yo����(	;��B��q$@ hY���׻��(�5WY��`0ڱ�l���PD�x�v���N�{0�d,F����/����b5&���T�DFE�!a�)�"u�{��6�ux��!%2{vi�
i�����2E�t�Zo(w��j-����w��Ķ6�b�W��ԟ�60E64-�Tef��^���c-J'r�0�rz�� 슠 ����2�c��,�
ob��`����E�u��BXS�f(U⎏7��s�c�����Pfs`W�Oe��Z��	��FU؃��v˜*~bZ����'ح�j�f��&~�lP|�8��N��}:FϿ�ng4�I��#ڛ��b|��"������p�`Pl�̻��Am��H>En�����������+���4P�˻�TI�y����=����"���<���-����U�M�Jq�s���-΀��J!�(u��d��u65�;`�������b�
�j��Y�o+]ʮP���p!��R�ւ�_�E ��q��D�~��^�8I<`�{#5$7�LZ%�����Zڔ��/0s�OfUE�G]/H6B#�T�;��}��&�i��g�O#d����-�P��6����[��o@>�w����L�3����Z
�H�"UE3��yT1��q!;�����V�)�iKa� _�g[Bn�J*Ȳ�No�z�����i͇	N��uŌ�T0:��ίQ���}��e+��/ H_b00�y�µ᎖R!�����y�!i��ᜮ��]��&�f&��'|=�o;��[���v!Dd5 �ٖ̍����[�U���:6���"|�Y��W>�ׯ�9��u���---v��%`���|��6�y³:eXR��3���)����I�����z�R��'�	_ngy��S�"UȤ�<��1��g���R��Z�����l��Ͽ��I���^��C�Kbkn����\��1��G ��S�Vއ8�� �:��V�c�#H�F,��<�c�q;`+VY��_�ZĲ��n�SӏY��8����5%��9�E�Z|�͕�:\����/�׏G"
�`Bt�i�鍡o+�Ņ{�O��< �KC``����=�s�C�^��b�o��'��պU͉��?����lY��M�Wٝ��v7J7�"ϒ���y�q/4X���v�`�#Ho�Ǳ$���Q�D���4{r�Fʗ�S��%i�z(M���Nk����ё�����/FGA	%9H�� -��G J�+;='`�U�<�+���?Y��2`��x��}F��t��o�#�1�a��6X���2��}|�99�B���᪼�r�.�e�*7�ׂ,��n�՛�����Č���;Mz��Jk�h����_t"k�<�+�
�[�8��o�HWjƮ���֟�����_#��s��ksD� \SG�>��������e;��<��@�8��8�<#^�Q��M��G�V��I����ނ'��5������v�'{�����|�/�[Q�����������Yv�̞={@@�y�)HT�c�J�� )��L"��\���x�IM>��������6�o��o������L��:؎o�?�M�@�y�B�����d�cH��_Ǘq�����1_�pZ�
`���w�>���;J��7�Ҭ�2��������A�����S-|B�/yb[?�<m�U��Y��'�r��1��?{_���m��Ό�]��e�.��4�GSrx'���'�v�x%�mËN ���?~2�5�������X��y�!*�٣���b[M��ｿH$h�%�m~��?�J|���k��yNr	�Q�����>BS?�ÂǰG��T��g�~Z;(��A��:��B�c�V��uID��W��yp�yO���ڦ�4�1��W����խJ�抔?�	(E��L�g<sVP)�D��S�r;�ؾe�����g�5�Y�V�9�egGQ�>5z�Ay��HT�QW�j��<$�E���"5?=;p��ݔ�"��%���\J/�����_�h?Bs����
M�Xoſ4�ѝ�Ӝ��ڪ9J+����_�jg..砬�~gi����<O�����x�������X�\�
j6�V������,�K�9=�Y)ѽ���W .3���RV�s�41�w�1�0E�x�?������t�y`�h�t%{�������~��~P!o(������Y�ҜPR� ]������_I�X�q��Q@2'������?�2���R�P�}�c���NN�ْs8���ׯ.,������v�ќ7�N2��M?@�?���&H	�,��٠�*X.��U�	���		��\��&�����,��(�Z��m
��f��P�d��{avRC>}�劋��`�;�o��%@�@�=�v�=�_?��k����E31���%��/��J7Pm���5��2rY��|!H�����kU?=��u�gfLүa�\EC:́�d��*i7-�Q�_��=+j�Qj�*+�e�M����M��	�A��y�g�k��@�k��~ D�(K��KL'�EX�"�;#��QC+��q���c�J z��}���w|����. *��U�?�S+���m�� �a���� ��,��=�� i�έ75睮�C��[��/Q���LOO���h��:��b��	���c�� 5�g�5�5��g��]�淐G�)�gg>]f��e�)8��1�O��PnL��:�l���5<����]���l�G��=��pe�ha��~��<��`$
��F��c�6�?��@�#@��5�Qg^��B���7����9�Gp�q���߭#i*I��͜W��4K}�Ӭ�e�#jw�L�����s?
��$b�#bWڭ��l�l�����Ȣ��|$�r`�2ͿBЭʚ]J,�Y�zM3ѿ?ބ�D.�&��wi���h�.o�/v��+;ލ(�N���X��R�t՚�ݨS�Y紜�������E�[U]�>��(]zn������ Hy=����=�(��Km@�)~����B  ��M������hdd�TFz�� }o2
���w Nbn�T�2-���mC����;rHJ�����+%�	�2}��<i�`��C�t�7��\O������+���d;�?�N@��	%vӿ?�l A�i���^Te���wә}���^�{E��$q߳$<���A�'��n����� ����|kо�J>z�ݛ����V�$�A�҇�ӹ�:-k��<�� ����힍S�;o��7})M�J��5�v��'�k���4���' |Ŷ����wV���e����&J9�z:W���3|B!C��%W�����c~!��x����LD�8ڀ��H�B} y�Z�~S�L���T��� =-Aa{
|��M�ԕ���B���~�Y2�H��O�� ��4��a O��S�v+E�i!�����Oy�����{�����l��*%�K%�Hs2���;jÇ#z��3�5}9� =�S����Ԙq�wB��e6����b
�`�?�ޘO	m�3B�1�@�+��rr�W�;#1�8�:H	W%9V+֪]'�@�o�mЊ����e�� t�+���9�NɎt�ջ\29��v��#�r���3�vÚB�c�#(���>:����yU� �(�VVVY��(�S�D-�ۆ� ��G �e�;�(PQ�hS�f��K>P[ŕzaS���%]3�L�?�%�b3j`�X	G[���0�w #n{^�_B�s�� �x�aWJ��c6���.�C��v(�(+L�qx�h�đk%�v�|�
�A"�k8���ޱ�oV%ܔͳ�ې�Aw��(deg7B�\���ux
^����i&50-.@�쮌��JM�
'x�n�򾯡�|�v�,Y�6����3�Z2����:����FA��H@W�8i��a&u��^xjJ	4��ehV3R`��&�{V�فʞS�2�
e��E��%Y^̩�d[�-��%u�ē	�}}���&�t�y#p5������`=6E��$���x��	b�O���6�{�=��M<��ˏ�a���_���6��"��
�BB�'�j�*��i��cD��_T$��U��c&��`�*�Fo�7�Y��|3MN'Y��������P����prys�	�8��Խ�QP�ޯ�rs��yقz��oP����G�1��yݶ$����M�J��+~�������#1~�KS��/�98RC�6�;� �=w�TY|'���H8>-�]��v���RЈ��4�hQ�%���]�s7z�����cy�`b�i�p,]�pA����l�D�aVN2��`�M)�>n����;,ymF�\�,��10�@W1��zJ-q�)���ݙ�߬�h�Av4����Eԃ�o�!����SL�\��ls��UCο��l_^�~�l�8؆W�}���� T�y���u�)�`���6?<�)������ �ٻ=��3;�7@�����eu��Ln�'qOz�DC��+��+>w��E�,>���O�*L�{wz��P@�P<��"�&R[��q���uAB/�:!W���wc��6[�ڐ�XT���֌��$����/C�]�v���hhcA�G�)H)V)��kщ?$�"T�H�#�����3\>�+;�����^�-��7V{aTe*WL�n�ڃ^��_&ڲ���t�&� 9!�3W�zo
�����/��'yȘ�1�Ml_ll,?�����7�ӊ������i���f��~G�/���j��JC ��N�F���B7�c�E�E9^���O�JT*����n*��؜Au2���e֢aɏQ�^�jv�z.@��)@E���NUG�C�HgN��ʈ�3�3�}7�[����A�Y��{|��̍Y?~��W��	��}G �~�J֖���W�<U�4�8AR���� �/ ��Z��t�͈?֚c��K��2)��~N�r�pQQ��+�^^s��_�dK���6竏���iNֽP��ۆ!M�4�d�5�]t���B+b��������۫i/LHi��Q�{���ǡ$��U�Q�)��C��c��ߦ�b���G���9���㍔��-}2i���,��9�#�n�(cM�=�A�\bkq�	�[��)vu��b�=GB]�����>\3���'�Q�!��)k70'���(ȹtg��bpd�'�j���v�V�M��䅵;�rw7�g+"c}��N.�B^&�%L�\]IFKE��OL�um�Յ��4�H��?G�Z�c+�ut���[�*�u{�~sۚ����_���t&>���kj�#yS��>}.V�}�
��V�Ì�u�eA��V��e��'��|�/68$�^�R��d�oꯉ�}�iW�C�-w=�ܪd_c��kf	n��3w���VM�sz:�����-�X�W�Љ|_qMs��_?pU���	O�_����rGv�jQ��z�� Q��xu�k��5����W+��W��y��/ζ�Sgeee��*���|�J	���6]:����5ve���E���p/~����KGKK�]���@��3U�/_��
��|��Y��o=�ٝx�|n�p�R�ѧD��݃¶���	4�MW;l�col�!{@qqq�����JT�Z<]�ݟlv�J�4��0�ӊ&)%E�ű�h���x�X����S��x�l�/О�6�C�X;x\Kp��<�zE>���Cb!�m������ !��o	�M�:�'�~�����������M�>}
B�;B���OG��o�{��ӵ��d�˰}�O�z aF�豮��%I�k|���^H�����!d�!T�ԮE�g���z�����Ż$t��h��њ(!14<��s��"��R�Q%�ߝm2_��p��w�ށ���<�`No&w�����)|�wX�q����$b��߭�1k}i@���hvj�kË����X��yLVS�#��$��W��Т{jġ=��׏��K���@��,v�UC�jj"�/�H!G��!i)7g[���&�HK�Ĵ=<<���]�`	��Xt��G�T6����m1�;�z,���v!��%_���k�Y�Nݥ�T�����3-)l�d��B�VW�kdi�;99A����V�W= "i]t�|��g��
%⪼�� 'C�j����/�f��o�10��w��h
���J���3p+�����+�K�#"�R卺�Ɂ)O�[V��O
���TS�ᆃ���L|3�����2������Z`1#�(@�Qv�+�sg�N�u��ٺ�����UA$#��RU�ɾU��Ew�>��&��C�h&�
Ʒs�����Yd;]��˃�h#BJQQq�Mן��ُgyF�������n@=��w�\��ǩ����O7$�;/@�*R��9���c�M{�$� �&�vp@^�d��ONNf���ԟ����0=@�m/��$BSиM�딦*����n�@ۣ�k�r�t9�%95�ֿ�2�#�����x�~东�l�7iI~�ؑ����s��I�����ј�X���Q����f����˧�_D\l� ���?�'��RXTE4��R˕����Ȳ_FMM�=Z��?�gj4|�o`����$tKIl���H�م?qT SH�<W�	 ��URd@��e�Q80�]�{�R��Z�.��b��S���C��] 5e��������w�r*e988������*��E1�e@2
��
*�s�DE@� A�E$I�X�JQ� X( YA$�R	*I$IF����t�s��9��ޟs�{�j��&3�����1�Z�/�h�S����;ݥ�%iHt�����Ne��G W�!WD71[C�iU55 ���R�֦^��Y�{͌���{BL�;�|���x�n��76�
�u�x�]^r����M�m�/�'���]�-8h��|��(�7�	Pd��5��O��qAB}�O�C2J:�"5x��A��`pS���ն�����
p�}d��hN�l���ȕ�u�_���Uf���v�up��ŎBo��))���C���"P��G���a��P����N�ԕ�����]�/ $���Pf�~�Ǉ�jj�?vm�����{9)�������p�R��/���6
�±�h���|��p l[:�����(Yߨĳ�7��g�����ff�,��i�	�o�wE{M7�J1�����Vq��Jiizn���{_^\z��h���,�0��5�*�NF�����n*q�`�Y!�+����'J·<��yݽ{�|�5�gֹ@�� �h��.Nj��-:�iu	�4��ÇU*�K=P��7�XI�'J"��7:��7��q��@I@�b�#Q��b̞����,���o\ؘnF���a����; yV��ǡ��	�g^\%����?��m�����F�ۛ[���w�!��D�%���O4��C)+((׻��i@� NMj]�K[y�N0{X��Ā��l���6L����l$�h���!�jOq�B���_���a��ڐz����=�	�k	
�Apz<r)�Z�vOy{��������P\T!�̶�����}���7�RJ9tu.���Dy�6A���t�p�N���ӟ��:z����������uTJ�4��2Z�/�N��%]Ȉ�X/yɩ��?F�q�raP,� ��(����]^�}�nb�7k��i>?~�Bsf�ʡ�rʻ
�֬.��͓࡝��,vd���0(���֬a>�t�<	rQ}����b-Nr�Z��9u�9����6�B�t/�!���<��� `�{�#]����]D�L���Ij*�Tu��/��t�y�g�B%����M6�^���* �;��L�����]���ڔb� gjC����u�&�nnn+�K�ښ먯�펽�utt��g��d��6�z�< 8��}	�hW+�2_��Ն��������v��}K��|��`��"��u�LϷd�����S��8
�B�;_U+����P8oC��p�?MKK�g�tV��<���ƫȗ��s�:�Jr<a*����{l�եw��D{�in3_;F��%��mv��j+:-t藽��Oq�o�P���u�ߠT\IP�ם{Iq���~­�3�z��nQ.jβ1h�uR>��{�~���	h����?���x�p	ڬ��mg֧��(�(������4�Tܞp��՗�{��:�{LX�Lo��������EU�><�s|ݷ����/G;I�ػv2�y��U�꺪��0�X7��ʚ��� �~��.��z���
��S
"���N����/*���V��ԟ#�|}g =�v��[h��l�N��3_{����(�TVr�0J��%��� ���|7�>͑�m �bߟ=f	�-:bj�k&�	

B��:٥gN�����������ݭm����`�_܂P7\��AGL���]]t�z�g�9��	,��(��<v�~,��jӗ�"}[[�� 9��赆���~�a�K6C���kٚ�H���A��4Y)�I��j�N��N�B4!ޝ2LIL�<�bl�\�R�P�N�������l��.hWp����Y�Ke�.�ԉg'��W�Q�, G]]B�y %o���Q� 1�.�\�+S�v���P*�C,��1�� Ud��)�n��9�L�L�2�?!.�Ƨ����;k]��O��$m�&3
v�T�i� c�[|}pN�%�����ggg��:Z�[��<�n�"z�H$�^X��er`�K�=�+�9�S�X�����%)�	ӋS{�������zܑ��<�2�� ���#�op�411A�+�G�窕Q�L�ϡA��M���90oA�������؉��X�QgRUJ�[t��܏FQd�.&&��5�;@F�?����������~�3���!UO�J�Em���$�䬔�^�a��;���٢��0�$��yg���~TYϏ����wBѮ9ˇF�o߾y0
�G�����	��p	 K4������߫>����(�/vbA�5]m��p~MCd�ʕ�[v�n���ă�`9�;>A)I��^,p�������9)%�(��o\�ˆ��7(��-\|(6�ڡ���Hɗ��15i��@�b_�/�]�L��1ӓ�0��~~����T��h��"�P�������*�ċ��VS��N>�S�c��w�b�QJ�ph��@ݾ�0p[��&����̇�F����/�όw�?��#C@u�[��{'�e�bR�)�-a�"�O��?��z�}k�CCf�~<��,��FH4�Ywȝ�؁36 ��}ū����]��n�?݉���(q�/���N�}��sx�]�9�������KÝ�.�~��k� �]s� �Q�0��E"����)1qq��欗-ٙ�n}���<���~|��>=�rs~��Q�f��^m�366��ڢ�:Z4=h���ޟJ����ڲ-��	`,亮��h���;MaKs]��mTV�(�]UQ�:/�ܦZz�u�H��8 ������W�v�(!p�ݻw��س���nq�V���@E�{J���4��	7�^>�%(%F����-���o�������xqq1�f⿽����|Z"]���'R<v#$ ���a@��a�@��H�)���'�ԙ�~��;��Hî�~.��FI�
=eA��g���F{�I���������2I�\��⑰�nY�0��S����=K��!����;���_N�8���+f�]�ho�vA /?8]Hq��y�Y�'��6g�@�'�/t�)J��l�~S%�tDT$�l��$����˖��b;F \�[^�07�2����u��s��},&xk�N�?;?E��Ժp�iz� ė�ci���$�<��Z[�iU��]�v��O�갧��C~��"��b�ڊHii�֎��ٳ^��[Z�RAA�oOn�|��N)ccc� ��a���}_��,����֦����k�P���l}r	�D�_�h���S"���fH{*� +*)�(++���馶�:���S!��pG�J42�����ɨ�>����#��"'	@lA07�4z>�B���0���ͮ]?jʋ���?�M����S����h'��+>�_M5Y	O�sjjt��U��.dX��
EO���v*I�&�H-.{���n�0A�Pq�������ʵO6�d�n���.�X�Ag��r�4�N���|�ɴ6x�{�c��f#�Y����I�ZI����ж:��|�;���^D�oș���u��6&��7��GBhE��a��ND����Fl��c��X.��?��:��_x}��0��_vTJ/�B���?
�Wd��ty4'!9yH,/�Q__�;������1��8q��?	�E�rt۠��+�.���Ru!`�Ƒ��ne=�=۶m�\Z��k��]7��8K1Kq]�b�/�E�C?&��#)��)��W��	)��`�����{�4��0Q��![dِz��U��R�����A�)�.F�qU��܉f���6�Ag+DZ�h,:����VԺ8L6�����_�n
	-�G�쵒cx����\gz��/�b�dz�p���0�oW�&���!,�<�I�12�O�B=���I9�/���SYC��m����&`X��J�>ϥ�9��ո,�ڨ�Ol�(�Ӄ���{R��7����8��kmà��68r,���Q���i��\��{0�:��䯓�N�:��䯓�N�:����ѓ�{��6��ݺ4��5��ţ�����t��c���������U�?w����͜�k�^��
����y�ê���_��o�o�p��N�[��V�~�����Ͻ����E���_	�%�����KJJJ�Vɭ�����X����(����N����&��������c�S�Ɩ�TTjW��ڸ�������I�N��&�n11�S>�md�uq���V�'M�V�'"���4uf �֟�YU3�u��~�����=�𵙡y?��>Ӯ���8��a��$մ��.�W�B��<�]\0�7��QO5j��knnn�.��Mz�`�}���ƟW�)k�H���&¼:�/T�:�pqq�V�2��l��ѝQ�UkP\�~]����8��:���TƂet�X�O���ǻV'X��c�=���b�����Ɣ����ʿ��K�/����8b1Iq�2�i!����Aܽ����$''����E�s����p�]eSS�e�����):F������!y�W3��{z�'���Pp�E3�;Mn�֞�MV���jZ�FT��@�0��������K E˭�w�ۅ��K��E�+[w�ۺ��e�F��[�:�L���ެ���?J�_	�%��_	�%��_	�?!�q,��zX�veeҽ���xh�'Iifվ�ȴ�cV:�?��N��8>�ƭ����O���s�*��_l#�o~A�?����K�/����K��;�$�<�R���9B��<?��˺���{�2>*h�c�;q�С#��B�_����]�_'��u���_'����I��vJ��#�9}P�l��s�N�|�^���������C�ˊ:��;���x�./|Q�n���N�U+��>��5M�z��bk|q���d�5�|�r�!�耧�����3��e(<e����Q�M�چ�s�Tda����!�%�{�8�K�֜yk��a!KA6����y���{��pݓ�X�G��T�y�g��"��):���z�z,~�GXNz�^=>n��vk<~	�+������b�y�ؙ8�Pۜ�3d-?}�:\�c�J�=p_��$���&""�L�JL^8����JZ�����ԑT�_3��Sxn���n+��D�����%8��R�ނ���r�@�
8�"��󔽐�n�\B���k��QG�c��_-����t�*"2R>_8��y�8����l�D��3��r����)��Z@!��U�i����ИCX/��`]�\XT� �=nx�U�9�#Ұ���a�Ǯ�Os?Wk�2Mk����7�S�����Ĥ��`��8f���s5
�)������8�,��o�n�#�ʡ��)��A{��o��֒7����Hx�3 E��k�j�CDr���ԏx<]�����H:E���oOi|�P����j�t47:���* ZD�\��QL��'�s�G����}_0*T?��H�El�!�`���[G�絉��tqr:��Ĉ��rK7e١���Oc-X��߮��!;E�l� \�_@�*�~&��ؼ������y����������J1

W�j�&���1qV�&�Fq9s��YZ����! ���U���-�3����_NV��l� .��dl�	��C�����tOn��A�B�Cb���2����#�����(����1��j�����+zm�4�&��ﭳ����!�]+B�"��_JRO �+�ayO(x�I�qe�9��a� sH:8�ow���h�y���j���\Ľ����1q����p	8ڢtA�9�$g���Q��v����D��L	��$A�h9/b�Qe<R�_k��	���v��}mNN+�H>��#I�f�I��b�wY�an���'w�"]�����r����?���sZ��:ϓ#�c�CV`ĜP�EƲ�^sZ�c?��i/l1g@�2�@8�g�	1���r2�b�!/u�r���p�u;���l%XQG��V�`�O���
�Ӓp�_���H����(�M���<�7Hr!���T����ɍw��z�p�_�v��,��>���p�����]��Z��_�E��q�UQ���Q�d.�G.�R06[�& +ޮw���,h ļ�)f�M\�u�q�Ć7� 5����2�"�쟝���7������!��f���,���S|x18C.���^TP%�S��8���,�F���w�<r�>��n9��J�Һ�bǑ��U|�!RL/ɉ����?Kv�(��9gD�j#.����,��i69-������X:�����x�w�������3��d���Zةù��,��(�K�vb�
ƅ��Ew�B�w:)ƪ�S!��,�q~z/���[[li�
6��0�zF�e|�Yh��B�6X��	j_8�L/WUp��v��е
ӂ���R�/�a�C�� <����gh�'.Ml�_����cd�m׸�J���l.��Nx��{6��. !�q�0|^�7Y����_'�\����Ts N|j�;�g�*%b�F�r�Z�KG�
���:�����.�
fB�����뢀�O:)��B?��bH�:�zV�̂�ܿ�q2{aԃ�U����+t�[���L�UV۟���8ƿ�J�i(F������ �%��WYp��m����a\sz�Z���^h&_\0�OF�t�@{
��	V�lbG��N��r����&����>�[�8Ym����b�?�ܽ4^�oGvy� �P��, �w�A��B^~���귰������Vy��<[��A�8J�*QӜȃ�������&g�"Ռɇ�OY៑���wf��'��ħ��$��〒����C쾝�r��j�������	�V~Аm
뺩������L�h�`c~t��t�w�3�M��>��V��8��cϥ�J�&���"������s �L7`��r���9��BAz�����~���y_`�>���M�`�1�ǉ��=�g%ͼ�P/�%(y����6��6ui�+K? 8O��7.�h���D�ry�Q�M-�zvo�M�L�y?� �cIc�b7��Ә��;@o/,X��y���Xd�qb���6ֶÔ�O �<��<}��%�7�fi�-��`��ͅ)O7XؽUؠ��\A������`�����a���s�R=�%>⛯�'���|g��H�ЫM/4�K\���\��W�}�I��>9���֦�ʣ���6���w� ��љ����k,����*��p�aFP�M�g�x��6�]DPO|=� 4f�:ݦA��u3����#,8���&��Rk�!R�V����=b���rWS�sL���J����A$X��y)&��~��������O��`K��j&&�����;�S���F`����DԼ�6�q���r}p��+�{dd rY�0�j�J���αm�c���Im��l
���!�:�g��%�7N�����L|f�1��N��z�+`;���������TCқ�0�Zd跡z�k�q
y`���i�X}>I7䔥�o�'�kz�Đ;�pݥ��(h�5=,������G7��Ɔ�c��Y�ۗ|]Km�7�k임�@��#�+�u������áa�K����@�G���H��Øh�=M�!���U�]�e�O|m�N��#��q���:���]a�5�Bhk@�e��@T+{�eh@�)��;�h{��'HM�ml���h9*6�z����S&����!�#1	�v���
��	�ȸ@��a+	�w����i�҈�ݗ�m��'fx��>�A�YY������v⵨�*�w��0�D+�Zr	���6٢Q�C��M6!R6��d~d.N;Z���e��\�s�YμfW�qW
�\>�����.���� �?�u����,�CO�+��ǧ�!4nm��pn�5��n&��/�;P�΁l��p��d�h�6�"�J���W@�R}*oB�,ݔK(3�}`���{�bsV��c���(�}��'�[�Ÿ�}��OQόb��Ȳ�b��e���a�Ox����C�hހ=�	�&��.F�@C �a�=��xp����'ۇ�������δ�|��7�6���0Қ��d�>����)��Oq!��D��,��k�B���rH�z�6��F7QE���d�À�BP����o��.��pֱN/�G��<�H� sK,��F7C^P�	���A!-'�;�Z"��� ��l��Bl��]��˴R������e���K#r�5�̸�������3����i�Z%�.�ݼ�߄���(z�ly�~֟}OT9��.�ԯ��G�f�r�&�hhvS5q~��s��n�X����(��K;��B3"��VD-2���"6݊ޮ���Sn���� 0,a!���������\�M@��+]_>����0�?��u(I� '�%�e�6w6�;V&4�	��";�__��u�)���_i��P�j���|nf����n�g���^�h��.���t$`���7���A-XmgIo��|�`�Nm���Ǟ':j��]���_s���*+��Jn�Q_�t�K}V�{���<�)�+8<��f��@^��@�|6�ЬCF�r�]�
��j>��р��֢艭!1Ff]���Z�0�z�?�tJ.��;@.짉����O�]{kA��J:�g=�u�\���k@G6⊯_/i%%�+<���b�#�Sh�	��ݏ�����lA�3D����~�j���RP�VH�d�<�����I�%
L����w��}�n_n?ǂ�z���+��ep����Y�S��R-j�_ތ�� ����3g��W���SX�˚�C�B�*�4D�pV�8C��{�޽{�/M(r��Al�G�[�\��.>#]+$:u3�'.5h_�"5���Ėk��vC%:>�r��v�f���'�>C�B�nW1ҙ��E<�����mL��pt����%0��)Ȯ��_M�q,Ԕ�a߲/�{i`�V]~�~����ǘR�A�p�3eB�8hܤ V��1�
C�1��ZI��WZX�>�'!i�*�<�C$����cx��#�YO _�;Ԫ/��� �Mk��{���@�n9r�0	�?��Ğ:��n�S�2�5���KƅqN���N��f#r�gwȸ��l6������!.�g��2������ܰb�*8����E���2{˛mV����{��Q��6���O�f�;�3̗��D�|�l�������N�ޕс"�	մ��$��Su�������(�W�7�o|�}(�3X��Dmt�Nb�q'-J�+΋�͞�U�����2*?�9�,q!�"�i��J)=y�-�Wi�?�ITWX�6r/a��.:���k��
Gq��k�r�uM��?�B������y0�����@�-IP��W*�}*�ȹ��!o�/��{�¯�X�����M� �S��
u����"���R,�R��0�]��;6���2���5Z��jy�g��e�ol���n��ij�� 1\�N��CF�o��>#�֣���,d<Q��	�IN�Ѷ ��~[x�6��yiݯ���rd��ŵ`x�]����*�����؆&�"��:����,��9� ~�G��������S�T�D_R"��k�$�両�Q\~��e<�Ϥ@|�A>�	)�,��5��g2�~*�I���D�瞫���j�V���������>9ՍR��߰��%��ʎ���02�C�����Mُ��ߡ��ˢ��΁��wq��I-�n�d�Wa�69��	D����-K�����E��q��Ap�<����f�S��W?C��~���~*�< ��	�6����� r���*8#����=N�t�*g��a�N���A���e=l�}�y��CW �m��yn�]���UM�OQ*&9�ǿ�q��Cv7�}W��,c�I"
����X�h��e��ot�ّ=�u[_5�`�B�����V:T��!��D��"w
��� �tr?����--�B�����1��{����d*�=�dԸ���HZrG�:�m�BJTI�nҾe��KȺ/:W���'�;Lv� L:��_�����n�����l�^&xe&=g�&-N� ���G	Lx6���T������ƵB}��-[���"�����+��\J��"�l jd�uS�_�X�cu��d���A��d�c����fA�Da2���'�r�5���8�\f��{yXY���= Z�~Xy[�5Se�Ĥ��o�P�.7���~�lHe�b�i���c|�ktg�>zzŸ����V҆k�O�'���^-s�ƽX9�#�l�*�[����Υ��

fl��
�Ė�?�/�����=�#6�wkY5'4�Ҷ��%��5���:�鞁r�& �q499?�:M:�q��"jJb"��1��EF�J�r���|��ŀ��'1�<-�w��؜2q�iO�4K������c���w[�ǘ�C�V@:���9_"��Ecc״����bK��������[���z_]�͗�l7���<�{�� �w�ǌ't`�i�r1�ѳa�l'׊qI�s�MI-d��12�,�u�=Ed��ђi�͸pq��b�����<F�����g%ŵ��O��?�A�u���~2I���V�h���G�c�k����N&��:�X6���s��@��A�bF�����cn����!�H���'�D�g��`}ExF�����nKI�"�FFݴ�3D���3�:}0�b�z�)Q�j�֍���ñkC���^i�
�ǰ�A��2Ϝ-��]�Q{�r�Sd��iG���n��OC��^7D6�Z��5ӄ�}͊w����ry�K�T������;�xVJ}�ll��8�O\�L�w���A{�+�H{fjP�;�+�$?w���>j%&%�*Ӓ���%�u������f�5a�շm��@�H�xll̻`9I�t����U����k��M�'�u�o��!�do��[)�W̽ON�\�15=��B�U�f�3�#u�L�
�z>nQO�B�=�>��M`h�-�5����ѿ\R�}1*����W��~zE��ӥ����E��-��y��m�v���:������;Z3���?>nD��]#��
ȩ���&����,xz$q�K�gO�E�h/��>R��l��:9��4u�191���{��������i|�9;����M�p�Zq��n`�J��+�q���*�e�l�ciJKKc���,#X=�Ӳ�!p�����'��Ƚ[�S�J���-�M�/�#X0�z��3M���L�5���$�Ϛ=ֆ�|z<o4��D��F>�LIV}�NTd��ǉ�B��L��6�H���]��M���㉿r0�;�]�"77��="��T:76�FyMLL����z���=���0n�B,EKG�O1֦cx�삠�����qvn.��2�%������g5�J�E�ʑ��i?&�=�o�6p�
�J`�������B6�.���c�����BB�Y�sXM��w�Qr�&���	��/M|C��MУJ�UeG��MN��]~'<���b���."0y��z���\�i_ff>BF_d��켶��fnn�>Q?�s�p{>���� G4��+Z�CR`L�v�4(���.�c��kkk��O�'����!M��kzu�91���bbb�q�#��*������ V䬦����N�!.��7D\@���2��I�N.�8�9U�	q�����t��e��\� �llƗ!���[���ϟUUDFՒ����7�r�1���{�����?T8�l�ZPw����Y8/:��n����ߡ�����&FF�ꞕ������ �= ,�&���%�A�˱�x㨘�8�|�E�$S�P�M}c��=����\�!��v&ϊ�����+'�^�\�¥�O��и1�+d�Ut�<���׸�Є�_м�2�^�(ڟ���-@�K~�5 �FH<����3����-��0���CLE��9}�\T��S�h�B����|BBB�bbD*&��(7��f������]7޴���Lk ��w���@���Ї�� K%��,����I4���Fsv�
;���N{ǯoo�u寨IܐX�~�}[fN�6WAP[s�D��Pi8z#�9'n_�o�~{��s���N��!�����RKG���@כ��e����>��K#6�4�ie�$����`_�'2y��/���^�y;{���͛7�a�;W�|�G���P��>/*n[��
��m/ �s�a+j�.�"�N��ǡ���Ӫ�[3S��cj�B����1F\�tsEVrH�]���1>ԍ�^Ou]]@�����[��åpOP4))�o����pT��i���~����`SSӨ6+��y���ݵ��|{s�r��( k'"	<�Dm�O@��БU�Mΐ���u} �ein~�'�T¦�J]�4��t�~��h�� �V��3�ǻx0X,�G����"��H�.�q�CF�y,��Àx[�?�c��>r233��Y������J$��0�X�]�(�Y�S2�0 t#0���V�%���E�4n�E�2����T���G�#5�Ͼ��?��'��TdT]���`���1�QD������
�Z�X��]M�2H���J�T�킮z~LD
��M����5��-e���^;d�mr�ɿ�.��JzU�B���ԼCJ���˿��p���]-P%�@+��]�9G���-C��%?)�(�"�nH�LY�g/~��wO��Y0�Ov{��{�/Ϲp��WC�ys:���:�mU��`���#G����7:PW�����?r����Ȋ�Ө��M�Ccݥ�[�5��| ��))(��u�Ƙ����-�eX��f�{��$ҩ'�2��1��J�srj�����zj�%�U��r��=��޺���YM��D_!�K��;�N�<<��Zn]}}��50���HaRS[Pԩ�q_��h�egow�ؒe�ae5"I��I������)��f�Aitv2L)g��ډ����}�o��"��u��1���$!�y�$�G��H���b�5S�]Y�M�íM�۷Gx{�nB[
�n�C�j���P�-��~�Cļ� 	���Mh#���[������ܹ��z	��Һ��M>��eVf2	[<@�Wij<522��5��R�y��{�@�цJ����z�F�E�8��@���?�,=�0��7�d�/MmN��cjA/;����2�hqG��S���J��>z��/����[ ze�� y(6�5��C8ڇ|0��s+T���S�k��������"c��ivP�@�g�.���N�s�n��;Mr+n�w���Nv`��z�'�٭w�r|�?����E�1_���Obr�7[1����#�۷o���& B�!
bu'�Y�<�DCMm�]� �6�st,��4��7���Ä�L�V��x\hZ@���˗S[�=.Wmpշ7N�tS���8����ٝT����6m�PV�M����ַ>�t�hɞ��j@�P�U?z��ᄀ���pj 4lq�{i$��CN8#d��X���Kʴ����Y;bKS���Cj�m��)����H�K&��>��[@+P�KO���H>Kk�@�s����!���o]��X����i�jԱZ�xxأ�.�B�CNK���DM���}�o��N�&�����13^��P4���d��}呚k��Aew�2���T�]�X���Dj	��+s�i�Fv�ͷ0�(����ଔz���������(�7+U=wK��(��?["��J��W�/Í��:B����w")�AF;�5�����J�,^��>�Vݠ�&��:��&'�ڮ��ȓh�T�K7e��k����Ԇ�<�ڣb]Yg����e��n#Mŗ��ًuwN>����^5�#+��.�8�x/GK5�uڢ�iӜ8'�v���m��2��ʴ�Mk)H�4���S9�&����w0 V@��,o�T������,|����$���:6��P3557����K=���yAs�[��qԽ(����kji�����zpȱ���J��.��~1h'��E���`wW&鸰z�ƓVVFb2ci����"����������kz&��s�[ȵ7�~��e�w����^ʳ�>/��� �� �B���&�TTa1N2�	���
66�������ή*i��Lbaaq���N�mjBX��~����Qp�YJ�}G��~�������xR����k���ׯ�y���"�yY�H';�L���2��L[988��z���/t�r�L#_�~���޲A���7�)�, �(�a��H��Xse췽�x �W�`�+��)�{{E���e�F}ikiYhyj�vȲ���7�t���j�&IpΔ]N �w�b�b\FZ�2)�_H�A��L��&�Z1��W	�-7>^P6x�FIz�G۫�/��VK|ЬGq$C��ec�z��v���
ɍ��Z rm�rRh�v�nm�M�h�˯�P�.�}(� PX���aڳNz����t�ŕ��2�
���?��2�Ҙ��^��2����j�;_t]c�Vbr�"�s��{��8:N�*��]E�[r�n!�9����"55n��ń��Yy�@陛��̚��g���,�����9�O�Bu.�C�Ά��I�$�I���z��6������n��D`HKD�.�� ����.�֩
���Ns�� ��V)�}{d
����tK�'[�k�x�+�4S[������*PN��w"�p�s�K1o�ۿ@����=�����Z�m6�����Y֝�7���E��L��ױuD���*h��>��અE� ��
4
����$�������h�g��Z�d$��u�'T���
l�Ҧ �ՑWs^n��cU�67��Ng�d!�L�5Ԑ(����<{="T̀D	wv�Ia�z�h⣃�1�p�*z��1G)�?al���8�F%�Ѵ��8���f�00�=�}�-""K=��+���k�xE>�G|���6�~��N�lh3�X�G�=mL�+B�l~��}��evv(�n�j�t����T,,,,���%�n���t�	1���7��X3g,�x94�Li�L� ہ���p��`6��L\F^�n�r�(	$�,p�jkh@M��ǘV6 ��\.L+;����4>��&�)�&�+Z���UUc�JO����6���l�� ��Dv�j�~��a`J׹�����?����~/�2��'j�M����Z��$5s��O��lc�4�!P�t�J���S���L@���h��a.�lZ��&��L�Z�88iXT�ӷ�E�S�p3��27�]����H�i(Jh���tV֝'����bL��:\:�L���w,�S���TTTȬ�"X)Q,{��0�
+�E�Z<���I��2�`J���o�t-�����P2?��i�U���"�0n�-)�![����� \��Ą]���M�6b�I�)4�n!U"��143;����XB��J�ejj��]`WK6�k_sች��WR��na2��#�#���0�5S��\�)��.S���a@ R9c��a�Q��`vww7L���\V��\���Yꠦ6���p�i?�ǎ7ͯ.���l�fں���J	�9�)|[Hi�����,�"��p ���e�(��?}���������2�00��I^��ؔ�W����WU��9!~օ�%Ւ���X"b �sT�����n�qw� �C
�k�ܜ�Dg�q0�d
���fT�Օi��u��)�*4���*p����� 3P\U��S$���6�J��a����S.�U���f��R� �.�����<g���^0��i���]��S�Z"��`)�B��d۠���D�*wF�#k����	� ih�2�7��MP�(=��F�a9�����TkI�7a^����f�Q��T �$��=��ʿ���m�����D���o ��q̏IèP��a�PM������=>�R��x���E���J�ؒX��\�2�M@�]pWq��2����Lʋ�O � HQ,��`i&=7�y˖-��f)�5.]r�K#�J�0v��r������W�hn�LII�#���55b&���->�����U#�0k~��+�Q$�uV���ٚX�+:��N��>gep#@y%$k�ǏgT�f�/@���9�@{́p�A�r��#j��j������x%%b[22������� ��%uu�Z�<�/d��c��DfZ�պ��-˿I/�j_:���JE��l���f*��t�����V��CϹ���=I�� �9ҌT���
h%���q�Tzf����3��5�o��7>��K�1�)82%(yN|���̀�ի��4J��]rJ�VCY�ꔔ�Ҭ�Ps���V�� �0zw>��=7�"��<e5�3u<Gr�a,������^~bDtG ;�?�829��R"�:��8fP�=Sc5������v@�]���K7��;����6�r��t����-\��0V�3@q�Z8<B��hqhhh��wS��m�N6<�[��Yz_�梁�_í�rҳU���%��ˬq�0�M~���Ĥ�S�=i��T0�N�ѻ�;������<�he� �����>1왮�eٜ��}�%*��o��%�aEg���x��T�P1��K����.dg��ڑ����.'��k�v�bM�o�Om1|�1��s���������R�3<����c�n�6d��I����Fl��JQPT,���|�3��s>���0�g�&o�4�h��秙p����d���X�����V0_Z�*����،��H�hA�D���΂���w��۾Yv9�˷�)2�8|�M8���.$�`g��Y�Lby����Υ&�����f�Xd��͎��ߟ���hLlF{�%T��a��1�_j��1u�c�ToqL���m�K��K6GY%Y?/��B�:-�;�y�^W��x��WeZeڢ�vxG�9�"�e0",��nT��5y��(��2LEؗ���QC��w%����1��O[,���Fs�M�S��j	���������F��[�����a��|����͛2-ڊ����؃^�$�.V��j��c��`A^̲C�㽕����������#��)������"@p���p�g��C{�2\O;}$�sN��d�d)#0���Z�?���RX��O'k=�ˇ�@RL���UKK�o]*�*�&��֥\*g�b��\�G؜����CK�T�C��:BRR,�}�'��u�j��'6��a��r�z��q�>ʂ����z��m���>���R�܋�|?�%QM�j�g�Z^�(+��㐿De�dZӗ/�����򳨑c2<����G#=.-�,��.�����@�e���VҲ43�?Y	C��"����mN��ab`�	��]��L���|I����Pؒ�����5]i&�Iꁵ9~��k���{|��^]C�Ǝ��J���>+�������)zyI�� -S�tN��L%n�����֝G�J��_љ�"��-����M�J�V�]֞��@�3�
f��I=9�?;��T��]d�1��(x�ºާ����U�N����R	Koa��3�L���Ց�����h�\����[i��ӳ��N���[̓���h�oh>���իW����M)��3���.d����R�"
�J��VV�ᄱ���|�������S��O>�:U�P�ѡ������#T_�����(��$��ob�� �Oc������p0(v�*�C>z ��S�-߄t-6�i�`f"Mp��&�,LU{E0B�#"��L���i�Z\S�g�3tr^QQ��"�!z]}pP����H��{��>�)0=kK씗�?�onn��͉�>�R߯�"��$,rW��)�.��R12�Yx[��o�fW�,�3�\R;L���4~�qgtt�ѣG��-�'|�2�������~___^A���ü��dӵА���E
���%��eZ��ӂ�ެ{������u���Ij;�C��s$F���5�7�,��$
n*bA�8W5��&'���rr�O�k�	j�DD�UOx��
&�UR@~Dx�T��JOW�����L�LYy�,���.��oE�����B�y����1	�a�J��/"�W�� c�{=���렄t�"ڎ�oǤ�i)~���0&�@�}������Rd�g3�Hi�Y����%��=?;{W��� UU����H����4������O�Y��e��{���U
�����VT"�&���&��h�����ՃW�ĸ�,�8���i@b+hWVY�?���:��Cg���������߿�cgy������5̣;gB�͹}�O�-4�i��7545�ה �ÏS5?;�Q����^7�5,���SO(*.>	Ѽm�L
�~c���f��B����k����>�lM'^P "ǥ�ӥk����D�s�	������8B@awτT�$;O"j�!nU�����*~E�4N�9� #6IUZY�j*jXu���Q4�f�b�ڈ�6�����Ϟ M#!!�Mz�4n�)b.#��LP2-�*�����5NI���rH8�2�wg��{ݐ���O�k"��s��J�N$�Tu��O���,p�9��GO�\�ؘ�职o�����s�;�kk^�sDn�dg7�v�O3O+�^\\��4rS+~�X��*.6���R.OWI��)�I���悮�/?ջU�?�,���֦TS�=C<o��뙹��W�?~�8U�*�N~#'�̮�IC]]�ʕ����g��]��J��5����Kt�F4O��@<�r����3�����1fM���>ȧV�,��SV;�ip;3�rB�>��%������Ԧ =(8X{�f��'��p�L�}��u���P:�f�QU���i3��S�)S	�7b�^F$���9iA�b�y�0�(����-�v��������m�?��������0�H���
��lS�MO7�ѣ4S�]� ��r��K��&A�x�t�޿iӦ #M`ZI�b�}����8<]��C��룁*�?-�!�Ѵ;��Ғ���/�¯߰ӥT��
�$ǝH��6f|R�}��eF��x@9$����L��c�v~�0 	�kKS9'���ܓ����{�!�8��һVݡPVQqP�6��! �U� ү����=�x�J���:6�8���
ŷw���aR�����ԚA���Ƕ$Eq��]��yKK���EEE�������������xq��	����MԲBBNk��v��D*R̈��W��ޙ����<�P^9�>���uu�ж�VR��+��	Dp�l r�[��)㌐h�_{�����\=�C���_����d%�C��!�:+G<��>�ߞj%�}{�s(;;;���ӓ����z�����ԡ&io+�'Y�������H������玄�C1#�� ��sr�ʍ�Q�#EћY8��ޗ��9T�ځk)�s�&D����8RU���U^VVXX(�9NP�O�1�755A�t��^���gv��wK�LrQ�Ӳ�����Х�6!{&�znn!l�����~H-?&��N�<����1I<�V~Ю=~��5J��s^k��F����j��vNR�����{�,'��e�ڇ���m_ߕ��@ٔ��ą_[%��|�u���ʍ ?���e��)�k��`e͕t��>] 1)��e``XW_�50x���$���<z�����±�k�C�}���f�oKBY�kX  .�ٶY<;�5�H��-!�^]=�`����x>��t�����/n&6��RV]]��ك?2F�o3�G�6�>#�VNNg�6^��&��#5p��&�~v� �>���?i�ʽw.��	�慄����:I��������@*�6�f흙�T�üm$��V��BR"{����6�&�B������4�b�萎�]$뱄sp8�뺟c�����y��<�s_���]��}������/Z�}�`$�8Ӌ�b�n8HZ���x��jV�ZB�B�$f����&Nv¡/2V��I&jn�p`P��l�V��c�(i��}�:tI�u�xAa�j�%ըY@�'V|~���a~X�d�ɿ�)��5���r��Iv�>��e˖(�m����c��}'0��n�A��yN��������ψ-��o�o�u�=��ْm�����8��>���5id�ΤC�{����K�'R�����h��X�V�3ˆƶ�S��~,a;*����{(�u�U���4�����Py8ef���nVz������==����?�8 _0���9i5��S���'&&>�3���nrWi��_���K�6��M�v9u[�nK���8�:;�0�g,�R��R��յ}��b�rM���;�-�לhѺ���z�ef���J6��Xl���fy�'�666G����#T��� ��&�������g���|6{�h�~M��;����R�w��B�4Z�@  >w�,��#	Uź�I�vj�5�y�z5<<��q����:S3�0��f���^P+�=�� �t'������AU���J�1�&��r,��*i��vv���iT��@�2��g�����vc&��w��3�T6���Ny2T>66Fw�R+�������EQ�-��ߎ�`WФ��!�K]]����Gj'�+{�˃؊����X۷oI��"��&VV��c�,��،����{f��Lm�]����R��S%�m�:456^����X�h]N��o5-*)n�25ՆB�D��v�\ڑ\o�O�D��ge�}���-��0'ҿ��N�B��M2�����;��} ���Wow ʄ.�e�am��k�8.Jm��l����u3�OQ8C�T�3=xv_���������ʌ<�@�/c��nx���(�]|r�����f�F��Ò�[6�0�̨��X�[h(z
>�V<+��p���3�l+%�y����g���ؑ��ST#v
���~۝1�ma-�A �9,({55�5i��.���5��?���a��
;��8ɚm߄?�(~����f��m]+����ג�&Fo��0ε/�{�uH��YyV��?��Ηa���7���Y��2��mtrr"
ǹ��iA�ܻ=~�s�Y+_��Q��㣘����['�p�@�]�wFY�&�9G� Q��ۉlH��n�dԍ(8��j�ؾ@Ȭ ��9U-]�^���h&)������S��ףYYX�OMM���8~7��l�~���Y��U�tOu�����L�x��!�k�[�M�B=9��l|�r�����_�R��Ԥm��7==�ʣ��Ԃ����;v�Αݾ}s���..۩���{��&�t��L��.ᄐ-�7d���Ǐ���\�&���[�BCCw�ݻw\|F��+���+��'F���>}��f�� dK���ZZ�����M�&���X��6�l�KJV��O�(�o���!�ܟ��S����-òb��{7�I������u>������|W�-��f��Op[y�����.,L��3�S����u�ЗPmQ�"<q��x�ν��[k�C{(R:v��t��ȹ�ؖJFE�������<pkE��������'����:��.BqyQo�'�X��x s�j>��u���ѝ�<����z���[C9����iCi����ᾀ�y��~~����ଐ*d������57�bM}��[�̋����'��NsF1���(*� )!)�5�U�P�Oo�el���@䫔�%Q�Gi�쁴E��B�>��ӊ����,���\��v������*))����Ԡg��!/���w�ާ[�^�r��ο?L��)P;!c�u��) %M�7Bо��]�_�|h>��S�y��<t��ϟ#-����[y��l���qډ�W��9V��bNYg��2̱0:�c��u��Q�s"���Xh
Lr�[��JF{�7E(�ǅ�.C��8;�6�A\] S;�� �v�]ٹV��7�v�3�^2V�h�� \�NZ u"6n;[[���:$kYq�(K
� W��*u���9� y�v�k�L��-j���y`���L�Ie���l�,VgM��F�=R�l�W�����i�Y���I���D��꾜�	�R��Tt��)3�� &8�f�'���h%( ?<�"���w$~hl<�v��9�U��?]<g{!��}H7���x�n7y������p��Ǐg@�T�{fA��.�^���)(q@��m�v)(�T��dL�u��1���Pzt���f�.*����=�K���] �&+����]k����޳g9���C��|{敶��	d�V�z�x�\e�=i��i�	�8�@7���Жܻ�&A|��Z?}
u�8�F����'��p>yAW�u7>>���$�[������~:8�����F��?����:X|@.��V�� ���>��j=,䊎} ��ay2릎�+��&�����Al�@�C�^i>~�x W�wU�r11������ؕ@~������P�ՇaD��0�p˅��ë��mV�UVB��o�lĉ�C�Tfϟ��8�mq������d�ȏy� ?<R�Y���F½{!�FG��������O5��SQq�*@p._0��88<�]nL��g�^��m<g蔯ع�}<��C�%�}�z�H�cU�O����v��HM�9O���q"�Dݱy̶���5��k��$({N��P�r�����\����ળ�����)+(W�#"#����4T"y͍N
M���(��W�]iS��k�o��������SM�1\�7�*���7O��O��a��Z��%�/���w�����.x�e��u�{��'졲 ����!��MUH2�J�ee{�{"B����wO�}BDB����䷝�=�q2��K@u�� -u��$)��3@< �s��?���)(��N*lĖ0��UhM�oR��'��IY����<���-C��޾�3���]"�����jh0"1��S�$�������+��u�[�����A��H�%I� ��/���Ќ�d��e)���/��+�Ml����#��(���B̢��5\�Z;s1nu �����������_kcc#4��(�2J(��
lQB��sM��B������Wp��I�]�A3�����is��'�k��C��4�|R�.��)���/_>���d��)�</��|A^�2�����*�+Q�vΥ-�\w~�'�[=p�g�sg�p�1ߞ�XұDMN�X1������ˤ|��P�����w�o�?���͒�[�
���j��]�D������B�=��7��[殺���P���?��o�K�|'!A&M�0�����>�9 ���s�)5�칧����W
�4h��A�zgGGi###���Y^�V���'Z~�A�R�w�=�ԥбu�� '�)ħ��Un���a~�֭d_��|S��^�9���C���Xjoo�fL}�_-!���.��O�*��]b��f`` �}0���+CjU���ҿ�f��nhI�{�r���K=��8YvN.���u��b����P����k�Q�TpU?��[�{���e�r����\�<�;��qTpg�	5xx��/�d	�����w �&&&px���y�C��$1`l�&\�ȉϮ�����nSH?RkKK��opŻ�]x�jk-�v����'�-�U��"�Jq����ɵ��~��]�eoȼ�-<9�c����P$pK�����PڡE��4gh�~c[ܵb��h��K�n>��������Ez�ڵ��g����[Ma)WU�4� �K]�Xߌ���C:Z�Aq���s	�o0�@���06���?}ؤT3L��o���+ZZne��v�
���FO7��Y��~��N%ԃ���y�j����q.�{�66t�>�^���mm;H��P�i���w� �]\W2��c�D�?���Ķ��E��C�ԃ�_�p-��ݽ��ҡʣ�Rf ʾB`xx��3e��frҷ"���gggg���y�����x&�խ������A���7}��Y���T�Ì95P�F��UQ�1ϗ��G��X�jUگ���������6����8��#��AT�?]S.+(+[\DJ���s�<�f��9x�ch2��O�/�gA��_f��qؤ�o]Od�AQ8�.̀"�*�i�I���*��
���LIU�SΝ`[�*@�Wc����ar&K�@P�1�>|8�����6��3�Fr
�ъ��}I���N�;�������㎊�5�s��Z~@e۳���K>�ؕ �Ѯ*�1?(O�)�b�B���r�Q�[{yɃa�����\-j-{}�F89wi�24���\.��;a{��`:�(�G�5Y���u��d�DF3ù�Om���ۄ�5�ɉ���:���@>��wt�'W�}�
�]`�˗/wd����]h[;�{aeݔ��\�g ]	�7����OL�(�/1�b�����4n��0UW�~b�����m�i��jrR	F�r��b���H|��a��ڙ`_ʇ��@��� D�YKHJ�*��5��슄Qw��[��d)�n���_/U��&�Ru%�K.�@���p&�5p���*�w9�@xd(�h�4�)��� $�#�}�W�.Ⱥ������mi��-IձM�m��Ȼ�$]]w e��X�PA̐"E�%#����v:'dfr�.��Ɩ� ��J�ob�� �Ҹ�q����(���LN�mk����_@���N�x�	�v�O��������>�J\Y򡇂9-���{�؀�Y>����#�����JY���t�8��Ą��}�p��m`bZOI�0Q��������=$���Y����۴�j{�^�.W�*\��AU�����4��ax����1|r�Ņ;�������MV�ώ� ������<;��d��� �E'����ӧ��=9�����.y[笠��
���Nô�{W�o��t2�	6����ND�S:ݒ� ��:���t�һ~����瞞�&3ї������^d@K(���F0� �<�m�j(���<�L�[���n�5#�1"�mK��u��^�����;r̝�֎Bp_@����秱 ����%""�K��3_�-�ժ� �}L�Н��[�:���3��UubG���~ZXx�t����
Z��nL�Jd#��!|q�To�z�8<鉌�f���R���>�(kTn\��m�1~n�;����e���wC�K
��
���\	�`v2\;mt���ӚA�V�O���������DuL����.U�{O��!��%$b���"���ܳ�ϟ?qL���p�V>?�@�_m(�̱ml#c�O�6�Ӏ����!�i(��;����Y,Ǚ�"!W1O9������3�ROs *��66���x�>d�,YEE�,|R���X���,q?DzI%����'>�Uu�$��s�������쟮j��d���P�!�Gvיִ�	,h� �@%AmR��6w`K%q*g�����k����4�3d����EOk� 2d� ��Y~Z��,�Ť.���bZ#!	��ӈy�l�J����4V�'�1��O��z�}��o$�J��#�����h1�,c+��)X�3����R�&a :Ys�/�pe�Ț�?��0��y{��-�����砦�Z�$A���4�c�ɡ3�xC#�]0�!_������ �4�2�i�e��N���U���9���j!� ��F!����!��>����Q2��|3L]���'@jڒ�� Oo�V>:35��_b��EAi�D���)�P���x+�W�Z�z<�v+=�چ�=�nBC����3�J"ԧ���3_�+;�H��wvn�w�m4�L�
f��� ��?���ѡ����ں=[���)l����^�v�H��4��,����95hB�9j{��" �TXI+[@�W��~�6�@��`�i�喰��ɦ"�	�wA�l�$R���ԟM�IU�*e��vZERJ�}g�z���w�b����9�o��ï�#���$p �d �
{��!M,��8Z�.p��=�����8(Z�E�~��{D戄L<kS���{�c��r���pi�]?�ɬ*nV����~$�}! S���TO��fPh˼ǝ�	��f�]O���i.}Z��0aU�Bs����k{��hU����;! L�<ht~UWg@]HEx!��8�b��FB�qR���i"�ʄ^]λ���CXBңlM��*&�!	s}	���Ɍ5b�_���	��xԊA�B�Ī���h'���*���;�,,�O��Y��f'�r�3N�g�^��O��/����ȭt� ��z��V��m��BWo������7��s�]�"�Un��_4���ׯk������̔���$����߆#���hM�Ђl�S�{��a)�Pѻ�~W����7{3k�hO�4��M~��A7��jTand�E��" �	:�l������p�G�h�㸋|�ր�߭���뙙��r���pÛ�ܓ����u�m���B0�dښ��t�0�\�����d��q��ʵ���x�S	�%}�\����e8��Fk�=UC>�,���U_�O#o��������b�ƍH]M䘷��	�fL���n:r��
q|�8_��P���*��Ʉ�$>�Y���Vr�[;r����(ܰm(-���¯<L��ʎ���E�]#Nd�y���6&��e��ŀ�?AM�f�/_��Q�)�]]���$N��A|�E""�޳���OG��ʷ�OzJ��fn�rhȵ9l0�X�f7t�1{{ϱi�}�]Ǩ+eePN9^�wj �d`q�b=y2�q5���3��a2Q,��ب�q,\���c!�o)�s���օm3ιw��v����,�����v8I�!���#��]���/��Z�<(�p�������)Q"2QxzH��8a$P�5W�E�&(����Js��k�&�ʹ��^��	��޽K�K�@:Q�@�eEǜqsۉ�=Zۧ�O�8�>�f��B�
!W�;��~���������t���L�K!j��kntm-;�xţ��K�^������!��ρ���eU��lz��B�nI߹�#F�.�#���ߗZF���E>�m�N� ro����ݛ�(:Na�fg2�w��f��;2��yʨ�9Z%"99����%M-��8���J����8��oX�pa�caS�=e�C�v �Z1�pP�T�&H��π���ϨMi��W���s@��c+�R"@�@�r	PPRZ�Z	{�8�/�]tf&����EWg���l'�ߤ�X�r6���NkL��O��oo�%���� ķ��s��S���^��i�v����|�����8�5�=���T'�����Uu�)::����l�X�
��]��e����嗀y���AZ��h��a���<��`Hdeq��=ggO(Օ�p�͙3�*[	*�jjk�!q�%[�V���Lyɇ|�Ɏw&7۬[����)@AEe�|tFom���{V�Z������>�����MćJNǝ�Q8�r���}�$j��n�z9�����m�Ǭ��+3+v}��_�3׸�U��j�s,j�"�"�C���0!��v������*+�X�`)ǋP� �4��7t6��Ђr��e�T��o���X�	�4a��=	p}�Z�57�:�R��H��8|�$T��SSSw)*;^� �����j�g��8"�M~�SRR:��k�R�$5<��#��5s�w|�����ޥ)�3�\	�g7�b����d�>/*@Sg�#Sm��S�i��8]8�70��Z�N쎗�=	�����8��x8F��"U+�,n����� Q��[	4���G�p�ٍ������M{���#u2�)ː�r�#v�����!ǎ��<���B�s����4�X�JY�%9��
v�l3۪�E�_ ���Z��	�uT���kϱ(_	�pO��,�c�.�*��4ྜ��$����P�,�� �Q��p�̅[ 9�`�����+� �]{��x#��	.����U:�F\<Y \��X��=��$����`���;⻁)"OT:����S��H!qj-���|Z����^�V�����遗��Rě��Y��o����9�g��\���EQ��k��$%�*kB��j�,�fL0�d,�a쁘�knl���lNtqv~�](BVR:E�8�yy~���{ÿ�����FqߟA)[�ؙx�F6�ő'KYJ������[�4�ݻ4���ň!��Q��P�׀Q_�h(u���k��9����n�sju%���������߹s5C?��T���w9;�b�2vO�币\5�"����'�{�4�q�_T���j��Ʌ����<xW���@�27�!ܰ�2���fj�՗/_�z�~=6G��wt����!����1��7{��#
T�i���c
e��t����"��HE+�MT]��BZYӼ�{{�].���Bu���N���$Q|��Wu��*�NUf�"�x��U�ȍ��{Q�7f�+�������5'�1�ٞt��"���A�)z��>�!ssz`� .u��%XOP�Y���z���rV�������߉F�}'��}[��Wc����#Qy���7��s۰xѢ����[yEv^{���E���I+�znn?��wab����WZf�:�*qK�G\�F��5�}��wAC;��-Z��3<����R��kr�6X5&��\K�l��G��GFܨr�@E�.=#���.}p�.55q$Q��@�y*H_��ĕ��]��d��nMMMA����g�����"l;;�N�5�i%9Drv�,�zP����Pb�A��2�1�J�(GjF����.�S���	�6�p���u�7��N���T���4�j�b���FQ��o/^īh�͘�"��[E�@��m�k�Y��~����X�h��W
��8������Qltܒ�3��>���-Q���t��h�F�ZPY֔�n��	[�b�D����ڎ���Hq�~�.
DP���֐�ҥp�ƞ='�o���!<�o�eq���̕H���q����{��B:N���c�&��mj�	�Ŵ��I��]��}��]�Ꚑv%3Qh�9j�D��t�O\8�%IEsS%28}���k)�p�~M�T2�r�G�Jx���,�یՉ*ӑ}oWj�Ml�!rr���zAb����x�x�;4�C�A8�9RQ�7Q�Bn2o�L}���9c���ca��O49����mC]2ؘ�M���m'��t�C:���G!�\N3T�իSSS%>Ö��&1�	j�I��\��gPt���*��F $�GU�=��Vq:_��Ã��:��m��x��t�Gƪy����_����q�im7��Ӻ�J�o�k��|{f���d���ݻ}�
H�4��(�#�}|�� hi��0/�U%i@���������])� �����f����>�]$&��*���j�7
���AK�B�K}=����gFP.�"�;��f�T����f��WVV٣�E�7��k�.���6Ȝ�é��K�8E_���s��J�䁒�s/"�N~�K]?hݦcK����p��9?�%?�߿62B�D��?}�
���y��P�AD�⡇�-��n'�ɓQ.h	�]��
�m�J���6im�o�ݚW��^���㟗ѳ_�0#������A��s�o���̞��>�5t�w�ܑ�@�12u'.�ӡ����p"�d����DBY>l_:���-̷�#n�y�;Ed��l�sJ���|�v^* p�RP��(S��9�c�ri�#�4����5��x^�£JԒ`O��VT�t����l�F��V�G@è����j�i	��������$YP :O���]��bRL���7lW�e�Z#fstH��*n�CzJ��u�&��3��7�𗊦"Ui���)H ��|{ �zV`�8�*��4��xw�
��gLŋK:��߼�����-X�ҿ4Q�..6�&��г�����vws��:��mIT�[v$j:KԦk�>C/��3�#�T����QAȡ0���X����'�_UU)���f5��3�%�3{����H��"�fRd���f�;	�����������}@�귔ym�{߸zu�ڵ�!zZ�����/�s�՝Ri8��uɒ%��xqhf���-�6�VM]V�z��MGp��f������Ȕ����|*�����g����+：�	�P2L�3+ܙ����dfŪ�/�T�`���\鬔��?!PxfZԦ��?"����K
��qp��q"5�!,�L5U�����66:(�ɉ�Z1"���9�EDp�a���~+"c/oy��hNy�1�6���;i�ˁHhN�����O�d�,ߔ[0��<��� �ɿ�>����A����l�BQ��������Dko�����CBu<&;إ�aɓk�v@[٥�n�}���)����c�%]�J#��Z�ۚ8�hZ�����O
�è�~;;L��`���B�C�pjQ�;jMq#>))r����2!LM���.�<��]8N[���5�F
E��!e���*|�.UU|*z�2}��<�{��J�'{Ī9����79��B�Ju�k��chGmB�l��Z����(����]k�l CaE��)>.�?+Û�-!�o�Z!ur�5y�3CЫ�5��H������
E$�n����g�k��Ar7	R�U���h7�'�R33������h":����rMJ�=���9ei��R���p(�z5H�U	z�Mėr [�KC�F��n��(�}��ɓ�.��u���Y�TB�!��	���~`F�
:�f��i�WD���|> �օy^��K�.�X�i(Y.��$WQ�5��F oh���*2�tHi3O��65��/��%����{�?~�Hɉk�:�>�q�m�H���1U���z�\�u���� v�&�M�FI��X��u� g���5h���5��q�9~���Sb}�����B}CH��[�d��/�q��&U+�@�p��gIj�)\���:��)V��*�ѱER�"N�E�5~���d�_���{�Se�����K]����=�uߑ��'�v�-9�ä�N�c�Z�۷�����-�� ��}�sM��H�󑓱�a�D	IL��Lq;���PBth�+�S��s'>>�U;n�u��t��3�����h{��MЎ_:���Dʽ9�V�-X'V˨a-���+��k4h���c�Q��	�.�<��s��q"6�D��S��."Nq�%El�MG��c���K�����Bh��Y�q�UҥF�8x�ࢨ�`��]��6	��<߈駨ج�A$�Pх� �w>�3'�?�%]�BBǸ�݋�����/G�����(����v3�5@]���D��G��G2a4�56����
��񧥥|��q���з�
-k�c�MNN�/ŀ�Ƈ�@~h�n'�����.�X�Z���]2,��z�Ğ����\��#Q(�dddn�>�&8#u^�ג���?�J�����1�T]_���w��s�O���� �7oR6�b�����^'�:��N�Z��#�P���LЭ�ˬ���.�.M�n�o�d����b��EkW��n�����a7oB�����.,#Mu�08���8Fpd�C,k~όq"���5@�T�Q���Ή���knlhh�>}�����$�(h溺��ˣ��6\�2��4u�l���6��h�o��%wsA��&�N�f�s	��PK���V'2�̈ ����.�G�)v+ձ�\%�r�&p�8����Sff'�����ֻ��5���3����p�����C��J�{�q���֖�sr�!��	�T"K��(qN!Hve�i���0V�����ܾ����G'�����)a�o�Z����G������&�T⿨�����~�������U`	��U.�8j=a׮�x-c^L��Ν?��ݻ��혣�xn����b5v�����X������wD����'ף-H+�o�Ɨ!�3(x$�Y�.����6���f�����R���R�;����CC����Ū�S牐��{�������sr^e�Ƞ�|f5փ�j��������fq�[��R��ǖ�gMґ�ܾ��?4�StŷX�Cm\�g�|������	�|���Th���}vz""_��&9����aj�)R���b<��>C?�x_n�j�s�b�24 l�0 �T�L�Ω�w�T@�'�G^�+O���-���^����kD��{#�����>�G�@�-�t��X88����~��5B�q��_�6���kB���>|� ���@VW��I�^ F)�j��HJh$�y�U�JR\:��a����B����5N_l���J5R3Հ
�O������?�����2Nx?r�������(ť��t߀�N,}'��p�xg��VXJ��=���Q��~�dv���lE�QE�TG\�]�@�&E<�E�֯_o�J�[;Z-�xj�9�RZ�7ć������G�l1�z�nS��7�j,^��H��a�z=|�.�tH�:��D\��e�޺uKU�e����M���#Y�����+�.�gB͘�iv�Ӝ[�&gM�3`<��[[[I	y�K��k,��3�_���'�j�u���Z[-?��:�M��|݋���+4u��j?"d��S��	m�.Lp#�u	�˸��}jj*τ%��]T���˺u��恎C��k�*��^N���S��N�ݱ�\�i6WxѲ�GDQHR�	n�|�D@;�`:��|�c!X��V8wy��O~� �]�o�ћ�i��U�����[C!�͔P�n�kǋW�4!B�bi�x��̤���=����nʭ���6+>A���&1/��9��EB0��;pI�{�r��}A�P�e$�Ɂs�f8}%<����O���i��+�/Bb-d�v��W91��9�����!P��
�F�k��l<������"!	]-.>�ok������'?��j/#I�>xff�xF�[�.�DC:��S���t(.��Ҳ���+Ҭ+��{�#��0q�bݿ�wW�LU2�u�ĉс\��y«���E� .�t�F�X�&�fdfZ��L~�]��KA�Ҙ ��klFi��0���&��b�`�ڜ;����>0��f���!||�CO�:��@�[V������o�i�43df$�<�E%2;;'���㩄Tp��W̦#3�<���qF]H�6Z�{V�1���!s�s ��#Q���R�_�L��e�\����(� �(20�8)(+qr�p2�����QF��ܻ^�/��2�4�vp�J�4T�� ��}y�X8I��0
��������E��Һ:::.!�V5m���'����Em��j�ά���B"�ԺS�j@QUf�	�s[e Y!$d�Pږ|�߆:�
�3�<�1�5��BVy��u囲k��� �#fꚔ�p�*d��V�D�к���cۻ$�9��M��sP����q��#��[ը�L��1(���m�S�J��&)�Vk��L:���Z�=�x��27��i���		ھ������H��\��ƾr�J�95 r������J3�>45]7�bq�xYV������ގ�ڕ*Y^`�|"C�%v�ŋ��aЌ/?�I��,���(�K�koV7�t�fq����K�'z1N^��_�K�T�)�?�(��}N0�ZLl��d|�#T"��ŋ#��4cl���D%&�swB.q�F텲p�
0����(OP���״��m�g��c�������j�T�[��w�_��N�$�
xZ^��u���V�Nb���!]}}���QA�,��9-h�F�%�`�Bf�$��  q�S��7{��<����e.�לhUz~s�Tw,�RU��JHU��}6��l&�_ ��ԩSWKKK�R�;�;'<3Z�����Sl�� ��vT �D4x�6?&��2޵sgm��V(��==�O���C�|��C#��g�eC����ތGH����9A��Uf� �c!p�-n,Y��W��2��V�������
 q�~3�z߽;�F�~	�L����q�rn�j�鬉�wB�kK�R���2������(�l��_T�*?��C.ke�5���$��ZZ ���p����1u������^uj�R��Z{��tv��L�)����M��<�'S�|�#4��7C0�dی����8Q�W�v,8�����ƍ�b��p�zzb�r)�io�Pl��
݊�c�C���I������>�R)h��!�� �����T���c4���DՁG/�}iE�S��Ӎ�\�_AV�f�L���qsۉ��l�����$̰�0�%��I��k�UEZ�!�+�2hm%@�}�;�[��oܹ Ҥw��cv�={6oh{���Z"2�^r���@	:::d)/5������C�A����
������
�(C�mp�yfz w׾}M�Uh]9���~�	d�q
c�~�^�M8cS�7fg�WA���&�(�����z'�B���ljr�s��ZZ�	D�ײ!����7���<<�d�`<�-�.�~#�t�#���p8��sA�`��k��<b�?�1Հ>���!	]EX����"U��a&�V-�T�pǕ�_inq5����ߓ����Ɋ�n�T�F�ڵ��n�Ƥ�\�q���n�,hQSU�cz��-m`"ll�*��}
�3�v@A�^��v/��>�d�d��G�E�{�����LN�%�����(��~qI�b�C"�N@(�/�d�������jM��)�z�.��ڬγ��%˾�jxy�F����C�7��ǥ�����V$>j��$O�Xy�rlOg�����Ws�s��J��{b�9������5Į�F��v�D��Dل�KL� h`|�3e�ЭsVH<'����Av�"	�j����;^��Ƶ�a�	|�	G~~��=�0ҟ?Y�,�.7����Xd;��MCN�K²�2�/��n�A����3�s_��J��J8��Ͼ�3��gB��u6�S�RL���ԙcW'ck��m���Y�d�k���� ���B��Y�f�R��99� 8�U˄6�n�$sy����X��7q���FZ�-��A�Q`�"܋�Rt��n�x������@��M��D�P�b���%K����� H�5A��ɪ��Y�|)ܞ♅yG-ɵ�l�'� �_���3*��3q�i~��nE�Z����%�xd	�[� O��-�Į�����U畗�u�����Z�Bk��r@w�7n��n�읗쑨;��5:�������f��6] �7˘�N������Υ �L%�M]B�v|�������BSUn�p&�ckk8�O�D�q�:��퉻�*ב��2�M����:>���
7���"����7�"�?CB
�mM�]\PL&%EA'\= ����FҡJ-���h�׌�:kW��mW�nI�X憸q9+�2�j�qI���,��d�gB�0QWiE��_��� �6�A�ٽ�hv.�2��j</oT��9�2���Ep�o�1�匰�	���О,���TE�#�LB)GN��������M$�BO셸�P�6�x�1mI�Ԟ8����)�ە��j�����)3��S�Rd�Q��p�3��Q��W8��iǯ�-����&U��8ea��-(��ړ�Í��׬�2Sr���5�+��y�H�L�܈N/]#��f���?�Rջ��L�)(���ڀ�q%�(�c����<ɤv#���t��|(��A)�R�$��T�F���ف�5�6�~c8�"�� �$��u�4��u
��'\�����N�7$�y�������E�)W&�py
�Q#�V"�U�4N䎿!I�Y�����E���d� |����xr^H4��w�5�Z2!����u��i8��<��ׅ�o��F�����'��\=r��%!�Q x��M�pG9�7�W��Ȱ̭�H�b�~���^P�-/�b�ƍ��s��x��wB�#ʶ
	���@�:�N���ϡ���ȴ�������m�ۄ�,k�X�?��F���N��<wF:aNkn"&5ۧ�m�Kh�Ϟ}����ˊ�Q��z[���h4Y�!1�Z�B�ş������o���,E��E)e���.Њp<�z�9�O�	��60�"鮉=p'�)�`@M��Z$��1�@�wB�q����߄=p���9I�<jg��X��z _[��s�O���x�h�dh����ʃ��!YYA-�r����9�+��X������
ߧU�4� 111��{A(1B���c�0B�3=�Us����A%�Rhx�b�L��.A_���R>����Xx8�SjN<q�`8�W�}��Bכ1<+�?���>�hH��՞�{�O��7m�������&&�W��(�oO�g�����f��c�<�U����fѫW��s�*F��<����1m���N���������C�U?~gQ�k�ѭ�孠�C�m�"�����*Jp�a��[��7�ڰ�g(J����M�%��V�kN�G~�����S�L�y'��lM�h���I�t������.b�}i���h�F��T���絽����G�|�hAǽ��/A_�8��ʖ-[D�^��2e}��Ny�ʰ���!��???f~�����t��~��2r ��1����Fg#�,�Xgu�V3WZ�pm�$\�w5e����i�A�F������o�4��f��	xe��)��A�L��(t�2O������{�1�%���eH)b�e��\����N�ŋ_�^p�kw=��K_��pN���Cp�eXX؁ȱ���z�V�L�̚ǜ�����H���57%�>;�����3zV���E����GF�����.���3�6�ˁ�����H�_�Z_X��(R+˘I��i|Q���a81��B����r�w����}<g�Q��e��{��}9��љ|�0H��U]"ɇ-��1��uk���)��d_�;��׽�C�>���⪏��37�jErU�I��]����67p?~<3�-f���ha�|%h-��gJ���V�J�,P���+
l+M_}����-�m:*�l��#�XAk��l�<T�zµyLdWz�r���
x$몒V��A�6�[�����gV������q'��-P���	�K�� �ٓJ��Y0�+m��L+�~M�������KbO|i����2vqi����'n;+]�ƳVY&������{��r��Kǥ�������[R1?e�G�}�����ܜE��?���d˂�P\j3�P3<�'/�4g[;/��Sz��x�!��'�`���3��C,�y|u��WNY�����ȭc����������6+�hȾ_�'?��?�P��3����2���ZN�W��
�D�@���}������V_I��3 �C��> �`aԙ�k׭;!����:���K�}�&��{������T���4E�E�	��*�[��ݺ'��m[ن;b}*%Z!۲��_���lZV7�U�⿵{���ѹ��K
���1/�#_qt�=��i�������S�K|�z$S�}{�O7g��6T��gܪ4��,-������_��}����eDF��v�G)B/Q%���֢�ۅ�!ML#� h�;VZ��ip텠 	f���5�c*wӏƍ,E�|�vZ�t��6������n��ILZ_�CZ}�}���e���E)�8 	�������^Tu�m��V���~VV@ℊ~��F���m|��@Gq���X� bҵ�d�����o���ɋE�i�\��d����^��)��߀j���2⒒�` j�*VU�{��x��e=�G7�z�sQc���;զ�A�e_T�S�$J@�>��ߴi�s�7L�)�Y!���_����z�x�JNWWO��ae�c�(����Q͹Q��d���a�1h����|hy2:x'�-�K'g��%�uRz�s�>��+�����c���)�6�šϑU���KB����CT�]�ee��â�AU��Bշ�tO �AL��y�ZU���
�8�v#*�X"5�/�	��lVCC�9�ut������'>�{��9`�cR��ѽ�oa���B����V���ϣj������ ��Bc�Q�H���,�9�Ue>�%�Ӝ=��q5� �t�X�0�C8��7�����Omz�ۜ�2��5�d7/�a��/���XYl�#P%2c����b����P:O&�!��b�Sqf��T	r|�Q}CCC�ݥ���-I/ܰt20Y����m��(���H1곹�������GfŮ}\N�XqMk��xBR%eee=S���6{��g�c֩[�	��lᘊ����#�������cd�����%�5{����5�͚��Y�l��
��Ȫ	�
x.S�Ͷ掎���9WW=$�9���B�h��<��!���!N������H�U��-������h���ր�D(eF��?�\2?�%��Ӟ�����j-�AZD]�r�4�>'����b�'�d�f�ɓ���X��_�8)��XWTT�ɯm�������z�}j�М���:���¥߄����t��珏��c�x,�/�1�9V|�m5 �)O��*4սr�"�5W�
�
9�������WN��wԷ«/��58������[ /х���׿���*9E�pߩ�]��c�����O��ޘ���~B����De~����S ����9������YOy�L##O�HJ���H��g��Y�,qnn k`Ph���..$�I��XƌF��U�0�<�G�8A�E&�z.�c��1����p��c�9{tO�ٳ���N�}�
r�{�����r�fP����~i�ˢ������~|�67�"Lc��7o�$���]�]o!�6"xϝ�0nsP`{A����P���W�1A���GG�~`gg7��0�Я"ө�����5;'��M���+{9;�#��VO�ܧѧ4��?p�n~��%ɸ�  �]݉;���l�>��\�U;̏)Ļ�s�⺔�jk��g�s�|VE@�����غT-� ��wo����c|����+�q:m��� ����Qq�!��X|͛U��R�8���rx.��5�J��~}do��y�"�c#h�{{=4���P� k7��\��4�����g���$�X�ӷ����q)"�m��C�Q�v��#9t�{ 8$$��IA���ƛ]�ܔC5Qy��JX���o�ud��h*t2��X� ��鯥ش��'	�%�ss��xA 5�����-���ܛ9z�;������c".~~��EdF$u'�_�#w�Ki�{�o@���'����kM�~���t���é)� >����V�f�1	�/��I��ҩ��g^�U�y?6�O���u�I�)�O?��
�?ܽ�f�E�Ϋ���
K���C��G���L--!I"�,z~��)T�L���:�;^{�Z03��6T����[��d�}�����p���i)�3�f���䕕��3�%���@7�u�V�"U*
��/�?:��i�ZJ�������0��t�2;`��i*TMb{u��/�ʔ�5�?�U���Te9@�UE��ҁ^^^�jN1�
T�mmm�H�P�-���0���{Z˼t~��'�r��c`�N�81=T>\PQQ�3�Y�֭wP�Ba{����a�,d�caS�~��7�T��g�]}�\ܾ�_�a��`c� 
����e�Sy


��C�8+�1ؕ��9A�\=4�f��n�Y��bv匜W��%c1���H3X�Rs��㍣�`��j��}��V����;���w��2����V���V:lN�%Q��RQ���19��Oٲ�!$!4&�!��(E���`0���<����P����������_�l�������������� ��tu	��M�j9=9=33���F��?է(2*9�C�F� �A	C���[5.��Θ��vd��?_f�}���f
����*�U^ً|w��}�w��'e���*��4����weҎVz�8xTI�y�zd�9Pe�AUƹOh�R^z�I?�3�-���4�� _�ŗb�?��xb�
q*jƠ�41���UWGq�ψ՚z�'00�TJ!̆��1c�Ur�A�J$7k�7�«�C��xj��U�'��Q�6��-�toA(�����Ը^%��I)�Y_OO2Հw5g2�Vr�'�*�ׯ�C����j���m�74ըI��.�3�T�Ȍt�X�I4�[n�H��_}h���h���
vZΝ2�������+���m>~~t�&�úk���uq{9`�Y{��C�������A<�mm�=а $�F���Ǐi.��!Q���������<
��.�<!���aRS�������L��R`�a�8nա�lY!��(�m����-Q���Q�U��BX
�Z��%�@���RZE��R�՛Y�_��Ga2�ȥ��rroBNp��w��,(���y�	�B��Z�D��>�?��I
�(���u[*H��}�US��]�������*�GJ,��N�<8�Z�z��2�����fK��|3����Ej�FY҇�G�G	��	d`���R�b��y�!�[�1�x�NUj�Z��y�'���9q�2�UP ��H�*4x|��άf���8@|�Ai�Q�l�i]�؂�f)��ԃf]I�xz>�;y}��Ǒ-kx�����6N��Of2��f�kv��d�k�A��r Q��Z�������B��zȂ�Ѓ�7�6���
�"�Zi.�e������Ku��K�.�c�X�h[K`���ONNV�d� � G�f�Չ^�<���`���p��� ��䙠��s�/���e���H� R�h����%$�0�N�����b@a�W� 8t��v��s��(�����@U�L�����8 �U��C_ݙzR-�x!�2J+Xʳ�!�'ԽE�|#,�)��Z ����~!>)!�2iot-ѧ"�e'۬)m����0Z0['2� ��]���j7k�KQ���j���ՏQ��,��;'TBJ�E5\H�`K:nd�_J�U	��}�Ŷ$PL����(�(j��%4�'�v ���(��s�k���P��?&A :C%���>}Zߖ\j����\y�2�Zmmm3�Y�FY�N�C2�TaSס�C� n>%�5����*p]of��������n�V�:��ф�ڪ�Z�¡� �<xpx�>��/�P�-����wC't�h�Bm��J,�R+q�$�
��Lp�({��-a��enn��&2����G��گD�_���ylU����t ��@��sh�������<�������bb�5Q��J��}uq����s��N�}����3�"Б�ѧ�:Zeh¥��6!�}�H韯e ��P ��<��R~˪��i_�F<�ؤ�~��i������2jc��TZ�-�������P��~��L����a��O�8 5�S�F�ŝvS%UU�`֠ܬ: f��N�R���d�]�B�����N̨�h��׍��6�Y5��x'Zw�X� {����e��o�n ��}��]�!X�s1쭲��/c�/�+(E�:��o���u:�6��t���4��&��3
E�x�)$���D强��k?[YE� ���@kL͍�&���4ܵ�݅����D,�WPȆ.A�B��c����F��F:�Ç���H�,��L@4�9�zS���C>�Gj����[���.��{���7o�xg��m:	J����jU��X��P:��{�O����s�?�EB�@���k��}fFZ���*
����A� ~b?Y�ȇr�M���Z�AYu����Yn۶Q� �,4̤6��9C����W�`��U-����{�S��+���r<�D�rz~0a1P�CY3f�م�H뻄k����9����)�����˒|�6�d6=7�=�vXkσ��gV��sj"���^�j�{~;+��5h�V(����D�lNe���J<��1C�%��ܩ�����2��RQ�]�Zv��ս��SuŌ��v[+ެ��L�ooGLS])�l�̞m�s�nDD��'y/<��f�/L�^�����?3ܐ��|��ͤ�w����D.)�w�����X5��nr`��ީ��p�n���ǪJ�KÑ��Y�DL�`���_-9��795���۷7cpW����6�?VI�g��H:**j?��V�%��Ol�y]����h�����"u###�ih�|d���2�����	�1cjH��U�^�sYs]9
�T�C�{��ڵS '���~�V� pn�c8D��k��J��ܳ�"� �nܸ87~P���:0��6��Y���2T64P�l�����`՘���m"�ܞ��&�ƧK�!Ս����/�srJ�	@�;����U����5P:1"���tM��g!�Ŧaˌ���/���el�/ P\��zzH�iq�����1T�ݭ���GF>�XE�������j���PN���V�0���y�NE�2޽�|���if^~�������Ix6#��`������.�a�7����tF�x¿��q���:�%>��t�1@�D#]S�R��b�jhp=��Y�q�RՇ@� ����8��<T8�|@`4X��k\^yy����3�P'����g������r�-����fb��J��:���g�G���0O�@��͛��.��bOOd<����Xg=����'�w��:8)\y��пM�B�;4:M$�ڴ���vp�$;c���]]}��x'��|��!J�#ǃ>!t��҂�����=8-�d�B����+ ]ez��>�u���.\�h"S����!�C��9�P!I��m閖��r�s��~Y�u��<�֣f�����	�Pq�|ɜ��/n��V�U�=�yt����b������}4c��C��.�.������ԡ�L��(�2߿+�vCVJ
\���v���Gw��mW�jy`g���Ή��GP��i�[�kxT�U�h3�H!�L��9��J��3��?'���8wz>�z�޽7�2�9��n\)�<�n��S��!sݱs�_�?�_� ��!w``���q�.��T�7��D��[*ξ�	�mu7�>�)�%�{w���H���`�+._L�� ��C�|!g[�'��N2��'y��ݿ����ͭ��>���؃tAX���Ha�0����M)ĉ�����%�}���-m8
aL$"r+IO���-[�0'�::�J�zWP�Z�5k�ق�����Y:rO9�F�@
uDH#j�3�P#bX`ú��=H���ڴ�D��Y���-�Zr���d��/����X�����S�������YK��!��1NHHׅ@+�D��T`���d^)��ƣ�/u���j��ﳜ�y�YU/��B�O���s�r��ٳgU��y[��>�=,sh	vuׅ����2.!�4aAc��r�� U�*���=1Y��'9� a?�{E�y'v��3[[JKKwg}P�Z�'=��s,�i��UK������s.)$�zY~�u�8a�X�n���H~�5e$��f3b��T�j�� 7L�����V�m�<��אg~uź�@YF8�|_��L�����@:������{��kG��f�Y��b�b0%je	k�^��Eꭍ9������P��QŴ�������ڋ�����g����Y�莬�2�(�-ح666���d68AlwMX嘛.1��� ���!�ckk����%�����8?�X���`L��!A��1�~��A���ȷkG�	 /�X.A,j0vR}=�X�,�O�n�۫&)�n�:���ܻ���\]���D"����|�]�8k@��T�����ذJoϠ�*9_R�~�E�;_?�!!�md��	֬}I� �@`�J��/���S�'q�V:��>��R7�b����.NN�7n�P �����܌��IzO胕7���V�!�{%6ԕ��W�=�� mR��pSj��/@�!�_�<
Z� �t�f�*|�0$�R� ��\ɦ��RZFF�����v��ȡt����5 �e����<�H�V$}*����c�b}�,m4mp�z��D�M/��UB���3Y�?���� �������{��*;Ҝ���4�;-llH]X?Li��7a������w3.����I���T3��q��u��*���g"aMI�ǻ�&ءz�,v���?Ӟ�h�����iƹs��f2�K�8��`�� �I�X/�y�r<��З��'i�A���i�^���{Xfa�I<-˸)UՏ��r� n�,��$�Dי�f�`9>V1&E�����%���مN�ȸ���$��/d��������226Ʒ�=����d��쬳��)$d��{_�; ���Xh�D���Ҏ�4�`�-OD��w��b�R�=�h�>�p���'����� 3&&���p�;[~)ZS�ӱ����.q�ϫ�Ӆ�42օ�b�۞����/B��YSs��e����]�<=�8��q��C�����w�ۭ_c��o֯�9>B�>���U����ps����G��.$�xA�ө�oL���U�^lJ�,�`���ަ'�΂ȓ��3��mDl(G*���q�J����R���Q��ʠ4�q��*���h2��^�`s���wW���*�Xl|�}�Aμ���d�����J�fy���3Y%y���Wa�??���a�s�H<T��*�`���މ=�K����K�3H�������q��j{>�+�#��d��С*��J8�:�"J{�[N�Ò94�9; I1����&��BAqh�W��JKWN8�b���eX�ѵ�S�x:� g���;��q����Ȇ���v�ٱu�&�+a��q�Y�T��J�kԁ�BƷoO��}�Ť�R��fł ��C~Ph;��	-F�����7or���t|SG�b�/����"m�5dk��)Dݩ���k�9T�'���cqk�#��*!ZJ��e3t�|@��E��[�=�(��4�T�CMرc��݃�� 2�|�7���E-���T~�/|��R�P��lg��3E�)&:z�3��E�lW����?�IZU>U��AC�?+k_!l�j�����R�'�.�Z>|��#����0�G������dƹ�Ϲ׻g{Br�O�y����
���:P�f��o�'�������]�'��b��\���"�Zݽ�9G��=TS[���C���:[�I,���ܼ	��W���!6k0]�!W�27x�ÁͿ�ִ���N9Ě�ۊ�({'|�ECaH�:�����,$ࣨ�Ekkk	�\�0m������	4�Vk��^_gW�D�(����c�̅q]!�O�z<�x�?���~-;��@@_��2�B0X�5���z����o�9�^\��� d��8������ �E+i���mRx�B�Ň���=7���/��>QlHc|HX���6�l�[&=�L�>C�v�gZ-�P?JnѤ~������dr�UB����n���� G���k+��xv�}T�,,,|�ZWW�����]�ڑ��N��ǟ�8;��s�κՔ����q"o�h�䓳�}������
e: E�BP��i�Xա	�r��~�@퍕����n��<'��#�W�@JJ
}���.��l�Z��H�h��E��v����	v�*믑U?Y�lŪ��㥥��9�
�*n��#B!�EP�wf��ː8�2&�!*A.N��^�1�	z8�K/�Ď�b)(F��b�� ��M�=m��F�yK�j�����-�k� ��N���x\����-;4�C,���[�d��=ˮ���pK�U�5�f��ҕ�̀�G,���.;����'dO^�{b��e�1��Re��!s�6����G��I4����<��LW�����V�=��� B���Xd}�|�Ԑ���;�����{��5����W��߃Q��KKK5	��*��פ�]�l��o>���X\[iW���܄-�������^����s<D1j3�0M�鱏#~���'~��2��^<�d�1�-n��G;B(faaa�A�*�	nS{3��,s/�A�khh���xx�b�W��1�@d�X�E?wt$�Q����1��GV����,���'�������k�m����o~�F��H�\�G����>��O��6��8�ߑ�H�3�}�nD��{�~N��[D�~5/W�Sx�5r)XChg�b�����g(ꉎ�oO��sW,�5��6/0�ӥ�X�0h�ֿУ{�3Bػ�W�2�Gw��[��P�ʟ@�=��V�ZݱL��5k �
 y/!��	�g{u�A�����'Z���ީ=Q�^X����"S33���["���wN ���Zk���E���"�������t@�Wϋ�J݈ׅn�2^�}Z,��W���t�9ͲJ��D��%���������ݻw�U�	�����tuu������
~�~����G�s�����ld_�ku��L}���o���>�g�E����633�6)��\�o�M��E�ʗVZ&l��s�I%���N":�0��"fR{f�O��La�Y_���z��D6o޼�Mz��&�N�����CO8��+����9�����Q��-q9r�)|��ʭ�g?dCqA6o�mnLa�%\V��g�r�^r)xնg�'����$H>����L�ӷ�E�#N �������EF�;����}� >����v��}���w�=��F�D��ps����(����udĘ��]*��x��Z�/�5H�aA�3r�QJ���V��X��{�h8~*�U�jY5c��=.�����<>����T�|G����U���jڋ*(pvs��X�h�����L`���!!V��Qn�QM���g�El�z ��En"���*?�1�{��4��z��D�w'�l�/#��)��R\�C����
�;!�m��yV��I��s�~&j� cdu�@��C��֫j��[<�W�'�>9�rҷ��(�7o��<���<w��	$��2 ����"������J{rrU��_��oA�d�<�r�I��F[[[^N�:T��i'["��"kb������n�Yw���P�`�[�+��&�?�{
/�����j�w��As�wt�+j~%ux�5���y��V����kv=�~w�pb	���4�g�E�똕�R�Ђ�,�~�wYt9���W��DI�TM�TU��p�p�����!<��~�H}��e�w<
�Cd1`)� �,<l��{�� � �x����BV]��0Pom��0!5Ig���ɚ����E�M$��h#S-�]0�o�z�J�h0�z��CD�C)�J�p�U�������PD�P��HF��6ke��@�̺mdg�o��h��fTYc��Ǣj�[/X��1�hWr��U�&�<�z��Z�KHHH���`$O�?�~�u7ci)��/�?V+��}(�cZ�]
hP���OC]�z�ָ1Pmt�a��Har	�6�gѦm�喋���8�ѽ�N�^��o�2���Ntf��h!��
� �/J�P�����Hm��m����j�W^��+�j �j�v�)S1#�y����U�'�ܷ��}[�) ���}�����l��i��DQ�ט���i��]�M��ˊ3�]S�5�Dc��������Onn����9�' �PO�R�V�w�� �o+E]����8�����ё6q�� x ��@|`o�W��i���n�x��<�P�>d�+��HK���̜��3�ޥ�Z������Y�!6�8(�����M�p���(��Nf'?��טzR�FGP��c�<'����S�&���Θ�4Ͱ����n���C6�Ц�QSx:��D��n�'�f��g7�K�K�$G~�N{���jdf���������^���������(m���Z�?�VTO��yE�	D��&�����l�/��%r��-~fU����O ���@Zm��w�&�T2��^8#DH�M0�[*���6��{E^AŃ���sm�:n�U^���������b����t~���C�(�3��?�M����+���%!.^��� �(��_<���O����|8'd1��:��5hb�W/Cֺ��u� ����9�R��;vm�SDj��C=�:T�n�(���A�4:a�Q�<�C���K���zj�"�l���)��y�M�/$�iCK��E�0�D�yB�����(ӷ�!����^8�EKK�(���24�>s߀��dv� �et�ֈ���ef�M:�.8��Hµ�,bN�����ߣɱdK	��P�YYA��u��g\e��JJs|�Q��#i���#�3�t�j���M������!�!����м��Z�M�i��ƹ��Ad[I�ʃ�� ̅�\ɡ��T�w>��h��R4T��ԙs]��X�4�M/+f;!��1�	�\���Ѓ��v,����E���\�֝u���Z���~[��~�*�<r�:��	����Ӆ�����6�-��p�v��`�?{�)�����߾m��%�z�u�w�����O�oX+1ao���H����ȍ��ڪ.�z�7��&c͆*>݌%��痑�/�z������h臦������Mb�!�惛'^�4�D�GT�P����+gS����A�o�$��փ~��l��4_�nUY}t4��H�UM�ު�Ws����&#��G1!��K]읱�(��x�u�f�y3�Kc��v�4����􁹹��uW�v��3����g4����sX����?8�0��~�H��L&�Ҙ�g��)�qZ� (��1�N
����=��,I���(����tx#���ӳ�	Ǿu�*YD �C���-��IYC/�MOK;P���ӿ'�TFN�f������y£��s�W����K��eOx�B��ҟU�Vꌗ����#}&p���]#RSS+g;\hR���	��&�t�cb�/�(>��ǝ:C�z ����Ü���̕{d59>�F_l�����4��B=�y��������|||^���x�E���Β��_�&��s�_/�J=�k�ܮM�1aj�r�7���'v��"�+k]S�����o�3��ծ��JTsI�~ɚ��%��r �0=��5g���^����� e�
I���R�I�'c^��s�)[B����՛�zì��MSJ������W:��9g��aUUՀ��"j������sZ��Tا��0�O���Ŧfff
	[]JiD��Ѹ�՗Q9ŢBB���4a$�Gi����Gw��]���	D�a���O79[��dg\wm�u�8��vO���̇�A��v����W/=p�m�������h~������Yb�X�5��p|����w���N��G9a�}5S��� i��e7<=��}�v�K�|NN��1�ʪ�D��`��3��۵��q8\d-ȣ@\wv&��\9�<���� {�v�L�[��Y���&&vj"�2��������0&&�	Qi�P��tгN�#8+�r��t��gyy�]��c8�|$�ʠ˝�*�ڞ�ե�$�<�� �G���$?tuu�����*���Nyy �!�yyg�H�g6?�ņYk.W`�)�°#{Y�/U��,���7�B�j�7ʊ��SS�R����#�]]��k˗ao9!>��=��DVu�}��2�<���3�&ǿV�Y٠L��f&�u�b��+2�y2|TR����dݭ��:�����~i�K5���RVR�'� �{��-Qa�Y���Y�	��Z<�;�{��0��g�q�~�����,�Aat�`���չ*`%	�9�L�+
��U ���D�T�#P��X��/t�6��V�&.9�\�����Pl>0`_l���j,�L�f�"uФ �ج5:�$�{4��8<�ٸ]�Ѯ%�n՟�p����Z�}"s�=r��������9�Ο��^x�����t�������H�~s��@�ol�(p>�6  G���Ȱ���Y<�D/��d2�<6}�����[��(�oe�`�9ͺ9�uZ8ժRC6?� YȆ�+N~�2�2���l~��i~��|��W���\&���@Y�ϓf�lbe���2�>��6Cs/��,TV����Q�.�ΙO�'Qx
��s����/�;��x�5ZV��fk1 6�E�d0�`"1��Pk�0�� ���)����X��3:xi!�����NO�@�������A��e)�U�N������+�����[ ���JP9?�+I��	G=Yݏd�kznU����������?vK��nx"ܰЏ�K�޿#R䐷��9��^��7_SI��K�V~���Ð��pU7��`]�İ���|Pĝ0�x�N�����&&�q����Se��3�HE�A:���,>5�W'�x��?��i�h_�Pd�������<�Jq;h���~폘�GA�PVV���Q�LN恐��籶9�F�b}�7�>��R����[}e���m{}݆1�*���*GQ\!�q�Hw�HYjwh�5��H�)�[�a�ҵ��u�>;�����\�&���:�#�˃Yo���z�L�>5���s�9�B
��t"�����ow�l�1B&�#ȡ�.w������@g�)+Rn��`��n�K���a"��:TK�S1�)j��x�)�:�Ͼ���c4��I�kUz唬���T�0�!��,.�*SH�-J�6�'���@�候@��ݒ2���WI�761��OL�i�,X��5�⡒?��Y��0��1�ẹ�����H�300�
L~}��9 �t&��h�/�mw-�A�E42s�&�j�$�M�{��J�|ͺ�"Qa\�)�\��"�i~�W�Gps�|��EP������ērR�>l8�x��������)��KƱa�uC
��h��&&H\�"�����ף7����f'�@�_7d������s�R�bBNr�a���-�O���]L������Ǐ�5�3�0u�w�P�n1�>�Z� �@��Q�[�$�ngJ�|K��Yʆ��P1K�x=VV|�۠��<k�֌�Ӊ��8R��  r��v�����hbz�Fg�4�3��[<k#I���[ϵL�:1"��Xу�I��Z:���ųeIN� !h��kgn��6�oO��+#+RR�=��������`��<�X�ؕ�����	��u���E]��>f�@Y�m����9�މ��yA�.|�z��[�}��.����>g'�L�g�bD�xS6q��-M􉕕��2O���ńLM�+�xA�����W �;���8��<+�Y�ҟ�T���a=�e,��~�"��P���?n:v�H:L���f��N͠�Q~y��$����G��I��Ned�, ��1��Yk@0#A�i��/���ksvr���Ҍ��F�����h��be��^]�0�:�3r��B>Vj"����V��1<`���fW~�]��T�� ��I+#���㮞�j��C����#�SGRX���b,�#�	`$�� ��r�f�e���Nj���	��MJ�{�/����㶗�<��ڂ�ܷ�ʹZJ���%~(Z����H`���$$$���#�mM�ϐ��Rԏ�\�5�����]��߲�&S'&�F�q.�����|���q�!�5�ަ��2=��#c7����qT� ;�{?).���n֝Ɛ�-�ܘG�<����w��2Z<�,����ط��H-�`Cl���5��1��3���e�Ȏ7��q�����!ͅ���v�'��l>:hLٗ�Y�OL�}�G�xғG�0Ca��1fC�B0nҐ�sԟw�7T���.�&�����x�GpۦG�w����t(��a�Y����*];u�W1�K8�+s�44�ꯇn��i=;�
+�ۯ��l�Lm`���IX<�����`j�5	����ԉ\C������&��D�z�S�Me;�%�AC��:y�*z���dc�$jT�E��yJ|���y�85�tTg-cb�.��T�&?~\�����M���)�u���b�L`j�kB^^�%��I���9T����ҳ�e�o�=Y��'�����5i���a����9aERVW�oo7_`��qݨA����(�]�>;c��k#�n19U�p�0�;����KVrv��J���~�h�Z�j�9���N�g�a�}�����Bl2��N4�Ѷ�?n�u�����8���z�#s"߰.z5�e�j�:�.��l��~��ݚ��	\��J�a����̀�Wt��S��{�|����zN�c$8\� _-|j���GO�ʙ���;L�����.P+����L=mP�;�&Qg��^+����?W`[�����M(..��AU�?��|�fG�-P��.0`��o�r~��� d��e6�>x�w^䪻�bIl�Q��|�%�e���C�(	�M72ʌa�ȁr���P�$Wy.�[�k�2E�����ى�B�|To�j���˞Rw��_��+�b�����6&-�95\��d�,�	�~{�0�;F?�I	�\^�{C��Fs�i~��G���[^�\!��摵-�1|��l��C�Ŗ%���&L��u�~�$��Ur�S�Y��-{޶�sݨ�����hV2�R
�����؃>���ц�-k����6N�����{��kHeW����&�n��
��JX6C���V��D��j���uW$�����L`YZo�'Ž�d��y�w�r����4O�JBI58��WtQZ�;�/[>f��ivb���?�h[�8�Xk���R1�pv{'�VTA�nl�4�׽�J-W� ��cc�]c({�䁫E� ��������1��Qd6B�l,�ຓ���Fjj*�{�m�:�-��uU .-�B���^>�q��
��R�o'C��B��Aڡ����3]zG$4t�õ��Cd#r���qsϡ1�k��컫כ(o�re_8�E���_�c��A�*+)�F��(L�ԫ���0�o�Qv)�i �����k�Efmnn�|�t��A���fX��n-$w�:��'��P,�e�i��������v+�LI(��{�� s��w�-�A��	!����#�]T׾YU*�Ys�� Z�?}Ux$?�������[Lo\�W�L��z�ԅ�.*��?�HD�� �~gU��e����j__�6_r� �Sq���,W����8<Z	���D�b^@�����d��T�s<���K�N�%���B�Z�W���8u�hJ}�K#I��V�\N�G�B&ygl҂SM�1�"�Q;^���l�����T�Y���0�Vn��G�-ϩ(�4BJ�
�s�կ
?�[7����Rq�Yߝk���R?~V@����1�0��v+�:�u\B��Ϝ�u�ѨP��PS&!����>����^݆�������K9���u�!MV#Θ��C\o�4��@F�!�Ԛ�L_��Dy�����=��j;��ֱ�u�4)��!�,^��� �Ӣ�:��f��� K�7��~��@�� �.�.W�=i���狭ь�AY�cv�p��&~.ed٭\�z�<|)@�H &�D��yj딇F��\��dbA�l��w$�l�z�^�b���Z��iA�e6/��N�������iC��oΎ��-F)v?O'��o1�V�SI���Ԉ�&܋�#
��j��	�:�浺��f��`�b��ߘ���V.��Z �����P��L���5�d1�$٠7���*�&'����!ӄ��.���I�Sf>Q$��V���cE�?���8���B��un�U_OOO��dc��<!$_Q�;�Hz�"67���3�0�>>>0dE})�&�Fс�*z�Z,��}[��D���э�"����a0Ôt��(�\{�Bb|��~i����X,��{�K�0�>,6(~�aܢ���:����b�;������-�r�vf�PQ��[?����g��H1�	�Y������!�3�����y;2�C�.�r�K��h����&	�K8�ŀ��Kȕ��K�`F�Q��6ZH���&��-��ie-�K���e#�1^�7
.x��ƈ.�[~������f���^��Toe�3�>Y�j��At`k<,�qB���t�٥��^��r��p����櫪��>��|ɤ����;�WZ�.������:�̍���d���NO����zK�Sb�{=��1D�2��K˱��n�/�h4L�R�z�3�9�0?�B[6�]�/r�����@�̵��9��!��;ɲ3O�},�U?��&�Ɗ�����f����B���e<=�4�������z��=��3�4�����`G��T��Q��N�ݣ4������]<Z��<��@H�[ɚ%��N։5�`��w[ͤp_�ȁ�Y�N���p�B�%�)��	��/�d�[�:Ƨ�+2=�� ���%��Γ&��8D�|%Q�y��H@3��#K˨��m^�$a�j����۷�e���j� �87a�?)!f$�* u������xc�����Z*�1�Sv�_�';OsF�N,l���S�Aff&�-�>צH�"p���e���	1����cZ�8iG��X  ?���$ѥ;Gݗ�Ks���xU���h}�n���E���$�Ђ:�z�v��~�������W�H�3��>��/8���&#���qw� 8��-_�Y/Fa�7�Td\��n����l�`��ͣ��������l.��� ߘ��Y|r_���.�4�K
F=_��X'��W�3�Q� �n"�܃%!>tQ�E�l9N���F�)�/��4���M'������x�����w��x��3G�ƀ����v����y+Z ���b��k�b<�Lt��(?�5yƗˇ����/(z&s��y �ԔӨ�@�uC��F�\�����\��%Y�$I;��?5�[K<���Q��a)}����~E���}\{��=uMp���^|����-�h#u���6���q�K�Tu�{#�dJ=?a#M�4�\�&�9����O�0�܇�۹�c��Ų��R	��.ץ|�6���AP%*>OL����b�sK
��ƹJ��v��ɽ��!Gre<�vC^�����Tb��h������\|�J��H%y����j$6�Y�v���4���'j�[��` 3u��4===��F���[�+#��Ej"3�Q$U��2`$��EB�U3�ѿf[J_��m�)���eaˆ�/��fX�=�HM�0k,W�L,@6�)¿0a��Ś��9a,�z���cf�ឣ�^I�',;@-������"�A���k+
�k�`3N��IAUY
�[�\,��Q��/)V4(�ߴ�fi۞�[���
�j�Z�w��{�^��~�� ���¹��k:�`�n��9|���o�y���Ԩ�G��|��0����K��O�D�����1�P�C���H�+�T>�jE
��UM��i*�5�S�l�3\�����b����'c��!�v9�Z�A�!� ;���'������/��Ҋ�1u&]Ⱦ��Hx&�ekE��S�͞?.
ױ�	�S�� �r��~�c��C��8p��:~��P��vlk��W�����|Þ���{i���>{~f0��u�s?-��B���ϼ7���5h��@u�[`U�D��Ba2(�}�
�-�\��9SD�3CS��%�w6�t�,O�P5��s���J�{7���ŗd�}�<�� ��g��Z�Ref3�Ni���R����U�.��ʣu�8d�XzGuW w!��|��ʔ|�D4��s��!�p�N��]�;�w�k�0	�cMw�_������͈ل�O����;�����3)�qj��zH(�w�p:��ڱ���~%�r���Nmc�Rt�bL0��}�^#݃��[h�:s�'?�ԟ<��0��/>��Z�3��A)��
x ���{���y9�D.�;�X��E7߃�~��m�"Yu�q%���w�?��2]�7z��|ȏY����0�J��9���:T����s���	%���u�%&�f��I7�qO]5n�3;F'��4ߤ�w"<�k~�]kjh��}��c��G�R�p_�:E��}�����-��-\��O�x$��zc6t��#��wgR��H�Xk�F��}�0SFhEڬ�˞Ho��~�$<�L��+A�Jc�i~z�3�e�1l+��yz��Y�d"��rZ�2�1�D�z�^w�V�K����_�t� 9��1���v>�g��CC�@j��� �p3��Φ97g�:C�;�X�&��R1H	�Jk�zr���+��@����G����R������ y.eV���֟|���?��}�g/�j�m��]?���d0Fal�c��e�P#���2�vy�����v�lj�"�D8��BN$��0���l:��x�𽷊����ja�\X�|��~5��A�%��C��A�W�p��I1I��%��-�sy(J9�r ���HpB�b�K��M�[��'�ո���dwL-�ֲe�ز�];u_�*h�!�)��M~�֐tġ���+0j�U��kE��q��.��c��#�_��twu���ƸI�;��	�j*
�Θ3d�ko�Z�IZ�h!�n�H.,�Mj_o
�T�����5H��
��w{�-pq�5��o8z���_Q� �����>�x*�A�l��$��i*@ق�r�1Y�;1w0Q�j!2C!um��e���R���Y/�fd�
�Wm.�h�h���V�H��� �O��a�������TG���@X���WF\s�WL hN�G})H#��W1Z;���j|��R����)��k�JY@�7��K��pb�|;g t�9�L3�/W��g����i�Ɍk�-�9��;"Q��6��M���?3d?[0�b�0��
���`����&<O<N�ӁQ�%AĹYw���V���y6G��z'���v�hf�$Cf���l����_�����I(���g���HOҗ��3����� �����=חH�bm/i�>=yTW��p��J=��;�?8W��V��c�wq*���m��[;�Ԓ�!�)�FWA����C8���\oL�v�r��s��u*F|�=�e�8�ɮ��5�IԏQ�7#_^x��B�P�HL�#�틘fÅ6AG�<}����l� �+�����QYj3�����>�v^ߩ�ły1m8�F��Pl>;;{���	巻& ���	���X��
y~���I9�B#���bS*5��:$�p��H"���F��������ݱ���B�.͋{@}����亦�Pz#$�B��H��'ǔ�֎�?��V�.��=����]�x�(�ȴp�h��5��Y
�p1�7O�[DXxs%����9XÐ䓢ƒ�M��ߐ��3̓ѐ��Q��l�ch�}�e*�\C(
)n��a�1QL�n�d�+�`c:!��<��n�L��9��ׯ�ӻ�����	�~���&��#J�&�o/z���A"�"��ul�'cWLmJp 3],��*}D:޳�[Ik����]j����{�.��F&�=���Mf�v��vx'��)�SV���J���F�.�sM��f��0M�p2�l���p��D��]��e�:3��(ٙf���Da:7��;iQ����ِ��(��P��=K�`Z�,Q�����/���፵j���П���7�l�l�}1���ۑZ����g(��w�t����p�H��>v	

��%�£h4k�맹�N��#��#Ғ�� ��9f�X_	��`�Rwi�U�9����)mo)s51����D�&e��e��̗���U�Z\La����mq~�,n�Z�{��6�n�ǹ�[���ϙ߸�ȝ��� �n]˽����SnO���> �o�]���]���]���]���]���]���]�_�|�6������$*	=؁qA�ڽ�ՃE����S��}�(����}�鍸 �5>]O<��^9�X׷�r�Ӵ"���S�CgB�>.?\饪w��N��3T�͒OoM�%��A]/x!V����EmE������n���o�o[Ł����ԼZDD�,��� !,��c��!��%ߌЃnTgt�\l접�bB��*!ʾ�jj��?�;ܘm�����=�.FvL�O�>=7c$5����Cʣ��&������4Fy�0���q�����za�3��ɰv�Ԡ
uji�~�W�ƴ���ٞ@�y������kI٩z����T��6r��_��G��<�/�D�+�Z~����]�]�OClC�go���?}O�.��L�~6h[��ݒ4÷��Eb��ٱ�'?���E�/�ut���5����c��u?ߔGƞړ�޽{��UR���
]?U�PK`:&.Hs�~Xj��9B����@�����3�����x�Y\��]�������~��av�ҋ����&�7:z�h��߼<U΋���y���x��b�޵�\X����KW����3qu��UT򚚚���������(�bm
���n�õ��C����277��pUEⰒң��K����+�z�߃JZ-Je˖,��[R��e�E�˾d�-WFH��k��%	I�-�l1!ː��s����<���^w�|��,��}�9�s��Ae���P	q�"�Sm'�Dp׋0Aѷ�d0��V������o��AwL�C�S��?ݽ�\�2rKȤTĭE�:����A����OOO�\���b���H>��l�o߿��GO[������0�KPRR�-�ū^�RB�Zf�R���u=	�7�m"''w&if�/k�� ǈCǴ����zk>~������gҳI��A_�p�ب�Ěw��.G�����߭<+�u�����/�^�#���>�%����=������0e�9vqЏ2m�=c�NZ�5�r8@�����P�
�ء-�d0�\�GOO�R������~mӊ.���[ξ�fX[ض��J\������f-�D���� ���x�b��EN��G�^�4u�������$����<UO;�'<�70J���X{��s��vN����uҹ�
ї[H�~�ܑ詟��e�%�`�}u5��{O֩Li���*�[{K6�q��4U�W�C����*�����W��OSjB,M�[�����6*A������ס_9��)V�R�s*��ކuuu�5�5&B1Ȩ�%���Mۋ�0�4��)�K��9t��ԔQߌS	�#�f"�oF�������9���"�Z��_�1�7�S��ÿG�r3���{z�0pȦߦ�˯�x����՟��Ԥd��1ͦ\�>�[l��ۅ._IҼ~��QLLڭ[�b��s�;��<���Os�;K ���W���'?%��mZ9:�����Ν3%C��}łvN�02;Kij��!:W�4�ɹ!!!LE%�㏻	��=-�G����34�a�`7u9;�Y1�Y���-J���C�FvtD�hK�zt����e�r��a�
�9}����EuJ�9%����af�/���)��ߍ�������?_=���6^Pݘ���'�^���]����n�O\+د��s�<���+�y��G>������s�P���TEԇ��#�`\�ͮe���׻�SVj6� �Sl�̞]�|�Z #2��o_#<%"�Ã���p],��m*/��o�'�c�dÙ�
GG��ч2��^镕��϶xj�@��(����KН�8��3��TxC�NݺS�RP�{�M܄�<:Č������{�><:�d����!'���zq���L�˶~*��  ���"�ɰ "}�'Ff���|FFƜ�1Ew���ulm3.����֏������c-�̳�ۄ��^�PZ�?�x@�?�xb��]�\�KE�K�_D'��Ss(O�'U�_����2�?�IO���x=�������	U|a���#�vU��~;���o��;���f�����Ь 
Q��ݯ4�T�M�1��k��S�~�C���n�W91�)]䁮�Y�۷����`VT�O��1�r�-6 }�Q���R��,��2��1ְi+�}^U*�H��C�/^����g�G��t�;RK�%jh.�u��ۊE���*���C��o��ej�����",Gp�O=����7*�xT���xt�!�z����͹2i~�F�S&<f||�_Pp�����M^���%W�Ʌ]]�>�	��D_G,@�2�n��[���jd�E���q�/�6EP��X��:��^�3��Z2$H�UoP[�q���; "�����g�͍�2��� D��_�;���}�SQy��f8t�&��m:R��c*�f-E���u��|]Tx�KCA����!' �jk����MP������ڈ�u�o��l����|������U��Tk�+���8;
�H��\��^�s��1�YL��/��~�J�@DWb��׍���ff�k�1���]��y��mtf&77�	,#�������ʢ/!���)efh=g������u[������2��.�<���h����ľ�)���r���N@-t��w�P�X�|�����9�n�\Zm43'�v�jiY�c�(8E��� �y��`�ݡu��Vp��Z�����"�W�nQ#�cߕ�u�@��NY9Z=M�pc��vt�%X��dP�B8`����-Kkv����;<��ia���o��r��1��@Wt��s���[G|�N!߳9�ξ�<ۙ�"\'-�'T!� xu �m�v��$�hyʔ�0Q4詈��n3?5ڽ�����7n�*�gj���y��ׅ�Nx��hu���k�sKE
�.g�XB�Ɡn|s9�U�g`+���.����a�� ���ƅ	��Ww�m}���'15tW`^��}�X�}(kk7;;:ҫ�QR�K���n\;�:�F���������/�սx썅frrrܓ'�ַ�&Z�Ey�j���4W�S�������þ����/D��.�Qd ����|ɣa�-r��v��Ma�r���@̽�7Z-�7��yV毙㓼��|1�'�Sҗ�-3�=��x�����\C��߷��G_6�V`����l�9/�b�?���swͺ$
V�mK:��@(� !!�g���J"�����<�"����2Z����ILX[z���`#�`���j�>|��@4Ǽ���e��3�K+����	ɚ�>��FI����"�6/��oss�h�Wq8�xˢt���<�VN��@`�u�������f�#bbx`��>�P%�F�[�0�zu���ΐ��C��$%xfT̖�X[[㺶p���S�@\V��ֱNDWG'���>Uf*��m�\��!��[=�#.P����]��kij�x�cܹ�chȹ9cž;�S�fU�2n�~�/��˪.ʹWn�`Ƃ޼��jm��=�oz��DRaz
^&1V=��rp=2��[�<�v!�t8̼��1��n{r�}h]Ry�4����E[`��f�^��萙�L�9���^�:��][�nr���<���ﯧgf�
=�^@�u����4[��d]�Ƃ�Ү"�����M�^y�cv|r��Q8/?�?�sK~aa�2@���坌v���i�[��p�}�.��N�XM�j3c\�z\w��a�`:::�:���������tM��m�gb?�>��*��@�So��{�n5Ё/+e�+Qw�>��·���ʁ�������-���K�~���9�)N+�-{j�l���I���U����*&FF���[޲������4��@�-'�t��Y�fyKƕ�jE/(H&��֛�������f�h�8% �!����D����<o;��Fƌ�\�X�;1.N��U�,���(B��`�-���2��I��y�ec��ⱸ���#Q���!�&�(a��vaqQ4������z�G�~�omj G;�\6�D�+P"�rM�mM�v� ��޽υ�U�;���W�;��O�)�K��)|������5��X�#.� ��XD0���ã �`PX�?u�ĕ{W���rTהn4�㺶���#����^y�>�챩�F F���^��~��!N|�k���!�p+��tu�ZFF��tu55-T�D3�>6󔳅$�L�\������?����(kgi����~��~)9b�(��B�K�����\U��������\��Fط�0�����ۨq]Ŏ��D�聦-�w���<���'GA�gܥ;{z�SS���7O_�YZg���*d�ˇqW�i���*\wx�(R�>�M��4˫^'��!�����L�2oq����Ϲ�ПF�ݣ�H\GGw�����"XYi�n�u-�ބL-p�*�Ou�o�	�!,&��g{0v��j���3��!Q
�C,ӓ��X҃\��H;7D0I�&�˭b���)HcY���tP��+d�Rs�<g��w8#���R _J2J��Չx\�6��]ۖ8 m�l�j:@|���]\ǻ�S�JJw@L	�跈�A��H�8<�{�T�c���G)�-3}���Kc���͸.AQ� �wݨ���m��}v��A�rsZ�s�46^����J��|���f�++�@���Գ���PQ��~�����������E#}����AVJJ}A� 8;t�`) �E.����qܔ����?4X�d�;1q�B�٨0�b��lw��mW�|@!���o1�G-+3���h���"���,!I/^p��;�	O��51��v��zZ5�3o:�b�@,j���ڧ�&X߯�xН�*&ff{ �����Owi���K�Ʒ�mx��L�\��%�)',��������`�龜��3SSm^Ջ���,�N��:^����[��u��a�������%٩q V�J�X�>�ڗ���� ��@L�xdxi��`KT����}}}��^k<Z�ʝl`棄n�,��8:�N��Sc�?�u�	��o��n>������������6��ي9y�#��)w��r��B��~���&+Q虁�F8�_�(��wW.��RПEc�F�2j�bT�砏P�W��M���,�]�X�cg�k��r�G�=��錴B�'Z�/���Y��i�`v~���#�'��`FJ\���|vv��Jȩ�f��t~�6��G���DX:�΅�-�v~:�( �Z�ā��N�T����3%s��J�f��3�
(�2h^C�qFt#kl���-��̜N5������z���1�S��rZMU�:t�*C!�ʓ�z��ǂ�HWt5𾢒���n�2�Dg�i�R#O��>�EJ���Ci�K�m���e��։�P�ah�ro��r������u�f\����>7�SAy�����??`�� E��[�$m �i80�A�|�����;ڝ�?�����%�]cc�s�N%�}}H���Q��KӐ<�^Y�!�9UL�m�\=����QVP�dm�"���C�G�764��>���}ud:���̬,=-�羰B�C�P2�~�����D���\SRV����;�Ae!~���Z_t���:�����*��}Ŏ:��S��}�}�x���<�����{�����$i�<������8v��K��A�ij����Т������A�f���q4L�ʉ��\�_�.�32b	�����bj�]��8�4��w�V� z�����b+�sl[��@��9:�yxY{P� +�D�W�e��j��`��� B�u;:V���&����a<Y&��v�O��h~�-DA�Ģ()�����eTV�?���d�%�ŏg|'bm�.���3}%Y/��D� J�u����Z46��|(ӐH�R�ulA1(��н� ^�N�gA3mϾP�g���r~ˆ҇���5gff2��+�^�{���а9R�t�@��gt���9dl��w������'C(q��<3'g&D�Ԗ1�$���A��
dٲ�����}�ƺ�r�g�No�<9��w�m�$�Nw��K� 4���{�ߥ���J%//{223c���wSy��S�fa���'<�ݿ!����َ5�|ǁrbȭ`��oߞ��3��(q05��[��X޽gOYx7�X�)fţ�q_��\��}%���g@� l��{�I�+5�5C@L����f����o7��BPfTT`�Z�LDCd�����:��a�9!fd�����@��_�t��lȀ��&�T��ۂqK�;��#\�������;u�������-���I�%mmZ��e��N���v�����������V:�}�LU��ւ�Ru��7��Ԡ����3�a�*%` p��;&)@��?���RRlM�CVEE_{���q�4���MHA�k��y��F�����v*�V��n��k�m�m�٫i���'�JO�2Tݫ��?�=J���e���wͣ�,�E�z!c�yx6��//�j\+���]*]���DHx�XU;�Vw���W����g�\5��S����5���D��K�uE �T n�q�a�D|t7�*����R�o�e>�0��TP3H�B �{�-䒌 y������4�y%%2^�)*19X,6
���F����tHH����]Y:�z���y=��Mx� )����e��v�h�7Mtp=�M�w�V�gpJڇ�'�*5H�n���9�Y1�.$�/ !B��R�J���4�j$���{�>'��뺹�>)̦���������<��Fju"��/p8���..�����H��[���7�AYlq�6JW�	��������>�V�j���z���V�
�I��v������q��||m�3}@E�M9�����L���bd��A���Y`���e?�Yii=jjjBO��:�2}{�<��n�������[��-�	�BLM��@�`��Y�2`�qq��Ӏ{ cs�?�`�����5��h�2�l�[�.{�O9���AAA\ǖM�km���3[6ɑ ��-,,��-,,0������c�~=B�.~�\l�r7��+�ˁ�PJ�R�`�6=ݎ��q��4�ǆ�(���Ye��}��Gd%+�w�v�!���?�}U!=ݏ�!J�-�wn��+)��WS%d��^
�ۑ|��=oԭ�t:�Z\𲷲zWby�.�8یG���m����������t@���,���(�g�Tf(O�<���rGo�� �Xp���)�����/�A�֕�����Wa"�}K�����#.=�E�%���?f-��R�u���>d�_jS.�,��{VnU_Ymhn��j8ߣ��(�l Ef?^�m�KK��/]����˶������ܹ����%K��	ʱɫ�繒��� � �!��h�U4���a),tc���2�R�������u� fɱmx1��� �+��@c(��ڟ�]�G<�K�A�l����V���(Kxߑ;�hJ��T(�ر/���}{���#�hJ���!��!�W���,�3�����J���oƺm\o��#!�ϻ%��V*��FB9��(f�Z���֕g^�\1�D�� �|�v3��C�=	,c�tX-ԁ��SP�j�
<�s�G7�:::7.��3�lw�a
?��u���t�I~�ϋ�@ׯ�	�p)Cw�\�bŷ
�:���i4\����S�L�����7�m�I~)���P��$AQپ��mhh����Hc�����wL?Ozݸ�
�#�A�2T��de=����]��[����T<�ܴ�]��[�>d�AK��'��z"-#uW���"e
?{��? ����x�"�͡U(A�T����������6�C[XE8�X�R2�TQ����ܺM,6�Ύi9�h�10�s��.�n���׮�|i���+#Sfz����EH㕡@�T�TR\�{2���_ܴ���]����{�ǧ��x�������SSZ�	���A�����Ɵ�b�S��߽zS^E����{���v�O�$>�&e�HC��F�� ��a�~C�gh&I� ���8X��_y�S�)*h-#�Ɛ�,���B�)~�B����_��H�BҞ�6����E
��
���A�gfj���oqc�S3 b�6��(�25��H� D+�@�Mjk����_�Ʒ�c"PQ�<g���44���732*{>�/�(d^�}��rJ:�>J=����ֶ]�0؇OX�����P�y�����Z���t߀�\TH�cnn�DK<�!'��r���7�S�1L��q���ݒ�-�Z;Tm�����=�o�7��E"䙱13��0����J�� ��������IOI�^<Q\M�K*~�;{������oz�����K� �_=O��m�(&�ދ���D1.� ���7��hq����4��!��Qd"�l���o���`�Rs)3�-v�G���}�_H;c����������j��\f^^k{9~d����^>^=�cu��9�B���vԘ;p7�ʲ`�X �܏Z���-��<��;���߇��9�20`�q��^��=�G�[Z[K�����sXԋ��h����P{9��d�xbX�(rDjj��)M�J�B+��IvW/�\�����Ȟ���>`�M����_	�НW3�j�YRҽ��Ъ��Uo��,., ��_e���v�
��k{�ɹZ����
C(v��a����k&^����_�ӿ�ʝ�y�f��<�r�p3�p��9NDs�(m�L��x�R��Q5k�v��c��
�;��*d�2Й��]\~ĵ�k�
���QX���߫���3X�O}���UC6m6JW�9U-ĂO���랬���۷o≈Q��L��������>�����?�>����,_���̬�y�w�%��Fm�;��s�~M���,�������{�8ǥ>��pif�f%�)��Z�������@[��L�v��a�55C1�e,��M�5;�H�\���!����=[��<��HƂ2w�u����� S����Vﰐڹ�z�۷�	��oa�8��S�U\)�n��=��� � ƫ��=�Ɩ���%(~����e�����ZW4}������{Z��g��[�ܚҟ�݂�j�iz��J�=ܿ_����湴�4@��9M����Z`��8�=�
� �m+ﯻ��4���(�DN�NBZ$X�v�:e��P9}�5-M����?����nnVZC��j?	�������rPx�kB#Obae.�?�ZGf)7�~����j��zwJ�i���F���V�Y ��̯v7�� .}�"����Y�N.ڢj��YR驧�!��F���x�<�<�⒒Y��]���g�[�����Ӕ�4��	�����t͵����	���]��UX�f4CV-�\��UT\l��-�[r���{YTbm��;�H��{�Bo}}=�y�W�$������Rn�V���@���R	����v�fr�������y��싅|D@�����/B��� `]	�u���
��C��.
�f��WY�P�޿��L�=�A��,�G�y���&(�����"9��b�/\�g�Π=w���'��T�o���l�q8$	M:>^��>W�Q��(��'j�Ѳ���s�t��5UM��y��@�W�,R.��!�?wtt�%�;9!�/H���/��F�����Z��Z���YY��>>>����V*[UC��-�A
�O��4���VbA�����������<����B�=�=�����E�h����ۜ�֦EOOo4�f�!�/�k^�)Q�sl�N�P��)���$�D
ư���*�C#`�`�B��B/~Hַj0ky���ʉc��pG�I'<[��u��R�[G+E�4�[J����M4CR$���,wbb"K���Ȉe�ͩ��U�к$P��;'àҗO>�C��.��fn�
M�����������:��@�`!��t����5Z��$�N�%���׻��D
��͖)�'�.�r�+C�Y�,ʟ��j�v}�[5�?����O{|�����pׇ��A��"��t��_a4��՘��3b�b��3RR�ɀ ���p�v�w��%9H�̝A�M�W�U��ds���G��l�΂�F�%���_/^'*ބ����Ń�v����1+Q�S�9L^�����')���N��w}n~��8I\L��ǡQA\H��
Ph�����^�B򉪹� #���8�,��z�bT<��A�o�en���7���LVq���UB�p��0�,�30�k����A3��鞨��� {�ݥ}��j���-䏐v�t�U��B�a`.���
�TT�1wi���r�%555��r�x \�.9t���� j�m4Ui@��6lQ][�Y�!�s�FV^u&��ҧ͆��E�S<C҅d�f{�,עq�Od�S�gTl�W�?��j����K�0���
�L�t��-�P0�8���stLX	����g������"d�����:��T�5�u� ����a��i֢��o����������NR�1�/��da��~5��˙:ۜ�O�ӈ�_��n݂J��K�î'2G���E���K��"��h8�V�	5�H$���d��}�"V�*."b���? �"53����������G�S؅<�I�=X�in��/,�Z1P�0m�Vڰ[�O����9|������Q��r������`�I�܊���� :*?�K���f��sC�k�+�QW�ڒ�]�����>�гM�7����:����Yۏny�0Y�V\,�%ťfpR�)����� ��O�@�ܦ��3��������
R$��������b�O+T��Ҷ�cA�Ν�]jSv���dC�RTG�Z�$���̂�O~`<���i�b"�H	��Y�����������!� � �ߋ��Qd}����0��i``��+@ϠL׉8LQ@'|��Y,��ݽ��j��u�LZ���% ����ɪ!<�*�Ӎ�%����Gp8�_[��_�.��R�G0	�G�à��H�t�}���&5������S-��оڦ���ؗ���grhӶ#�j��>�����#.h^=��������]��#�����m�"��3��kg�>�����0\���HS������OVy��SaIԆ���9���YT���{���͉qځb<%Ƭ=C'�!����#5�	�����?Y4��Lbecs$Ty͙���7w����'��>��_�<����t�^yE��)�a��������'?�2�]���B�Ho�<؂�,�B��x��,�\�]�����)�J�F�*�6U��1ƕ;����WT��c����r�R��n��Ο� (Q�w�PЦH))��*䋎������s�r+O�/. _�:_�j�v����K�|�W�1��>b�
�qb�$Fw.^± gel�e����/[�\��F���z.&��顗K��;��XE�_����붶��ǡ�j����O�4M-���g�+s�g��#1+3�t�Y�t�/M�T��e��n�����@�:V��ˤ��oYbՏ�IGY�
G����6�'�����(E8(>��z/
&�, �:.>ޚ%D�Jߑ.ߴ�#u
�I/�!v��=�$�/�����"��Q��,�TU?��vX]]-&|���0��,<@�#��H�Ñ����_�'G���27Ot��2<���u�O~���"KrJZ'G_�m>[\Jʖ,y���ޖ�����䱃��1��ƴ��9����?.���c�U3��i��bT�̜��E3x�vF8��arವ܉%R~ܥ��|s���6�!G��߅6�
@�j�\*vo^w�v)�&	_�:$vP��ħ��N���Ҟ�Avvvߩ���?��-�	Pۀ2:� ԉ\3M|�$��NC I���/��sE(���0�_���k�!yD�I!���=�f�����=T�#����o��+*��Dk[h�����ݧ4��ۡ�f[��bç��P�-v������F�	v��k-�eN}�<v����!z����w}u�qF�cSS�QwS���D�smm��V��k#�����-��w#A[�������0N��2PT�T�/���7���k3@���&$��1AY�ĴŦf$�������C<N~�듙���iV�x�����;U�f�T�D$�U�/_���s�[Ip�Փ�*��zu���.by�4B�^2�}����9��<��@9��ě�r䦧�ǈ�6�I���T�OyN�8�KH����8���`��3j:�
��S��r #�F>=xo�]��"jn����ts{MW���%����Gmx =��f(��o������9D���4m>��{!�k��>y�)ƚ�Q��q�W��X�����?���ӝ���g^9HKy}�j�?���\�avW���\�cb�z�h�9�\(�2���ə;���T� �����E@�^�~?��+__I�p$�h�F��y�g��,G8�]p��!�L��k�E��ꑮ7}�97(��j���ŗX�e�c������dVR�e���ҝ:K����yo����׹}r�������%���E1��X�ll��~~4~&8�XzMM`������٩�@)op��
tIJC� �m�l%ZYIu��۷���1v��}���O,=0_{۵eO<.�.t/�+��+ ���A�&�u��D��w���A\�M �Q���7WeC�����Aν/��a@9p�u�^zz�����Mn�ޯz�\'���n�{��.?�i���U���ZP%�rFL�^,�T_W�ef&����X�����L�����}	�}d1		��z�8H��AԶ�K��8K�	i�*�g�p�6_��x?��*lT�s��9��..5$$�af�����K@Zʫ5��,������`
�S+F=�qXY�k��u��������o�m)R)�����7{��U�S�qK�]�;M�6/�j5���ps
op����
{���I������ߜ?y�����ey芠���
��mZ{���x70ٳ���y��l�n���k,!���s�va ���?ѫ8��fh0N+���I (�{�p�=�D��`��H` (̽ T ���zތ�S��쩙_K�=`W�f�}��c7��8������?�����>�4�/^�lb�`ge-�3�{��'%@)��T.�f dy--�$޼�ǉ�bvV�Fc>ie��w2����h~�p�>?�пk]s2`�̬��U+#u��Z-����Zv2�Q�	S[�|8�j�0Gt��WyWGG!o챩e�U�lu��.������'�Ur�-v�#['�ޤ$%�Y�N�]��c���۬3�h�.&�W��_m�j����(u�/�7#S�`(�н��U{�:�Q����i�P&���c�M�ITMh��ɢ�,Zd�ZIQ�Y����ՏN;C��Ҙ�ܨ��k����f��KK��װ���=�9in��0��}O��9���.��BOf	9m����g�L�X��Q��~W���X
X�b��)��RCP
��T/k�^y��P�=����}Pk�6�R,iؑ���>���,p}Ui���, ��G�-�0��Ra�˗/C�q�������iX�RWq�G�}&��T�V��aj�sWɋ����~����;���5��T�$��##�U�ي�Y�'!��d�}Tk��7���g��mȤ���ڮ_`������]�����)������#w5{��3��}o�/~����{��{,`w[d�R�����q�ǒ���H��6�w��%/��犖[N�3����>@���O9�gC؜x�g(x���&�MO�n��PJ؝q�{<xp���$ǡ�A�%�*v�~�Y���ʟ�%�_�0-���36��u�m�7����P�������Hh��h<�_^%��=�6�?=�:8���k�s�hXJJ�7�Q#�׿̲��^���z�Md��Kn�&�������U�������g>��̣����9��e�LLL
���z͚���t���<2�䵸���n�7B�����S�7W:����[/�p�8��Bǆ��oWcH���|��U��}3������νa�9����1��C���Չ&���ש%4�����V�Z���%�����4�M|���\Rc�d��>55�Қ����ݭbĖ�;c�Ɂ|s~�U����Z"�٤�X�o)��ײ�gj(}5��9_�|9��mb��WxfJ6�nk{�6ݎ�-�����;�R��7�afy���o] �Β�~�{4�O>Q�#3�#xz�]�ЋU��n2k�2^'ńu�nߒ��Yo\NQu�[:[Nx1�>�챾��8���)��m{t�� �����L����-)�t���<"�{q�BD��a�s`�N��e�z�w�S>{*b�0�IQ�y��3����슌eԙ��|ك$��y�{Jȭ�-,��s~w]��Q���,6n�؛��Y�jU3�[�M~�.ذ�tBK+�^���iwq��oqxUD�q����^.jwz��u����D}�}3(HM��x?%Ȕ����$�0Qf�T�6�{N�:5oH4H�)��{�.<8Lt`g*�i�,1�3�z�J��Wџ������G������.��=��OL2�<M+�ߘWP����d�?��!gZ�w_�~��t��T�-+d�����]9{�) ]�R\�0�.=?�X��E�j��Yma�ۑ��	����j|"�����F�_e���Lkb�8���1� �x�R����ڸ���-�T6���+�^�u����!�ܹ�޵�����v!%��#�K�o��/�o�&�� GRA�~ҿ��[;�[�����
�
�L0���d~��Uua����`S{{�6�2�-����6��l	��;`�f`J9d��}C�;J��&�F�`b�@���K"�5�v�p��%y��]��-�XU__�e�v����1��ͫ�-o�;��6�.f�� 0a�#O�t��u�U��X[���h�.�#OD5x���#i���Tt=l�+^���5k��G��R�a����h���<첷ظ�,�C,��>�A���0�����v�v�S����Rm������UKˤ�"N��knRo�*���l�K�y�(����s��f�x���4�z.A�
��`�2�G��Eq��o�vuu]6�Lw*a#�%��k�w���E������gu<f�Aa��-AMCÙS��\;^�Sp�z�8W5h���36�M����5\� �%��6gT�D[���Feaᘻ��^�`��yӏo�Ὓ�v>���{��8g�7SO����@�V,���%�W~x�^FFF{������cfڔ9�@p��������UEE±g�D�.������Ӻk��[�f@\;{���p9��8潘m������+��H���A$`���lvt��/�ޏ޸9)3������q��Ys�zZ1�t8��#���3�~}��DeIߒSr7y�Iug�����eS7�7��w���B��D�k�������"5p�ܚ{!��W�Wj8mZ�	z�I:���'��5Rr)Us�ί-6�il
�w�t�e[ll�ݻ����o,4�I�r�3�G�|Ōs�31U1��� ����9]ōM�3#3��/x��.'˳�]�>��]�)�iF9�n���[�x|`W8f�rI_����{��9-#��&�h.q�/[���B+������)�R�����Cr��OE��k�'�]_�����״���4��>Vn�Ft�m��V�E�7~������6sw�&���H:��{� ��}��ț���H*���˗��k�(�6j@��n���y���Q����*���uE�%�z��3�f�?����־���3T��ᗽ$^b�) _s莗�D�l��y�t-��B#�
�ے���ծ���t���y� �ے���'ܷy擺ES,�����rF��Kۅ�!�m���9gzI��Clll�_Q<�Wg�j���ӛ�.�<0P=���u�]��r���a���Sp��1]���Z�Кڔ���Z��۴�߶����Zt�)G?����W�����"�Y�������z�
cQ3��%�)j$�}�בz�5��5� �H��(�N(�����������Bss3x֩$��V*i���U��<CԦ����������xR��i�˱g����홗ް{� ��$Mg��ɔ���υpǜ�z�z������Z�`��|���L���!š��!���u(޹L�4F���c�.ԗ�ڈ}�ė ���W�d�����([�_�zs�_�)8l.p���WQZʲ����nhb�~����������{6����� ��n������h�c?SP#m3��\�K>��� S���S�[Z�;:t�y���t4����D ^�oi
ۧ���<�f<���i�[g�6c�J՜��&9:���S�_ꢍK�&�[���ϊ�>�Ȯ�_S��4�Rc5 4�Ibb�^H������}3�2P'T������	~�A�j�Ο\�s�h!D�R=#e�S<�?�7�OU�aF�R�54��2&�7l�׼ߡӟxs��a3��#� ��^XH��!�2����qo_ѥ�Q�sJ#0����������C��?��S�5�j�G�$�?��y���H;�0�@U5�Ø�Q�D1"��V��	i��P	��5���Bϡ���B�5k�7�;2N�����֋�S�@��R��{�>�8_�����Σ?��>D/����79�^�&��x��Q��ov����ѱ��K]f0����;z���ޑH���<�J@��~
#c�VM�.$����jl����6�rU���NÃ:U�Y�n�%�[>}��U�b�T�N������,��!�5���%�������]���v�'���<�^UXK���j5��� �ba}v�:%n�@�z|��'Q�X"Ba�����`jj�k׸��
��@Cw�Z�D��,�/�7d����(���/�����V>�������T�޷"�� g�^����9������3��7!�����9
��6����5���gm�@�=�_��_�L%R��4v�#ú��F�v� �ɚ�Hm�s6�A�-�q��|������1G#Χ�/�����fo@���Qs�
�V�E��`N�C�4.Ҵ�Rr������l�R�Yl./,�5x�}l��Q�	�&䣚δ�F��X���T���É��A��U+ğ��?C�6�0Q�Y"S��W'#sc�c�"����w�ȸQ�%ǻ�c*��ǈ������"������Γ�7���#���"�~�x>�[gv��o�ҍ{f!��7d���!/$k��Kg �k�4⨮炔�z�Ib�"He�?�;5�(
�\�b@{\|۾�0����VN��mtp�p�+�0f�X�F�B$Kxå�#�R���54 7.�����(i����R�a��v7q���N�7�3�	'��ܿ�3���mvd:����F���bu��km)�ڜ�/�"I����:�JUA��<"�n����EE����Kg>~��Ms�H��m_�IS�R�N�����[Zb�Z���kn%���)b�f���-���w����^���h��J�³j[
�e�vG$ԏKgd7�/u�� i��/6:�w=+r�Ntέ$����-��VƈF�P �����#�s�攳:/Ǎt�q�F�Zy4� m�{����{�X�B����U�G9!�R�8��A����Lx�FoT.������J����B`v�~SF�$�2�0�
�����>�N�iص'淹�;�?�=<�$��/%�8�^�5���p�l�!��N��"i�)"��[(�R�F����1<0�p�I�#�!F�D�s��j[q�U��l@��U�S���e}���zT=��x��R�W&
i��l��d�c!��l��H��ٽ7�
�����n|�QPa���m^A�M��~s,�K�>d�E��G.�QُC�&����h��Q�.{ǎ�����z�x~�#xx�EGY����� �iϊ�����\\@#"�͖�>8ȸ�������<�����}1�j�5��C��،��`�X��v��Qڲ�J`X!�����{����T*R�m�I*7�iT����鷟>����'7���ݒٷ��Ș�e֣1l�&�6[�;u#�!�s��n��)�灆EGG�����~���Kx�o��6N��ߒ��mBڿ�g�M��T�_:>>��3V�Y�i�*4kԱ_b\�r
����m?T����;��L�@j��!26]�2�E���O�Q�B�8b<��vl�J�|A�u�՗{�X�u���:�rG�{ն��*��c�&�H���ze\uh�q����/������06b�1}����<�3��8S�p[�mx00���D� 0���E��;���\��bbt�7�KSs�Xl�ۥ��?\���� MM��-����&9���.�m�
�i��/���҃+����Prl������NE�ݳ�]~W�i���`�fGN���]*�%�Ner1���J�xK�X/�{���t��q�g���g�6�VoYuvK6I�߿q!��ͦrR��?�����'rKF��!�2F����5N��s���<Z�N^��/�<2�G�.X���P���˙��Vǵ�K��Ϗ�Ќ븄�`Ѡ,i%���f΁� ��,6��R��W&�Ŕ�E�����&'�-*^��*U.�/���G�H��:z:c�����v�F��r��R�M�v�N�����w����Db�� :��su R�ơ�'�K��E��Iu����,�~�P&��-�X�o�<�&h��&�;]+���u�H��<��e|�8Ƴ���$N* �s���j9�~����M��y�{ґ�_�����_.Y�O��O��1�ׁ�M����?�m�y��t<�)tڍ l?�X6�P6۽i��e�#�o�)3!�W��a��V�M�D��)Rq��ڟj\6-�?�V��L}��dϤo(rt.3�������:���ЯM;��p�������9����`Wd��at�X����;&4�-�Lj*;�h�}�;����O�_�6�h|�b��W���`�����Դ4eoS�!jb�"�ɟfs>Up����[�SV��@n���2�8���(�^�o�3g�@a��t��u4D^�Y?�O	Ϗ� ��RzD�~n�f)��W&��ƪ����Ǻ{�Z�DCQY�����GE$#��]���<���d����P��d'�{�����>���}^�筗�=��u��{�s�<س&s�z@�q�`AO�/�:����#����ƾ1l��une璻c��+jv��ݹv��{�ǖ:�I�Tc�"���{��.�k�*G*G*6Fn̸���(f��G����4�1@��I?�kT����uZ	|-0'��9�m|�a��ᢦ�|�#r�#�"C-�D��3�0Y4��`��J����\�g�z<\uw���%����M���W��ܙެ&�p����9�ğ1^+/2��b�]�����&�br���m t>�C /n��a��t����釂��W�sH1��mee�����k������"k�b��&��BL)I�'��k��b��Yhц�o'�b"����\������qhB�J��a@�XBn�j�T�J񄔮u�����/$�޺���(����"�pL�/�Vi�$"obգL&������70�c9o?E�t<��D��{y�-�_2B�+A��4*	�M5!U��U�����jf���/Rc�A1Ld�"X"|��#���~5�c��u"=!�O(����]���}��\T�
��N$q^&��E�%�
#���\̨2��C�1u�NJ�{�n�d�.��^�@����}%�g�^��~&� !�;V�bG�0LѻW�C�KHSj������~ʯ,orA)��0��þ�$���	�B;��N�G�~'��d�aL{�Hq�ڹ,���P�+�j�j.��R���?�;.&���RІ���۷yLg��U(5�*n������3��':��
a�ݸt�3�Ԟd�&�#�b�E>���e����v�B!`�%(�r/���r�3;�nr���c��$!�:p?ӗF~�=>>���U�)�`��I��~������w-����}9pᗡ��:��EMo���'3*N�=A����� ��"�s��&��r��h�'$�Ø1�V�	�ʄJP��ޚ���'(�+o�1P���pc㕦*?�m���X}[����| v�O��&�Ҿ^���^�Y�t\nb-xlw�p�����􍳩=�ō�V������	J��Q����U�<H���,*�`�2���}�>�&<�:/8�Q`��s܂�z%o�N��R�b��ЫD���7�a<���g���#���bf�����|:�����YEL.��(��~��,��fΓ=�.�b���Ƌ�����)	n��M�(�HŠ�ld?5�bl}cl�!שR$���}�Н�^��Nn�[+!��LxZ}_�~�U��U�]'Q�ƣ'�]QϢuP||S����p�)�)(y��(x_�- 3�n9�y;b�s��0������G��*䑆�4��\��y��\�_�xlv߉p̣�bc���ӧ+���y̤#��(���3	�oҫV7�׸�[ösnQ�b���֭�YY�LŠ�1�KX�8~���,����Ezkn���_Z��O�/��3�(���z\C;��ܱ0�sI�#E�	��V�wh�B9��?&��tP0�?�	yL��ɉ&6�Z3�lrV�����W��e$�>�*�sg?������پ脱�#G6��u��e${IV�֐�3��i|��Ȫ�n���;%Lv�h\�=2���{�i~�$����=��T�[q=�J9JW��:,r)�˹���:�&EF	vs���Osw�\�mK~�d�On0T)�<�%���0<6O���c�� f*I���mL{+&������S�LcI?������	jq�nQ�%��#�l���]�d����ܘ�UX�u�}�����;
�O�n�QN[����?7U1�T��D0ڨUp0�Q�P`�S�ۛo2�{,МH;����ų���I�6�Ԅ�X���]k�����I�	$x�|%}�ki�d� &{/Su'P�ѯ�+_-˶�B�����r)ʁ�$9w*��c򟝜h���J��)��-����ZL.7�j��5.6���zJƝ��|��9)��	�D�O�XV��vb����'�YZ�Qn�A3��GOL���^J	?�m��y���ى%�k����B����Ŷ�'�ʛL[�nَ%�Yc\���k�$�N�C��En�oR��'���6���4��F��xWP
���x*�RMY�5Q�w))!ۦ�|��V���*�cOp$�[{go�N@�M{�O�؎�ib��W�Dj9�wG�1b=/qs�;�u(���\�~����GOH�8�t�?��QI�- k}��D��Tl�$�kMM)��W���7�`ҟak�ZR��[	��qf�����4`������X�6����t��~������H����f����j%н�=ֽ�l���}�8Ĳ���O��!���m-���*�����(Xz}L���!��ర�RK0���l�R��_ܪ�Qq�LPW�}n6r*o�+���g`����>�m�`�iI;V��|�>��.��S��66�O����+�^���]��e������p�-�m�	������lł���0���(����$� TE<ҜM�S��c��n��x���%.$��ؕ}l�È#��mD�ƆômO❰
���hZ���jٳ�9&}WD��B����{m�����HF�?l_�_p�'��ݓ��x�����{|d�֋��Qу��n������t?V�Qa� __�@;K�q��[�K8���΢��ע�)���A�j�� ڮ���z;!8*�9�͔��	�t�z��S[>l�ā��tO&��:�j�F�OW����N��Z�u�E�싷
{�Q��� V5���m7Wc��<�n�Q�o$�����������ژ�нIu1*.ȋ0 ���b�S�����B����Ln��<̟�s�C¸�lCG�I�ku�洴����b �p�&����]� �R��H�:o��:�mM��?G���P�:C[6`������\�V0�)��BC]]����W0�`2��p%��b6�L%��
U7尛k�G��X#�݇n5�WP�]�^��Oe��hW1�TQ������ŋ�*���ϻ6p����Og�h�]�jZО�(��{��^��nQ{$�<}�RKӜ��8��-~�Hs%@�" �؀ln~��_�i�NUUn��O#蔖�q�E���\Ksc����������R;��1�\��zaL��yN�\��T:�}�^F���Ke0L��qs}8�xgC�R���x+�Q�>�޼M>X��^���ܖ��Ϲ��bA%�mP�	���R�����kZ��>��r�EtB�%�cS��łI�k隉��}u������s������4.J��!5zj�mjҚ8FXoʯ�?_8{���BI�rd�}�e�눛��֒���5�,� ��~7ġ�p���'B#E�ï�H
%�N)7{sd�t�!~҄�mNcT�d�ׇ���r�⪪�ህ��0���N�������'�m��S���檻0Ҡ� �1�_e��@	���6�~@]�'���`�/�����[v�~OJN6��n���m��������U��Q����K�t�ä��g՞��,��>ϡ�[�ՙ�+�)��u��Zƛ�!�>���

����0�#rl�O'�%6=��k-��ln1D��wߏ�����^�Ȥ�n6GV�0.D���k�g��d�f%�kn6����|�A����;x~��BT����+��f���Y��z�x��k�G�̎�w�n+��ɰ��-Mr�ΐ^�u��VcDA�����/Z�2�A�Ң�_�SGL{엚rz�f�����5ʽ��lOz�^�R������묯����w��yf���;�.�} I>���۳����-,,��Dh�/4�o�#t�7|t�H<�j��O	[��fZ�..��btX�j�d��9G�i�����ӿ=�j�[���)�������W���6�ʷ7H<3RSSWF g[[[%^�w�B(u�H�et3a
����ʛo�x-�`�ky�i��E,��xE�UsyqR��X����.��t��ǭ�x-�nt�fK *6�j� ��CFgg�>q�����_��*���'1��{<���κS��8.��RZx)H� m
��Uf��^��H\�z�|�n^RW5���Cp��A�����,�1^rn�����o=�v\���<��Oe����dCL��U�|��N���c��D�BA�����Y�[��A�V�Bڷ����������_�Hf�ɜ��M�b�BHn��oq������9��`Ŝ���QF��y2��3=�~�3��z�,��$�s��w���I]�l��22<,_�X�˥ߨ�Ǩp�z2���VKCg�����.¡|��s���c��y�I,�8:F����u�(iX���2�2=���CH3�M� k
߈��kj��EU9R`��='y�����P��e���Q������S��C"�÷pm��"��)��^�E��XÈL����xY{&�z(��/�@�r�ѢH���C׽GQ燙���yi瀋�֬Aq��9��e���<�}@�i}�>�[�ī��� ������de�MjK3�N ���P�7��P���`��U��x���N�_�UD��jj����������Ϝ/��	7j�G^���.�2,b�2�d�kPlJolL���mL�����ws>v
b0gz~I#K@�ҋ-j���nQ/<=�[f]��t��)e#tF��r�|9�1i7_�Y\�=0�aDm�p�Ս��M�NT�k�E+��-�x���t�{�/}���������B��':�,i�LqQ��G�H���h�2��� �;H�8L�J��
8���{Lb�������}�\ٝݍ-'~r���z��◚�X/��1o���F�ψ{}^�磍�����!�I����cű
&��?=A-�7��X��x!����)���Y�ېfA���D푙?i�;����;!��Jm�
9�jҊv{�lA��bjtp߂�xC9��kW�lG���K}�d�H��Ԃ� �9��ѣ���	�܇e�,�t����F'K-��22�ҟ]W����>��0ʕ�)�M���B_>�B���lÈ��������%���e�a����N�.��:���𝞼�W�|�[��xRfY�e��_�b �s�z���|�D�gk�	���Ap��]���Bu�����|חEC`K�Ս͌Z�����;�jq�hq�z$�*�4fZ�G�2�2ii�Ŋ����#/�\&͝58/^<���|y/_�W���m8�eG8u������,��kY�2:�(My���4��v�$͸{�������-`�T�u�/�\юl� �}@�az	��������xr.+�ȡo[2U����}R���A��!D&�!z^�Oܛʓ�ʊ���q�̐Ʃ���'����7�wVc�5�y\�m|��V�Q�i e��/Pj��x������t���C7ϡ%�O�;����Q��!�kb��a��+���mo�F�7\~JF� �U�=I�_���/�&���A�����`��?\6޼O�o���u�ten�Ҏ �+����]��`���.Z|�/b]{���э�]�K�~��i�_��o��51��*��>�6�O��q&��L��>T �a����HP�sB�������]v�s�ϟÚS�'-�;�'U�:F�I*�����~������z�B\����J�ka[����!�[��D-�Ȅ }�l����{r\�7[u���Ð�!�q)Nx�|*'9Q�8n#���%$�_k�#�5�~�"(FE�\n:�(}s�s�!3t�1^뽘�)J�ii��Z��9Q��*FX(:��,��x��2�	22�򊯺\f��_Q��0Y�P�2|���-<��R6�S 2b��֊�|U��V�2��2��%�*p�Ĳ�afǢ��� ���CCC���5��Q~�)%�u��tL^��<���x�`6 %�k+�-�,-͕�jLx�x<%O{�w?��G�$��7�����T�R�ٛ�t�Q5�,S�uKV��i��bJ��Q�6E ����� ��m���B'Pn��)��3H���@@�>|��׶Y�.���^����گ�{MkX�=�{�w,ɛ��	�ex|�zy6�DA3٧m4�R0��F���FohJ�Jjƶ���ӟ!��������ߗ|����0��->+hH����)��8�k�KY+��0J�d��3>���O�t%��j?C�"�7m?}�򌁟_�\�րә7�Vj��������T�k��>x~7���Nx��0R��.���Ӊ��ۅJ��/} wtToK<`?�a���Ą״�m:����yMW�Ź� ���������9#~����ڴ7R��c)�����\�垐5�Q���Y��LNJ��ح$;�/�>Ik�� c	���F2��������C��l�lٹ��~-�G�Vx�Ix{M�^��s\�_��r�U���66|�Ϋ������}�:����dLC�igZn	)�N�2�s�������)��4��e0�d���6;�k�_����0����!��k�F���1��k���H�����R�N��f�


�����K�[K����
�s��˟�
`��<��m
�a^�j�PҠ3��~�t��ŋ�*��� h�Z�����Ͳ�z�AB�CP�� �=�т%+S����-3xN���l~�X6\ ���x�Y���6�I0�La�7��Db�;�k�W�zVYlw*����33�رU��H0t)-��s��|���2�Tx����詐� ���7�r��Ӿ��Y�1���~�eo˰���!���|�d-�څ4Y蝑��/�JÉ��\VV��xS�m���4�D�~�Dm��>��n�#3_8k�C�."X ��A��erq�ˬ�e�׉$�KN���۸o�1UY:[���5��~M��;O�������M�ƻ���=j7�

��{0�o�~!�-,I��"G*ʇ�/_��:�`"�kA��CJ�!d��?�15�i��@yTw~NJJ╫:-C7���~Bk&�Ğ����4�g�(�d�OOg��ED��V���4�Ʌ�)_�`� Θ�dm�m���GǙW���T�����2�MH�H������9����7G�7p�%���B������ƛH�0�eZ����*>���[nl>'�`�=0��39"����StE�Ϭۢ�SC��&�V�;��+:K��^��sb���mug���,-HK�k_T6�jA^n.{o�R~ ���khی}n�B�˴���,�"}�>�f ������>/��N0���R�cM�����c��n���qcY�яQ�G������4����]|�>i5�^�;Ӏ�z��q8���&�:�i<1� �㼸�?ߵIƋ�Ĕ�g	�)^8n�l���^-�Y��Y��#O7�I3��{أ��ivc}�x�b�<�5H���e�2d��+3�>�2�i<�@]��Xx*�_��ml�	9��m�-�$9�� _�׽5�����i��[L�MM�7�
�,��'�8��򉗻�J`qkE(4����d�Ӄ���v�w��S�=�6c�/��5�m��b��2;<�Fj�J|0]v��V�~�w���Z4�6d�T:�E.^ϼ��]F-����3ގB�u�q��V���#��駪q�HI+~�~�R���а�k�~p�~����qO�!ćЇ/�=��&.��̓9Ξu���#Z XS�аF����Z2z�9T��[[_�T�۽ F�2����3�OyR���ػ�zYd[o�9@����%o���r��z��oj�:?
�O��3���A�k����y��K��^c��q�3ޔfff���u&�����ze���/��8����F�0�wIIb)-k[m�s��S��s�]��\x=��?y�!�̵���D��2����?{M~��΁Q��2�<�ldhh���|�P:�aK�kF�Ǔ"4>���)�;��Jp��kM\��B�U8n�:|)эibjs��dz8��jG�qAw�M-Z���a|t��6�s���i��|�������2{b�Y>ټ�n����fJs�l<es,%�~�)���q���=܆_ѝW�)��;���x�������
��{�����ɺ�󩏭Oݣ��+;�՞�ͥ�ر[��;D�ƫ��o3G(�	�T�AAA&FƬь��KBڻJ�PÑĴ��QF둲��tQ���K%���T#q5w�Y�f��L���`֜���$հ��&�����k)�S�˵w�5��)���D����Z��U'���4��y�����19%���$�<☼�˚yzo&�yϐ���o���P�~�}��r|�����"�6P�]�*#{%�ޢ�Y��)=���#.�������=+^�l�2��Y����U�9J�Ϙu�A(�h`��:�1� Ռ�u��X>|�6�cF��_}�%w�����,h�� �g��oSS9������%��!ܑ!�r��KI^M7��������)�i�H�5��Y7:nv<~(ZL���¾}����[Zp7��D_�=nue�9���ɀ4>��c:p>W#k�Zm�,(5��3��.ԙ}fE���P�[���ʁu�^:ʒtGv
#R2�����6<6w�l��@��;l���Dl�L�eF��G3U�HO�8��Z	�Y�}���ų�	��8=���K[ߠ�k2�&�s�jVϵ���m���E��˗�����u�R��N��C]'�,��CQU��%S	��a;�� �W`:^��L:ka��+��s�!!-�h~��Ӛ�'|�L�5��l48l�?�Q�U��j��yuę�&�>�Ȣ:lN�YV!R����7~u������n#���{��xg�����Օ$Ag�|����Rfo$��AKr��7�qR�lmm����@=��-�`m���?��#Og?q-���d2ߨԖ�p{bu<͈yyd��������mJ�������׺lzi<@I����B��SS���BK�K���Di}9���VH�������	�W��؃�Q��`�%sai�����=xܳ+v�T�
�L��b��ل簐��E���|���,��X���@��j�N%�4����t���sթ�;�'�n汯UԨP)1���h-��}<���{]N���qn������2����K���~-�����f���egV�W��$Y=Җ�������\��� �(�����Dt�ي�=����Ys�!�	�����,��Ũ S,Nu�6�h�>�B���)-y|���{e�FG_��JF���G'i�Ěy��ԌU�����k��3Yu_�J{�;C�&�t��C�';pPF��B������h�i�ō��y~m��#��=���ڑ3�$�W�وP#σd��|�e��Cՙ��Kk���t��]NO��d���d8���p=�J�$�ϵne�}��]m��6jN���}��l~MY�=�Q���P���˼���E}aǓ2!:��O�s��ͻ��ʠj�@&�+�~(����9��Kd�
Y�$�F�Q69QBJ�'=B>���q2ac�Y��)s��}|��!��>'��O��"L�ê��[�c�G�m���S���3��Ůk,���T&�4� �gÄQWxz}��l6�׼�����h�^(d��(�h���W�l��裻2;$#��g�@
��c	���N����9�*�l�� ��)�{�:���p�O�I#�t�����,,C���<@�����g�W\��A�)?�|I�2op���k k���Բ|�T�M��|Mx��"}�=̈(�2�aW�x�������+��8�o��s�!N�5�|��(.�����5����n���m�Xc�\�pHOK�f=�s��cNn���{�u		��J�n�-,MuA���|#q��'I�c�(#�K�/���z&���ߪ/2GԎ����Ĉ�n��I���J�vG]?�d.!H8�c�lhoo�����I'�� �^�#��1���i/��m`�kYj��	��p�&yg!!��Xb�~��}2��{_ǡ+�{�r���p��W�n���FP-?jF���Ĝ� �]~ɨ�;̓u	]{ak�B�߱},�z�>��������edn�`&"������ U�EG�qb�_
�9GJ�#��s=e�F��ÊN�j�W4����б�5�#Vr" �7#0Q�k����w���l����цh���cc��lO[Ϛ,�5�z947Ɣ����V�K����0��ʳ��"*o����ܠC���/��[���
�1;��=�i"�u|rCs�1<<L{9����HC}�0��E�Tv?.�$�?Oy�o3�+n�[����ț�i{�m2 n��Y7����p�㛜 �z~#��3gc�)��餤��9&�z��t�:ZR�V����G�3�]��;:SN�R`��^t��������s�	�Y]�)-�nnnD�C!��:�113S`�5:|OWUU�;ƞ���)�0�I&Ӵ��"�~�g��d�bPm4�0|<.�]c�C�CS}=ǘЇ�w��ȓ!�3�[9a+��ؓ/X|����=���6���$������s��M--#�x'QCta7��O�K���ΑkS��ODD.^�(S���2��8�НoH���*}�>�3�X4�	��kϠ<��J��h���+�<�Y�[o�d��'A�Ae^���8住��mt������n����)r ��D36��CXJ�%�ȹ���M(L�`: �OJ���~�?{m�gOc#��//,.�g<R�L���Z�^��j���'�cA��m������Ջ��P___��56(�(vW�xNU��١�͖�sS���F(�.wO�'�B����7����3�<�4$,3����OЍ���i���� �����fV�r�f�9�5%���2�A��T�&Y-�e�h�ވ�r?wb���F;b
�޿Ő���BMt���=�qYY�х�i�*@ƥ�N��Qn~��큨P��Z��ˢ���qRҘI
��G�_ �##�c���7���W`���4��W�$�x��#���f|n��˪�J8]��h���J�v�(C|^�ڶ��jг�y�����B�d��v��
G�N�T��}��ζ[I5Rz�]z/�n����
 �s�c����}4�������d��g��-�A���������rv��U�;
Տ��A��9�����[Ǻ��}�k�%�����x�5v��7�ᚐ��A�����+&����L�<JByͣ�@����C��	j��眢�0�#~l���#�z ����)�����n1q[��H��E���u|r��c��Vp����G"�+q׷�k��:(��A6,Tkn�ύ�Z�mx�����ш4�H'rHt�����9�@��f2֞_��t`��nw�ˁ)� )�LL���mo׈HH�������N�k��?Yq4�۸������(B|�n)O�iJ�vqBE�>̽Ш [9p��4xA��r�횕 �C�&��O`�����N�5��H1�w] ]ݝg�Atf򵏵��b�x-r�c��vŽ�N ɁG�`�; 
$yDhހ9�)	���7�|:h�����r���k�=E�]�QR
Z ��S�o���Y7���Fq�ģ厓��X��*���Z�is�;;���@lR
X�\[��﯊H�I�y%}d>�Ň��{�sOr������3COOLJ°���T��`<�+譣\w�q>EO��L^���G�g��㣢���3��!D3��&�l�/N�q3��=��*�6�47����?��{�Y�Q�ڔ����|PÇqt��N��@�5uu�wl��d>}Y>P�v�9CV	�D~�y8��̰~��8���/�99�	e��t}��w�#�D/q!1h~���3Bo��$�P�Hlll��M��}� 2P�1����m�(�gGF]ݾ#~ثAV�u��Vrŏ?�||�v �%��oT�Gm���߮:tHoq��p��8��b�����uu}�4��YH���u�d�+j�>;k��`*3N�Ԗ���uX.�3�\&*1�#�x����x:�n�������|���9cV	�1vB=�J�8TL�b ���3�A�@�ڽ���-�WA�� Y���wo�J��˨]���_�l�TR�]�h�			�D��my�s��$*�X�rНp��L�3V:-�l��2(��_��*���q���رN�x��P#DD��\	�>]�~�A�����-�lH2���+@ѝ�w陵�[��oe+����7FV��|�1ð����]x8�9�A�%����x�}��0�iq������0����9�P�����ysG�t�ɓ]5z�V�}��QL��
`�g�/j����Ȕu!��y���I)Ǐ�C}�XX�V�Ft�|�ʩ��C�Cz���"L}.���f/�������3V���թ�W#�m������J��b�s�D1�m(	��K�R�� �	��3�,�q�cc���F��hkBy�?��� �ş�y\f������w�sǓs�?FlHA՞	�z7N5B��N�R�C�$�rJ?b� ު=)�nrz�Z':c�Z�gW����J�\�.--=)��[9��J/w��w���(��#�X�i�_~GP�+!����X].�����Ж�'{ж���5��-�Kk���[�kZL�p�:�N}&ˎ�ˮO:��+�<�EFJZ���Q����S�*�	�.�%RT_�*�I�}��!w�ڣ�E�lu1�0I��4��c�DC�JX�Hu �2�SˠR]h7HA�����ͻ���|��c��O޺��q��-%qb��O��JG��҉E�ռ��X�����k8���^�#{+&�Į�� ����J� -�ڮ�̟?s�C1�5@��������y��
�K�Haa�z�J��k��:�{�٢��^(5
Vx�����fӄg�����)�c	1�>1Z�Oع��@��М��\BWƂN�:�ݑ����t�ܹ:�gJ����9 ¿�������r�(�u�s�=���Fe5:.Q=2�KI@����R˫�|XC{GGC��旕��tGWz(�u�<��(<��b`�'0���RP��sG���C6X��g��S��H��9�_���NH��N����L�WP���q����OM�Ał1�P��!]�9]V�2�+�u5�G"�\T���(J�U���妉KbVl/��h�v�Kv	?i��/"Ym�*�]%��N
��!�0*��L�lD�UbT<�������'�QS"�����-6rs������WD�Ń�cM	�_ �PbO��0#C���^O�b�6��ţ��^�xFO�3����N-�Qn=�in��$*z����ĉ���/3h+!X�|=�$�sdW��8�/���_��D����z-��P���Ꚙ�f�����@0��4=��'7����~��Hj�F��R�A�������ht�V�(E��X|�G����m4ᮭ��3񮯗�n� ~1t�U4�koL�#�mV�6\pvmJ�?S�~��eٓ��Q@A�U_�F��A��_�d#)�Z��k��p��=�4�1 �9|���F������+xy�̶`34��zD�&_�~�]ܯ��|%t��NJ8?�C�|�E%F�v�-0 ��S=�4!�AA�V��C���l���abFX��\�^yCT�u�ۻu ���c!~��������|��mj�|�C�m��-��=˴��d}��֎<+��0D��]Kj���2�B9-����G�D1Y-�����իW��|Gِ�P������Ru|�z�H:�rZ(V��nQ�¨�� �¥��yVr@PZ�-�c�Kݏj�O�_,�q|�G�Ca���r�/��@I*���]��6+��F���L�5B|�K�[����5���Ͱ�y��4��j�`���W3�ޯF��y���y�/num��)<���ϯ~���	wu�򁭔����Dd`+@�o�.܀���`I[�޲�5R+��Ԧ9�*gm��P�����X�>��Q��W�T�%��A�9*�v�A���Qů_e��y(�+a3��X/����?�r�I��*I�����0���;��e��+������K�%y�n�w�ܓ�=��S��wLLL��6�+%7B���jv�4�4_�1v���2�Iq�C�(�ت՞e��h�SN((�(����:nN�I��0�0i�
Hj�G�Z��h������Fm�pJ``���Sg;2�����7_ؾߑ�2�ٖ7B�#sz[��`���'����(�ee��ra�º��� ���G���-)ö��-�Jc�~ �ՅǤ��k �[��sef�2+��6s�<ljj�v�N�1�c�[~�M����dy�%+�`���/	��4��z�iM�V,��q��ͮ��~��U>O�5C��V�m|���|����=�?��19�s�ZrTRP��Sޜ���N�6��T�z=e�x��F���|�/
�(	����~R�Ь�g���:<��F��wxTwJS�����ש���$�n+�(~���ӍP?�c��&�Bi�����-��#�	����<Ǡ�趝Fr(b7@S�s��T�N���QV��J�6�&�(���d3�b����d���\}�S(R����9ȜR�O	�5�[ݘvLinV�qœԲ�Qw5�C�լ��(|���& �M�9 1`�������ث@%�v���؇7��7�g���.��;�U���cĜ%pC�]�'ʽ�b'644�ՍZb@�����4�g4�#ٙ�W�t�>A���^����w�%�?�Z�շnbK�N����HK�dy�Z��������Eս��cAq�
�}K�;+vB.Ǻ��������!렞�Ki	)�UA��²ZB��FVhE4N���@�9�ҟ��\ʲ�F�qQ�STT(���S���t�+W	ԯL����.%|0������ORQ5����#u%u/��+ U``22�����_�����xG�rJ-I�#�g����������8B�Io��@���.�����EGІ�����8hN�z������N�<�]��� /�k�(�#o�~)_���#q4Y�k��#J{|C ��m��K����h�
=��z��� @ę���ܺ��z�GbV�m͕*%d�i����|{{�|�����h)l���'T��m�lB蕇
;j�������]��)�ո߉C�x���ʞ��6�H�h�:��f�4��v�և.T��ӓr��7__6E�٦@b�T�ʣ�mŗz			C����$��h7Oܛ
"��a��Q��+t�b�;_5��˖q`R�����˰R��u�����d�\���s|������\����������O��Dh|ʴ+d���Q�OJ����+��29è+���q�?��9�L�`yf`lr��q��%=r?za���F�����f@@ P�C�g�N�M)�K�����/E�x�k`F��䌇��,��4 bk�p��ݛ�S��#*�v|	��b�����j�ƛ�T>�{N�D=�d�7���ߤvX�V�r"Uy�	Z�ǜ�$'�����ӥ3��J����c�XI���k6ڠ!$��z��Ot*�>;.���`��3�̄�@�C:����@�t)Z�^���
���'���!��q�U"E,�I��� Hх-��|�v��]4����\_�����|'vj���6s�פ'�R�-_RR���4�����`>�~�?�4�]�v���x`��."/	��	��� @��"R>�� ����F�Q_�f�FuЅ��qڿ�Y�#����w�F -���&�9II���鹌�����$��xy��̊�̀'��]�?Sz�L֧���LV���ɳ�Om���Lsr-AI�N��Q>P(�e؞~-�KL��)��T��pA�)�4X`��[R�@
A	��–��OQG'6!1Q�0ܤ쎝�_҇���JJJ�z=hioOpvv6��"wNHH �w+�l��@C�C:�Nww����RHq9�,�q_c]�^ZK����0��q6����4�O�Z֛��Km���B���G�'ڜ� ����/w��5��$&$�fs��:�2�UH��'�n�B5S����QuM͈m�C��"l*�n����M�ލx��ɢW�WI���<����Wkn��;8��u�ڃ=;>�:}�@ثءm�H��ڔ����sz��r%�@�R� �B���C�bo�U�d����K��N&%|~KNu�L �:l��<����c�_f��䱛�;̔�RPW�W�V7�>�_H�M�^Bv�2�s(�PO���܏SN*�,�ߋXv[���T�?�g�_A�y78NEE��۷7  .^���Õ��N��;�N��.l�:�1Z,�aʃYIPŀ6��5���B~oSR.HW�?011�D鞦�Ǥ	pi'�+������gY_"�5�Rd���䃨����Ea���G|*eRB��X���B�(�Z�M��`�_G���D��=x��L��	9��6P���^%ˤo�᳄-/�!r��Tt�� 64Y-;
ʱ��06m�A���}�e	v��1i5��ߢ������`�b�'b�;�c�9 x(�����t���!�<� 8�v�ѡ0D� ��Ы��$"�k�_2���>;T=����w'�*�i��1y��l�ϡ�������74��#c���J�;���:0֔8 �5�9e8DO���'��ْ�a�\:t���7�C�|��R�/�@e$�<q�壘��}UZ]V����"WL_�]P���..g��
5uttZ�~Z���Flfs�7��E^E��2���/Cf�OK�/-��~��;Z��q�5d��;j9EE�����~���_%���A%
L�d*!k\��U�{J>VS�J���jEb>v��3���j��0EԎ܌�����pVf
��*���Y��ݩ�<�߾}[ Q�*2N�*�Y���uy�k�5@� a�J� �H���&/[8�����/[O����aWQ.(Z��Q�?�Y�%��h[�r���oz��h��'#���"$�����UODzmģ������,m���B�/��|�D��|��Ѝ�b��/7s�ߧ
~)o��H�t�{��@XĜ���T����4�໨(ZTa�|ka�bi���zrϞ=��FA�2����L��L��4�F��1�r,ʯ2�������>��蜝��Mpp��Q\D�'�Y��k�8�M�Aك`�0>��F�egy�=�0A[EWQ�C���Wa��~��c|a�˲'��CO"P��������{��	���(O�C�y���߉���=������P9���M�T?RRA b�3�YA�>BC����T}���0�4gi��LEz�J�|"��LWW��S��UEw��*�o�9�'e޺}�'R������c�B=yx�Sߏg^��
`�s2C�jc�h3�L�+b���Z�L��Κ�!�	��T����������B__������:R��"+�ݷ�1��y:��31� �@l�HM��������w���?7y����4��Nԕ���,�n/�J.))�)ݠ���NI)aӫ���x��v�5���]�e�3�SU,���}h{�����z�y�������1�A�A���} ���WVVFg��1j���X��`?��u$a���:�ہ7cIv�3M.�6H�x��'0�Q|�yF��U�4D�E���`	����i�����<�Gю;����V���(��9�`�P.�����ee��b�-�ey�c�A���8�3
\:66��`�5�G�X��|l���Z�+� Ғ7�iF����������I(�A�>�rNj�@(����u��R�$�]haQ8�k�-~*�0@%�V��vL��h	x�X~���KJ������8^�����Bj�=�[��~k�����^�Co��"_]�@t6����4���՗��)�W�K5���fc�`f�h�Л�ٵ�LR�4�ڛ����3C�w�x�@ر�x�X�L;rV��+� zM�T��'w��˗��9���t�jI9�]z��X#j�(�O��������=L;~r�]�Ә�e��)%��v=�Rx8U�#㸞=��d�@� Rb���^w���%�͏��g3;�p�#c.�-%��(l�Þ<م��+���-��p��O�K�S��$��Đ�Gl���ag'�u �����\O�^D?~�3���C�^��y�������춝��	{�'A��qff�׊���&�ik䋼)qV6��M�������.���`逷�"��\ꄯ��羧!��K3��e g��O{�cW���߬� ua�ʁ�PiA�����v����7X����*:�B��J��yYL3���3��u%Cm���ϥ��W��������:ᗢ~C[�Dr�Ŕ	���iء��,��a�V��z��u���P�s�)�,�P���"�8�.��Ѱlm�0E��c{-����y�g���N�$&��OOK�^{����ma-%�|�ܾ�{��P�M%�`%�2=''��R��E��'���
���F5�Qt�D`���[*r(}G�5�9�%板���,9Q��������P����HQw�4��X��iӢ촐�)�Hd�6��:���D�۠���"[�d�B���`"&M�n���}�������������s]���y�s�s�攚�e �'Nq]�ͳOJJ,�`0V��8�&M��S��wϟyׅA�B���{�H4��}:t2q�5�uu����7﹤�s{��Ś]e�{��~��܋������.�^C�O�ޅ�}���C��?��ߋ�'f��+ݜ�?��
h_�\|��|���,,j�[<�t��F�o��׿���O�P�I�	���
^��OwA�t����"�|V��{xb��i��N��
.�9��]�>~|�}L��-�!g�B�|	����q�����Skk��}�i�������;oL�>D��fU�c���p���"_±g��f��K ֑����޼A���B�I7��ߵy�1���M+�x���s}vh�2��]'!q�̻�|�}JJ�ϟ�rL�o�_
��=��s#Ӳ$��>��$�Dz��mI��p���m�>�:pP��?���.[������~����As�i��+T�Y#`�Ho#�j���/��W�������kfM�Bs4š:7$a�����#ϓΟ���7�Zh�e��?��4Ȩ��>ɱU�
%W�pGY?wh=��WY1̞ff�V\=p:n�=ڱ�н����Id�y��|�zB�L{��$�[/2�t�t��+t�<k��u��eK����A N7{ʰ�) ��`�̥�{+%))��ҩ]]���/aKu��~p���W�*WC��(*)1��={�2-��q��2?��{�n�)�$y�bR��6�h|_�숊>�A,+�mdl�g�Rǩ�b���@��'O>��B���3#�%�����R�"dn���mϐZ$�<L�T���7)�j��><�+�ܵ�ӻH��?ʴ��j��z�/����4$D�	���v�+5ㆇ�;���_U^��ڟ]�A&_��
��gӿC��3����rh
,��>Ϸo�f2�6*NxoLE��Fv�@�8S��,6�[��NU�d�+*5�T�6��Ǿ���쮧�ѩS�������o><��)t/����B�f��-cx��e]OoI9��9��Xwp~��	_M�I�n�);,�<�����3��NΛ(pd���i#�(U5����l/u�cf�)�Axe��Nq�[Y�	���#k(�V�v��\V��ٴ�Pߡi�aYl�b��;3�ЪȕKh��u3�\M��E���χةCZ�_�~���ϒ�`i��/ڢ�t�!eI�?P&���%��̓dOC��n��O�d�]�Ç��� ��T�sI롛7o�}?jQ�~4�<�[�y�҉�CO�6�z�z���Q��FC�����>��=�~�a�;���^g��]�S�~vV�Bt��|�QĆӑ;7[��9�b7�����1�Q�#�I�9g��]��5��ĉ�p����7G�bb�_�Pܱٽ5�3��rc:;{W7c~ݶpv΂B�^ZZ�"��k�Ii�%T?;5�R೑��"�FU���z&;�����bˬb�Yo��>>E69�Vo7���M]BB�_�屚~���y�l(�� sG������%��]���}������\�Bh����EP��rAn�~����""��3-B*m����@dN�U�g��q���P�\h�oim���˽&���T�.�ϖ�H���[�O�Q�ir�h������p�����:��A���R��` 2PRp��682�ao��~����<�ݏ{�5�䷛4��A/�;*�Y���,_��6�/�,dMZt�O�c:����ʭ

L�K�i�:�'���,b����&�S�E>EE�i�Qs�_�L5`�״>2���l���_{��;�TAT��l:u��w���@�uu����N��P����_8|�S�����2�x&���
ܦF�F��]ȍ���H��]_�7�Ե���,R F|懶b��{��rЇ!{��~Gh󈩮����C��_mf���W��|F�<c�~]s����h�p?�W���O��N�������eq���b��5��zǻ��(6����%�$^Y��е�W�F̍Wm^�����q"�H ht���F��X�����U:hB{g<��|{i�z��fDZ�Hy��f��l�r���,���F\O��0vY��/�S3(o�\��\&y�.�Vj��Ϸ��ii���L����/��c��Ɩ��VDPh��
C�Y�l+P��I����ݲf�(��{�U;�<fD����ŴިrZQf�s+t���^=�l�*պ�T|�DMU��Z�,˰n׵�þ}Pୠ��n_=�d�\	}bD�e����I�[x�p�z4[-#--�0S�ٽ�5����3VV�oֻ��m,��,+K�����Wf�9�����g{�f��x� MK���5UUC��^~F�Ӄ�� �4{T��8�� {j���.���_�=���Вl
}u�e�ʯ�,4ڱ�MKK�6��v�J(�˄���p�no�b]ج6����:h55�YU.t��7*kMo��j�x���ܡ(�Lh��jv�N�b�����}zb5�C��>."x]�͒�\�&kkk���y�ed���S0�,g�%�r'ؖ�,��N�N fF���>"~uX�5�kѽf+��Bn�,��5������Jq�,�jr5E:)ŮP9'?���PLD_�Sl�-��J𝬌����nK�,>��ْg?�|��e�������عxv�9�b�%�J�b�@�����0Z�QɅt)-O)�FZ~A�q��MI�������ʗn�]k$����H��;vUGmDS��T��Yi[��"��]�ot�1���Q���*�r�q��Z��\�M=$�g�t[ǌE�agl�����b��������kb�f��+bD�˽���f�ie�EE>+ŇA�Q,U��%[B�|�z��@�������d�-ǾK�p6�[���T��9�|2�on|E�g2)�8�R_���u���!_�[Wӽ�fʍ���WS+$f5���ʻ{� [��	��5��J��+�/;X��~��xz�}�kj*�f�N�H:�;�:�	Z�\�<��=3���/xU�d>�8\O�,�B>э|���0y��jϚe��1���*��N�)0�I t�|%,}��&#s!���T�GQ/�Q����;���\��\,B��ٯ�d8�m6����3�����
~$�W�i���O"	2�c}�g˂��G�$��q����X4�-�l�<�%��|���EƖ�k� 8���_�~��RN����C>m<�B��o����Lb��*9ш�ٝT��	�q�Q���J��ጮ��ж��dߥL%�� ~ii	����\.�=;���?x�(�{�2�������l�x'�`1�Fŗ�f��ƤYE���m����h�tS�K!�tg���#�:��^�,n�����D��v���P�A�
��K=,h�ۀǭ+p�Ӑ�aI��*u�~�q#�G�N�퓏J���jEW;^�M�Hr�K��s{n�J�dv<�R�,:~����s��z��I5���t�.��~��r�
�x0OOŔ�ҋ�L�V�'���dY؟��R�/��������1e���W ?�Ft~5^�����v��Xx3�6�5V 50%��(Χ�꓇$���F5�'��c���%�@�\��G�bl���[�4��8n�9`��jP�El-���p} J����j.�}�����lΪ��S�!�E^2�\Mq�Ʋ0�7+mС����X�%PʺDhU].���ͭ.�gǜ9���-����557w!sg$h����yЕ�뾮9�*fb��.V�&��Kw�6[i���%���Kmħ�B%�vf�3)I�]���~�7��/��+�*/Gr����es���y!��?��;�J�d�y���>ȇ7a��V�BB��+/����S�V�#�}|�fg�9��TYI;i h�D���>,���?n�.yQP ���~aC��_����&�=R��|��*Ò����]J��Gd���L�Vȣ?��.=��}���6��b��w����n���g��تTFC����ujB"K/�i�����G����P{ׯ_?8�hP��^]�^s�Y��?�oH���5�-X�WүX4�h�#���J4�E{����|tl�U5�͐宋Xh��=D��s�F�^rL��l�3 ��PW�+���׋Iayyy�H.�t�X:>P.�Քa6ؠ+�᥼F4L�,�$Z4�Z#�������[�+>{����]�����1j#_XE�)t���G{�#���^���h�2�����^�\
+r�5��?�#:�#4C �h����\yb5�)�zlտ8Ut�T���%��d7Yn4�4�mq��0�볱T	7o��g������3���"��B>�
��j�g�}`;�p'��H�w�����ć��}�QQO� �S�q�p��vW�@˓C��������U>�`^�P�V�!�1�"�*K$ދXB���A|�v�`���^���]Ǭ&q�J��s�����ٹ�����Om9
�.��<�@���=��h ���jAo�[�ԋ����W����ע��T��Ϙ�o�OGhXX�������,'7Wᠹ����\`��3/�1I췟^PRR"��p� �*�F;0vq�7�GD��fc��n�L�`Y����Q� `
�T��>��A#����xQ��DXU�� 
����͍�q@���@p=8��%뢲ɝ��MsS���b9�-AJ"]?kd#>�"����ѝ�j�Z��?ӳހ��YKۅa:`��г"��{����Jk�f�f��q���R���nk��6y,�~��c�xj#Mt`�f�ޏ1<*d���K��C��g�I�h��<�t�P�������U$��ua��0��Te����:��_�ܒ ��ljߜٝX��>V��Z�(Z�X�y�����_�����~vQ�˗������L�JOL��Ҡ�qFd@�C�݆��|�6/o�h�����Mv��l��1�p�
�1�I��6Z�VD�B̵�םxX����DT�f|��I#��r�@�^��y�3r+yK��XA���Nsb&S�2��4,�]A�1B�'�Cۡ�ܮ�213Cڤ�wڋE�pV��ݬ��E���-5�o���9o�9Ya��*��TV�Żv���B���$�pz_��4÷[�+��f���8ͭ�2=�t�����y��g�M���Mn88��.Ls�
�����eB��k����&-���>����,�Zjg��9��!���,��C�`���i����{A���\5%�[�TF`1�CuXk?�/ x]���J���U�9d��f���]=���Í��a���"��-!28��`g�#�0����&g���W��NߛϷ�"�e��&�J���ţMfHJg�N^F>�>b������/���N�!%���uˤ�����[�s�w�::�`���D (!=��v��:&OC��X#�g �E��}}�(�o�'l}D4�j�RW���C�M!��jܐ*��35/��zB�[�T6Q�&����F	T<3����q�=�L��*{�2z!k`�989	ZrB��Sj�c��M��U�[w�M~q�����:��+{R� �Z)c톱�A B�X��Ǥξ��p����xvH��G.��������:}��ę�2��*d�֗�ȤN����W�a�aF}U3pj��_82�Z���-!03��0�e��J�f�;ھ4�I��J&Rg�.N�|�~SI>�	����c���s��A�7�{���ПiQ�Y��0N���|Z1p4�����^�fBZ��6��hbzbx�z[V��܋ə�V�?cR7"���/�rB�taf�ƭUFFF����+C������w58��a!�_��/��N����RȖ�. ӻ���|����A �Ρ����&R�nZ��[�!\�	�eMDx��C������H��E�E1������g�0$�8a�W	��/�]��:�C��k���3NE����xa�Կ�|{W�R�m�߽2,+���(���Č��0:������j��eB�X!� -(_�!��v낏}[����aA:�z.���WW�Rg�R;�H|��ya�o��U���+r�V`o�a��MC���^��V�
YD�b[�ཙ�AY�X�di`Z�͞��������{ȣh���w B�r@�Fŵ1\�O���� G�K$��K|��?��t��X�h����	u(�`�!�Pc�w)Y���s�D�	2���$5��a%>J�VeRHW���G!H�YQo{L�B�R.�g����Ճ���7ЖO��KCw��-�ҡ(��OS��@ 1.ž�R�1&!��)o,�Τ6R��<iYV{	��m�1�@}�H����{��v���T^��:�P�����U�[���@k�Zc��V��<&�_����$7l��p�gU:��a�*�Z��PA���_�DLf��Zo~����{�0� mq5�*[ qM�Kwu��,�������[c��$D�󽁢ET�2-��0&5��}�E�%�l�	�P��b���،��z��h���ҳ϶�C��YM���#B���~uXmd�=�%P�I1,X��|��Xy�"�7�2����BVA#7�i���ۅ�n���?2�
�&6�6I��T���R��s[�?�
���T���Ŵow���J�����Y8v��p!�֗�{:�Y~&��5�6��06�V��}�-��+�I���Q�������s��;N\zCsy��d���߭=�oρ�����!�ϙ���QV'���6{&��c���㥁 ��݉��"U��\j����ˣ�!&n�`��oe�@˽?N�a�I�/QD'�@A�s/�Eh0O��{8,�t�������T
����j/4xX�i0�=�)��;��mr>LZ@xK�ݡ�`5ǃ�B��<U� g�󓰻�84� W�B֝���s�%O��s��w"��{��r���!���>�i{y��V�!��W�F��a�L>�>MK&^؈n���zM��~T�ݣ� �Zh�a�9��=�T�]$<#��\�{�RJE�����!��P>����U�9��$.�F����c�md�Tll=�AQ���zx1�a*��'�>�<#U�<�����r��{�zH�J��>B�~�p�/�"���r���������@��w�W��pؗ���o}Rԃ}�6���8��IdxσyZ��|�����_�kYs}O��Q߁�ۭ���)�~3��H�/XB�v�.V���{>{o#��#%z�סd�`������6����?3��BJJ4\��O줔#�X�I�=�@	�6A���Y(�����7��ӚJZR%�)iis��^�!����S�*PwU6���x>�})V����|1��rix�9���z��(J����-�0W��b!c�R��J3<����3 psMo�#4�t �۞d��m�Sf!��XAyP�����<G=�B|!���E��_Le�6�=Fhm��������e��E����=��{y��c��������Qb�o��掦�cr8��|��Gx	٫j�2������V�Q8��rU��w�W�(-�/���E���=�@0��^AE�@��(�e�0����¨	0;�7o��0<\�� U0��\��5�!(���N���-�����PT�E�=�B|�*�Y��Y_�������h_�J�Gf2m���u�x'8 �l&.�
�V.�ɧ���\�)^ (-�ּ�������F���^Ed����O}��V3*:����w�"��l������\uW]U �	/,1� �S�Q]��b	x��M���R>h���9�KvWk��U@c����ۄ�y���Mqɓ���ˈ~L^TT4ΑO��[���-�ar���PQ�	@dlT�@�KE���fm�3|	i������x���T���;)�V�@�WP �a�H��!j�P����"���e9�Y��ɿ�e��JONK�G��j�Q��3[Ξ����z���� ��/Bh�&�"'�*6�e_[Ȣޅbƀf�r��O4{ ����ٖ�j�s�Wj�mZ`$a�G������$��p��#ڮ5��oϤ���$���&�s1m
�q�]�O�.��� ��ٳʿ��\��g�� ǯ���^���\�9P��X4�,�$��[N��E3 ���V��!\�Ҷ��*&uˢ�?w�4�A��,ּ����ݖO}�1ߑ��+,؀�|��͚����u��r`T����OV
.  ���Ѫ�u���\��o���|���^�#"U5ፗz8�H�(��g����,��^A,1jF���DZ<�<�0J�1	�7M\0���<V��ym{נ2ς�b��FF:sA��,)���,?��� �N��OӶB';�T[C�y,0�}[�&'���<��d�XHY��,��ZB�*(���+�7b6� u[��%r�6����~+wQ�d��f�ӷ��ʃ8,� �j�;78O'fK��, X�L�����C���?�E�nw~�"��#B}&�&?�0]C��d���']�q�1����V �^{Zw��Ql����z�w��B:��(
,������!����'�Bl�
��e1�<���,�£���ַp �``�^�푆%�=,t-��nf~��R���"�K��9`�[��%4�v"����D�	i��ُ m�K�����N��~!PP52�F�v���r�5�FǢ���E�
O�H�pl b��F����5�@�f!x 	�Y ���fH����	��* G@S�b�-(v�ᒁ{R�?5%DDm؈����A���&3��[P��%@�Q�I�%�� �,�.Q(_��w *	c��EA)�k�>��S]��⊢?E���o=���2U�nOJ�+��z{H'=m
Lbʍ�E�؞�y���7S�P�A�n׉��k�\�-!���P%�D���S�� &�"&���_'}<��]1�$}�*�Aޖ�pi%�t$�$�b���>�,d�qEO$7H_U; '�ٽ�{]��5�7��+܀~�O½p�Y�W�p�/�#,m��Y++_�'4s�@����s��Cք��!F��KKS��޵F��S:�
������G�7��"�S���eEb��PD�Vpm�Ij��,�Zw�.��u?E�,�/E�d2g����L��-7�n���P�b'b�)�"pX��"�け�Ra[�̶�Gܼ��{۞� ��'��hP�ٓ|Gί��c�Sߦ�w!�n���5�/��f:�4�V/��#�٫!��]�?ձZ�['���� <��+�*K�K4��BJ�QQtfvfi��~Q�?���n�1�̜y��F�޸�&0~j���5%�.tp��`N:\Pvl��%��Np�U�r�".���%�R�1����Z�U,a��7m�_�����L��ۨ��̊>F��h�hK�OS@�UH�N��N�8��Gf5Qг�tY�&�I(ݳ��xm@����������Npf����t�6o(ż�PX̿)�Ǣ�|/A�@�����B��hy�'�7���_L���"�� ��D<�w���͎�>�`n�%�Z���p��}����uut,Ü<|�Ù�!zT6Z��Ӛ�XD��"F��Q�FA����B�=p�^��=�@�NN�ߗL����:��m��<��psԹ��;�v����0���;[�k��;��)of��H
oN���1@��3�<+����<�n�o �<��3�tͳ+n�����)����4������?h�ߔ�M��Ԕ���vi��49�����bn��N������:�<������m7%Ο������o��/M)�·��*50��p0�^c��^>
W}��{�C�����Х�.d�����"99٫jO)'xw{~����}������1��C?�#�,^~�<����	~�GUph��ck���ח.]o�̓�:5�}!��G��%���em�GS�SN���ܜ0V��Y��gZ(��gu$�T4�M��%>���]��9.��GA�}�h���v坾��YB{�v��W�B��c�������~cᨁrҡ�16�-���'�,��1��6MZ��{<������ڼ�Q�?���>ބ��?�3(�稷��N���x#������`�k�k�����8H���U393k��D�XL{���;t!�2��6��x�3��G�Y�͛����Д�n��w�4��O�%n3��J��|*�u��v�C��L�4y�}R�w�(�K���\��-�wԋ�&��tV6������Ŵ�OI2|1yO$A�|S}��7a1�x�W��,���Q�&�חx>#�
[�O�7a����.��df�I	�����͙S.ڟ��2��{2��X�ЩX?/���Us�J��bӝx"��?_�7����� O:�t�k�E�����|�}�R�D�~
�S���?
���(XL֋vށ]��~��%�����ze��N���3�C˿<DN�^~n�m"�u�o���2���ny������kGd��y��Ky7��?�J�����?���g��_<=�kk��ԄD8� �>�SQ�	?��E��uM#�\��}�� J������)����wZ�o��ۏK
��x����8r��Lv9#�+_��ZB�]��PP�m�ޡ���D�c`�������Ңh�)w�ܒZиvA�a�$�?�%���.d�W&����ʫj	�bX�y���ff�@�V#�$�X�eBƲ���Ft�T��1���NyJ�*%�N�>I����E0�^,&�}��?z�iwKEpt��� �q�l�3?<<�vtr*��= 0^�q	B��u����o�����.���r>����q7���,������7u,ڌO5������Q��c��/�P[�A���Q�d��HUB�?���t���*A������L]~;��wh�h���x\��ܼ}֔V�8��t'�Wj_XU�$!K�e����%/3V �˯;&��A�ǧ�6a1
y|�v���ڻy�~����n��sU�b��_�M/�iiq��"}��7˿ՠ]��[�8�ay�̕�Q�1�/�H�t>���!�Qj�Ӛ���}@���os�ip����2�Y��������F��>�n�Y(�Ï�Vp^���`@`FYoT"W-衆�`�����i{���x��r4-��9ދ]�rO�l�-���s&�����du]zެ?���z1���a꧂�"��I���~�d��2^RT]�n6s���zM-Ai]��#5|lGq�����r�^� N�(���#��ި�H0˝={���wI{Dy�d���Ӽ��#ɶ��%��^-a���l�J� ������8,�J�Em�6�n�DM�4�t̜�n��>�P��:�5m�����D�KА!�B����u�)�}-���T~=~��U�ߠ$���_L!��S�5i�%P0*t��G��D*e%:��E㪷���_�y�߾ ��BZS��&�/������tQh	�J^SVYЉ�k
���x5���ua������'�wp�1� �Ŵ�Gɤ�����.gXٗ��!:w�Y�[q�xϾ�W"���K�a`�u`��`�,�
%~��ؔ�6��_��+��_�~�~n���]�z�,//�9gi�hևf���,ֿ;.F�[sY��{z���B�I;SS�� {{�g��%�Ѵȥ눃�c^��q����o!^8...��˯�B�β�����;��F3_[��zG��Ƿ�]�G�ߓ#x����g�PЫ�0��#2zz���A�6�� �\���55���f.[�
zC���Z�#��`p'��9��a�1y���I��yMj�J�i_���N�[�p�g�g�-d�Z'jiWD��Y���Lr�r�z�Z}Uͧ�4��o���΋Q�/zc�'&&:B���a�����(-�}ݛi�ҕL���V8���3��i݂��v=ƀ��n7Xv$K��̉ϱ�U0V�ēL��V�EeƟ#�SA�Nv��֨&��5������N�|��/5�i�kwuԶ���ZV_��6Ô5x/|!b�;�F|�A��^Y���S4%��gS�A~0ӺX�4���=p�pi�=���0�����e&� �TO���t !�Y��t��i��$�LVv�qb��G��G�î�=�C� �>�lr��������|�4�F[�,���5w��yjTXT�vw�yvW�R�R��6����e�wvc@����NiM�`ɐ7q��IȆƞ��23�h���ր�f�����gr-�g�AU�9�aG�c ���+���v@��h1�ѝ��3��U=��H�S���!C�X*�9���/�Lc�@Y�&�X�W���U���I�}��ZZZB�
_s/vuV�f0P(�섩AV}z�y~y| Xk��7�͵Y�CXd�*䁣�YH���=}�`�55�J�@���ҫS�~S��I���U��č�y�<i��1�i^�;�g�5�5T�83.f��6М8����hݳݛ��5X)�<����L�t��q>}8,Z��5�kbi�^�CM@�ib��K�&�cl�܆��0d"M���f��ԅ�����V����V�2�u��+a鹝Ú�D��� �	����>9�o^���5X��������N�5���D��ּ;���6�*ÜU��0%��u��.�hfV^��?�)Us�ҥK�>-P����|+QQ*n��7c	�u4D���0��Q��Ty��h��Ma���j�_y���Ȟ�9�����?�%��X��%�ld
u��>����ߍ"�~�7�!Xs��8U�']�>�>��q3N�=3Ů�ג՚�'�P=wl�^�����xX߼�{T�߀.B}�$/slj�,�4y/=�L���E]K+`�L�e@NϚ��Ԯܤ�g�2G��t!�D>�^6p5^�_���~�2:�3Ͱur�]i�JN��N!�>�<�L���oAB�����&Cw��Q�2tْ�SX8������L���ʛ�6,�'6�]��q�t;�^7X%p��u6ͭ���HSd��/��b��q�:gz9Z,�[��l��w��MK�6�H-!�H��1:��؆��I+WK����)-���z)/l-T��f�l^�vIc���� �,�
�;у�� �&{�)N���5Qtu#�¢����X2�N}�gw!{H*++�}�}�A�@V�'C�<`<����3�JʾX�b����2=>��
_��d��B��>}���S��ѬQ��Ǥ!{�K���N��k��֣< �=��ƐH#G����).�ye�I�[����KQ�~�6q��S̵TI�M�	�����~	`� ��C��_Z��<{���Y �];�^mМ�(�JK}����`�X�E�p����m<w`h�U}�G�܁��Ԥ�;����-=== `�$��6��s�������s��}@�3=n�'�~���uX*`z�{
���2Q �^G����(���$,�F6B�#Ѐ����.C��5�EY��M����&|�U�I��)h𩏣pӄ�]��W�����Eݟ��W8����?�O��F4���A��(Ih������(7�.�2��P#���PY����2�׳�>l��W��!�F�ͽ�(��3�	��k��¦E]�_�~��u���+}��1\l�t^m��ҷ�(�䬲�1V�>�ϵ���n?{z��C��p�V�����7�Q�r+0��r��3����a&�9�rZ�OB;�c_c��H��-%y�w��߷�~Oc��AF
E�P�`=L�ꃶ��"�څ�N�0�Y��{���[��������m����n/ŷ:�ܱb����ML~%�pp������(��[�˺��Rʍ^8�Xi��Q�5��C��%�%^C�I�j(�@�J�12�������(�}���!��-k�K���mɟ��-��W�@�I�hF4hf���
�.�TT�C=��$��Q�ԀV�k��F�R� �}S�
� ���m1�f���V�t_�$
/A��Ð��9�L�)��n���[��IHJ~�G�]�g�ÈW��S�)���^{�OЃ���P����")3c�`A�tK[��T��/L�ϩ��p�rBMM-OE�P��1�҂�YF�6m�<3��z`}�rXߚe4�rQ�V}9��9�s
_uv/��j���Hp��ڂ����gA��c�jΙ"�2Q��UfM�����AG��e;x�(Q�~��*�6AD�Km"�']�̍���6fU��P݄�1�sz�d��k�5��@���j��=�U�dV�摻vU%@EWCĈLi��h�?�	7����2��
�V��1=�Ll�ѯ��V�ڲg��j��TR2�c�4Zw�<^�PqK�ak��O��>��ҟ�ּ�
����u�����e
2�'�l�$�4�?�9Y$ؔ ��VVF�8�Y��o�}�Xt��l2B��Tq|*�G�/Ͼ����K��5ss����.�ӌC�D���@��t�*[	��hǾ�|g��!�$�O^������I��W �,�$U�$��/����r��O�}��f�|v�g����Q�@�(�G��u�-Wj�������}��h�k�Ǧ\��{�� UN@�;�tkS����^U�L���O����
�f�ZWf^$�?
ι�b�
'N�;��'�Al���.�q:=F���߃fc9�KTϹ0\��t�ji���|�@�q�ӂ���;��s��� A��ck)��a~'Tɓ�پ�>}"_�@��bS&������1lT��W���XL�:�$���e�X��d�j)L�ٱ��}ך��2�!ٹ�1cu+��'i<����<�T��~�����i��lG� i�ް(���/���`���R&r��08g$*Ůt�L��w���� � ^�p�e��c,8?c�ax>�Pk�|%�*�&7��؜Q[��9�'�>���v�'�]��sI�Af�[���Db;��B>�px�I
I�k��q 7NE���%}�˯@�(\a�c+��Sؚ.R�A��}�"�/
��'���}�h!�Ѷs{�\ў�����2��ln�Z`=����h��
tғ6�Zq�$W�%��h���7����Ӛ/��)�%��צ����dZ�~{}c8�p`�K�]l�L�+�����"��~=��u� ��i��t���â�r�p�l�j��t��V$��R�~<�*�Ni�����® fMߋ�����׭���K��T+���O��Zd'c��-�	�����n��3��JNf}��kOk����m�n��-hj��hv�JY1iȍ���� ����S��5���{/�9�N�
�D-Qa��T<�\��ZF;&!!q<����-"��Ϛ�XL�cz:�A����B*Z�ZC[������{���l��#dZu8�0�D$�m=��e����k#�T��M"R�p�!R
p�z@<+>�xӍ��I⿽�h�H�H�f,ӹ^���S�h&@3�N� ��k��ӕ�'�[�9�	����@]���S�<p��x��^�1�/��/��K
�ӽ��'�)K	��7Z^�ӻ?�Oo��P\ʕ��n�̶�ї�Fo���+��O�Q�,sb��<]d}4c���A�p"ǄO�p3Lw�k]��LO�Y ���ȩnu
Db�S�!�~$�;NUM������n�Ѥ��/�b3@�<~���mڨ�6_E v�H���N�2�^�k�؇�?� r�6�F_g��ޝ|d!�:�5��bGbG�?lA4F���1�����u��4o8-��
���L���	��EsI�c�t����`�=z�ś������ϻA&���L���-���l�!���Lgf�^��ͼG=�e���I9U2��M����:�,(�|Q���.�[�a�ID�'͎��r�$�W�/]���]��j��fS�u�E���P%Mz�9�������l�N�.�Y8�q�\��U5�����0�s��&��_�?�N��^��&� 0��IS�|�6�7{��]��Z�d�N��k?55UJLz�j�Q�3~���1,#���E|�i!�H۠³y�ORAȞ�V̳�߃�LQ���U'ARކڦ�����p��kEH�@�m����+�zj���ܾ7�(�G�+8�C����ҪFE��>ݛt1ݣ*��� �Q��'��i���deHr��@V-�ܱ��z�Z��2�ո����Ya��E����Wt�P2�Rj����.��|���h��eT��r�&c����X����i.""�%^��ޝ�ƛ�H�A{~�6�3�g
�z����A�G�m�9<'����h�����-��YK,p��P7!��� S��{� >$�[�=c�㉤�bQ�o���+�x��TV�`��d�����	��(�u���vq&���2�+��Ϻ�h&⪨�ʞ������
�tO7j�xq��>�쏄8����u�k���~nE̋�y������ q�������J�DYFW��f7���~��s躛ڳ/��S7�J ��F�z,�B��Y�R����B��"?��\�j#���{=h�ǻ�i���d�Z�Md��IY���f��=�e[eJ���O$�h�Z�����3������g��?�=��d򀊺�ff���K<f�*p�юաVέc�ЃZ��|�;��a����4���ܢ���20�̜�~vY������N���!7�<�Q7�8��};"qޞ��>>����t3pX�8�R{��4OQj7L��xT3z�_�8�g���s u�h;Cy
�[�m7^�{cl|��#����}x��S��VE��.��<���B.�}��Jl֩Hs�\��Ɋ *Ԩh��BeB\�,UaD0���-��DkY�B�����s�{��T`i�v�?n�D>"z�	�8A&}\
��Rl�1�B�.H��� ǘ�6n3zp�/u�E�X
�bE�4��>��~�J�
cX�1�䞟���b��:�',@��s�z��1}WMЭе�9*>�)�=7�	t�3Ʌx	0���K�c�*Z;�#���}�
؎}�2�VW&Ϙ.ӭ8۷!��]��Q9�B�T*+N	����qjp���83W��ّ ~ϓC�/�Kr.�7��!�O�w�R�d�dq����}����&ɥrxɲ�h�УQܕVH}E���T�eLגIj2�zP��������v��l���
CI��"|,L�M����Lf�%p���6�Dg �w��5��0kɟ� �.C��@� A��
��)qk֥��"�$����jg�@��#y��I:4���Y�Ā� *2�ھ�^��� _\H��� ���j��U5���
#�61����� ��M&iI�2$�w`���V�I-�J�� �LR�����%$�Q�I��޵�`����<���NB���ND�0Z���ǭ�	d��n@�֏��I�k�͞�t�kW�g���Xu��_����j0�b��:�F�����K�4�#���T���mܯ�<x����#���2�`Ц����?Ae]@�����\�}�o�S���!G����
� r�����]܂Ԩ;T	,��6m�B^spO	ZY�m�n�, }�f�}	�{�H�w����ߖ������!����D��f/i�Z��b���f��(��ϗG�H����VAB��ln���%�?���뵸����@�b���9ovJ�N��䑞n�	���Ϋ��T�$}���� �W���܋e٤!�XI�B�H���S��ЃM�q%9inE&_��\��uF|�^�?�����i�'_�nuvH�+Ю0��X�.TA�B'� Ө5��H�"�VTTd�^$x��vŰl�;#�S��I����Cq]��jB�U��k�q��f�! ��t��wO��T����a2��Sa�v�k95]�`&�5�Ї1<�p�⹫���+���]�&�G�����B����{x�k�L���c�-�.*����[�X�RzC�����V�Nh���yQVƁ a
��b��ќ�b(�IG�pX��;�b������e�q�"٥�1mRh�ź�����,���eJ��h���%
���}�,���vq.�����q��wR�B�J�h4�	�}Z�WO[��)�Ľ[�� r��T�`1�8
��[��P�!�ֳ:�N}q.��J�OԘ"���C�:��H&E�}dlL6�y�E���������/pj�L{��s]T�m@O��rE�+�e:�bf��!���<��4�8oSm_;m�2Л�Ye�'�L�-�}'`{c��S�wyYp#��*j�*&�j�/�!��9WLw�l�S�� �1,� ��
3��j�$�Ǿ�c�SQ��-@��i�n"��%�_j�(3�N����xiKX�J;���`L��!hOv2������m333
��Ѹ�� ��8o,��]�Ӎ��]0�ڿt+�]�&����|��zt+z�74����J���h�G��� }L=�I�I��޵&�l�9i+Y]1�^:d�RTxhX�� ��lgr�t�z�Q��� y�����T��c�Z`���d�"�b�C�E���u��
�'*���N�TD�Oa�Q��!�t��?�S?͢t���u��g�Z$�E��f�'�橡�G ��w�X*�,'_�����a��u�p���B�2����-�O$rI��s��(j��DL����J���9�CN�E=����)���{,�`���B��
���g=;���w���K_?A��3��t����d�弐L�~7[b����畗CH�N�¥J5�ȋ&U�&�\\�&L�Pe���҈$X����4����?D�vi��U�4���!�APA�%a��
���	�q��+�"� Р� � F�$�������eWM�TMM��?4���}��s�Kr�<��ƠM��'2���=W��!������ku�X;u9ߠ �o�5:i����Ѭܢ"�)cSj�9p\#�z��o9�e��,�ވ::4T�*�$�'�������_�LhV�+��97>42�f)	uq�����`������2hP
AE������ӵX�9�\�`�ms�O'�To����.��K`�.֭�ov�B�5z���:47�����m��|�CRe�"-�G�4=8%L|h� )*�D�ۡ�r�Rhe-�"��"݁�	�333�����_���^�Ű6+�F� X�"���O���D�Ͼ��~i09`M�c��c���n)���4p���6i�u���KR���T��y^3u�AcڍB܅��s������C��{?}RO��O�s�h���P�e�W�As;'�U��T�n��Ƴ��<H'�it�t�;���X�;��t����Gտ���S���-Po:�w��\����I�o@3�9�ϟ�=�j�-�8+�)ڦyS�]�-��|dg�
v~1��|i`F�mJ��Fe)g��}� �4�~���L�X��5��x��-����XJ`���d�jO���b���&-D3P��I"~L��g4�vd]��o�(��Y�� nL~��'H*�;�������|��ZO����SÐ��*�E��u ���~�߇�
� �J(f���޵1I#���i��4w	�[7�:�ʬ��r��Խf2�q�!z|p��+"�Aޡ��'��Z]]��5���I��^}ceip(�����6r$�W�Y��C���i98=����i��~��Pcj���	��"�����b]��&�q+��b�G�;I�`�H��9֎�*��Z�E�����!�<�B]_�W��S�066vy~��i�_�6V�?�fИ�Zo��gǳa����(~� �RHP�����t*�\��$�t5��ѸKpX0�)�?��]֜[	�3L����7��|9�µ���_052�5���B&h�'�M��}η�N�b�Wśf�1j�f �C���Q),�DK��@	��g���^���M���*Ć;)p���v�u���P�,�\�s��^@��|�������k����###��'4F���G����~�Ih���b�ξ��2���n86��k]�(����=�N��m�7XgD�2{�^�*��-��<�}�W?��UaO�}���4T����ƿ�`X� ���l����KGڵ���&>��X�`;;a��\qE]�_oc/�A*�ŀ[	G����9(]#��w�V2p'�qP�;�h_�]�n�>\)<\W1[%�yҮ�hX���^#��Δ���A�{�;��p�v�-���֚h:��.����!�;0�*뤣����S�r������j&���V�w�^�	܊�U���\��@�o����܄,� �9�/5U��uu��v&��ָY\�t����W�#�l�a��gw��ЖR޳� ��+���l�h,|�7<	�Z�x�~~��O���G �k�~ɣ��AX/FjdEc�;�[>K������[���4+HC@�P)��Z���!��Y���*;�	�tPRw���[�|�����m��v�1>�F"5��0C�_g��2S���-��rK�☽ٔ�rIP��ל���9M�R p�@�n�ؿW�f��{�bF���Z���~:8���xI^����[�M w����!�W'�!���O琤��Ҽ-�s�3��S��|�.���
��g�NR�|;8�� ZOD��.��[�Ei��P:�k��=&,EͿ����5��(T����`����T�POiI�ͥ:��L#���� D`�V�&�+qde��U�1t52*w���� �E/�(�DO>�m�U� ��nS�°���R�6I�nC(��w��e��ޭ��3K�`�b���������}�0l��_��������t�jw�?�!���}C~���t�Ƙb��K���4�Ǻ���/:�3���vCq��'�.��7��p���m��+W59-�>0��æ�ˉ�r^�ƫ��䃶����I�P�����0�Έg���������f��?��{��j:z�o�[�.�V�#���aNat�4V����J��4�n��c�rg�Vl�� ?%�[�=(^�IƜ4� Wq������I,����[ 
���y� a�I��	���b�z׭f���+�CK�C���y���X��@�DvV���d�q�~{�4B#]"yټ�d���6�5\~3^�Ix�Y"2��i�0��GK6S�l�n4��:�E��L@P��d֬_�҃A3>j(�����1�}��İ�� �, �Z�~X��w'���hc4���(�{���_�U����\3���n�+aN�p�.��f��N�L���!g���.��3�\�5U��A�����deА��T.��~���D���͌���^,�����XY��f�����%�/R (*j��FW�Fs���`�=������l����3(#%`(tC�G)��\��lx"v?N_�V�9GP�X){rk�dq^fT��d���X>�c ��'X�0�Þ����fH5��e�3�H_��cT���R��ߓÌx�:��8����V#�����Eu��~��,��`��@0���n��[�^���m&�*l��~y֪�pp�������L<~��_�P?
xw��*�@nb�� 5-+��	x�\wO�+��g,�Rb���	
**���C�~���(�2����5��"c;��*����	C�#������`��P�	)_�Ic-��b�?���ک�j�ik� ;k�6�@kn4����Ϗa�,1�cb�1,���c��MZs�ʧU�ޜP4!^���w�Lԥ���q�}�ꕒ�/�[��0gDA!�p"{E�?��N�s2)�Q#��ɾ�}[��s[��ꩆ��id2�5QZ��,�,�����N�Th	�p����T�$`�Z��fs�e�P.�4�ɫ~���@/��nU����ۉL�E�se�F���7I��`,_���z��Uׂ�Rv�ZYQs���=�K�˄V�~�L�;��̊�����'CmY�"_C��w̆˷��	'�Qo���F���_����+,*��Q5�X5���Fw8�J�''&�� .켷�(�Q�	�,����9Ws;.W���1��K�9&5E�,�ј��}��{�wY���&~+���G�H!͹��>ju��+n�a4_�̄w�����s&�&��'��u�x�~���-���@0�[����Ɗ�5P:bJ�LfJD���d�n���T���N\r6�?z5fԾ����רg����W�P�0�/Ϙ"�u����x��v�M��Z$H���lBxtw�J�r���K�M��1��<�1�U855�B5�Ue�Q'�7��{c�~@�6��@f_M��;��nM�&i�[)JW~�2(��z�oO�����rB������ܢ�mB<�hѷs�o�?D�!�����DϪ3��Y
{Ҝ���������	��_C��۵(�[��$0�?	^��R�T�uj��>�M�?Do֭�oÍW���%;�?B�wxdY�lo�|qT3���5��]<�R�~��sq��,
��o]]��5H�W�'=��3�3�ڄ4h��.����TtQsmaw�N�/[�s�+�L콣���� E��R&g���I�?�NI�_m��OK�:Ύ����D�+�$�lHY�<<�菮�e '^�NO1��/V�0O"����yၫ {��٤R�د����<�K���~�t�A�W-�i�i�-e�F�t��ϑa+�Y��X�	H8ƟW���݇�B��ZG +�Y�8� 8ߪE�{�xn]�[+�����c!����ƙj+Ʊ½v��0F2j��9��q�y�F���ɣ8F��#&�[�)l)��\F'`�j�-==}�+���yCaa!g�]�l�3�\~�����#V��W��EEE���.�m�x�R���&�U���;�/�p(%7�%���ӺaY��RGH��K��m��K�4�芨M����O#�uz1�c��;3Ir�n�R�L5��rnr6,zwZ�����ɧ�s���ׄ��F,���mhh�aMԝ�-���fo4˲��U�{K�+,���[�B�fgg3�j�Ǚ��m�/��	�\�<<b;v��N�g��'�+%��"q+:�ӹ���L�Է���s�g;!j�]�s�C��������58Ty��}�_�j�Фo.��w�k%w�41�iM�V�n����զe]Fg��������#=!��"�]ᠡ��X�Z��/�.ۮ���m$��c������(Z
5_�Z��wu�}��ZQ�C��{�N�����r2�����P��fF~p(AES�'Jς`^���i!ƃ��?�%$r���+�R�� $%�����h��5���Ԭ+���P�w��=���C��t.���ּ�&6N�vUD�c>J0wʂ�M�Wg6}j,�f�|6�u
�͞:���"Ӱ�<�-�Nɯ;��N�%P<P��.�B��Z�-��Ѭ D�o����	��y��6��4�D��a�iC	�Ncp۝����J��8Дc��6���eV0D��؃�y�s�?�{����V|�h3�-���t�v���$��Ӝ���6��ey�����%���^�v�q��V��S޼y�֢ڰ��3o�i 
�@M��|�-�P���t*�����)����a\(:����NBb�H�)��w"DQ���s��jP��rwK��������%>�r��L��z0�F��6�y�|�Gz#�%hf�0�Y�FJ9�y��Ǖ�����z�ޮ�%<z�8��4��)��:�����-�Se(�w��r�ՓO]�D%�,�����mp�p�U{#�EE��Y'�}����3X�x�C-?�4M�s���᎗q�X�?*ydEZ�f���_, $��������E�*;׳�7��7�y���~~_�F����Sc����T�N ��� ����Ӿ>`�X���'������J��TU����&�������k���(����}�&9{�.�'PK   ���X�$&VAS }d /   images/f915906d-fb0f-4209-a242-05d71b94b060.png�PT_�/��� � �����A�9�d #9g%H�,9��0"9Ð$#�a�0C��3|߹瞺�^��[��U�]�k�{u��ի�ou/������S�caa)�Kkbaaoaa�cs��lq���N��XX���V���&@�t��w�r�t�|�b�����i�`��������Uڞ(�c,�W�^�;K��i<�B�Ր|b'%B�Q{]I�s�iJ�嫃\�oa���ͿVA^>@�����'O��U�Ka�t�z�0�5a�-�Zw�!Ȱ�^�~%��e%e��������9rֺ�m���6?`�/G</��6��>���%���~���#�y��7���%�_��%�L�U�<�Km�.P��&8&r+�ͼ�_��~d�N���a�c��v������ #vv���U��3�y����>�X��p�>V�6- Cr�O�ˁFo�/���n�*��v�v2Z�ny���3����hՐ����G�w>F�4w�bL$_%l���d��5��E���%�Ln��P�8����ܒO�]�&�m2�&�����'r�c[�����`������x���t��GX}i<�J�!��Z�?�>w�gÝ"翙zv�~�\_��^�3w��,![s@����-Fa	�_}1-�^��1j�ﻝ����}����-/,����jֹ�s��㲎��x\_���^P�5%+F�e��{C�������R�]=�=���N[:��8��mF�UY �	����P�9��R�&��f�.���Se➂\C��xn��>���٫H3h"7�}��p����6G����?
��f8���\&��ɿ�����U⫬ed�=�u��t(y ���a���L��n�v׭�^a䨑�6��� 4ت! ��W�ڝF��+g#��O�l��&��8�yk!u�W�]<�QF�r���@d:I���"h�n2mֵo ಑��~Fߑ�E�9~��b1^��Y��D�	gng@��[��$��/.������a��\�nW�u�w�>�b�?aۍ��-��1Iw�vs�A�,;�P�s��L�Y���o	xF$\KbwZBB��^&��6m٬)5��>�p��՜�T���N3�G�=��0�A��{����;g"��>��c������X�]�e
Z=ϋM?��?&�T�W	��3��!J���&�M����4�2��!j�k{+�B5N��},z�J~��/���e�V�t�X=�Y:� �\b�~-��2�������l���Q����̷Q�狨�����3��}���=G"���b2C$�)�k�� PH�X��4.�*.:�j�)����P�u_�Lißԡ�PԆ����cϑQ����V���n[�0�gt�r��&
��W��%����B���J������򙎶�\V��{��s��K���t�οs��2c��c�*����%��'b`����'�b�$��O�]�AeS>�i�l��=f���Ɖf��(l�̌m��;�_���D�q�I�߻�q��
�)�w��N[@v.�i�6;��J��k-�TnLd��V�<bҀ��#/�\�L�|d`V{��e���]����3~Ÿ�_O�0�j�uJ���܈j�gP��Bt.�n/�h���ƌF�����Y;���J�x��դ^����*�{�Q5�*ݚ��*�q�Q�v�J(G�D���ذKL;#f�Ni�N��s�? Y���2A��h�&��,�4��ֈ�ky�{�XqM�0��C���F-n�0��Q�#y�Dn3���x���N$��6X��1l��A��@��%GI�p��b����p�Ձ/��Q�)�
��͔k��쬇�O�삂ȋ�����4��
=�+���%�I�m����%wL	A�r�L�~c��h ����ѯ(UH�ců�h���=���v�TV7pE��Z�w��n?����&h���L��"�ƛ�l�������5�	gWa;�&��	gJ5N���ݶ�� ��5uʱ�}��lᙬ�٢5��Ǎs����8���\]$�ۣf�I.��'�����ƺ�*'������K�3����Dmf����51H[�f�6R��T�z����T��kP�R����U Ѕ�+U��K������uCGp��y�-����QG;�5�#��WO1n�b�Ą�mE��޶r��ά ̂���d�ap����Ӓ��j��)�}k n�Ep��%���K�J��Ք�;[�_�#uI`+��6]�(|Z<�\g�y�˧뒹a��;��mJ>N�Xν�S�kHlQ �$���``��l���Lb�D��L��L��(@�~�j~��*1,������arS�Y%����4i�*1w�q����7(v�$3Nd&\yr	�����r�����1[)�u0^?�Z�ġ�&=)� �ܴo�hy�th����J�����D#��ck�U�vq� �IvF��G��8> N�c���O�CWc�(T����㫑��-������o]y��:�f��Y��O��<w?d�}�	�	���sa�C������+!�Vf���R�[y��qF�g�� �+@ZC�+�;o`��2Ua[��2r��Z�:�Z�<���9 	p|�-�����8�_�/C��:LZ���T-v 
f����f���IY^�P�,���#`Mø����%^Ed�Ty6�@�{e&(	Q$��V��z42?b�D�N(��ƍ�V�I̔�[�pҌg�m�V�=K�F۬&�^_�T���9}�?Q r�?�y'��>�qW;��-`ǲ�=>��e\�������=(�'{�+��h�ꀝ�r�=*B��ȧ���{y �ENЛN%�$����+�&����@~�q�F�-$�xhd�S-�L����L
����+/�2u�?p���H�Uo�\�|E� �Qm��ȑ��fZ�l�eЁ��,Z��w\�웭�\k(�8���5(T�jd��u��Im%e�����2����=rsI۫�U�������9İ�$Kl#B�+�wn"�Fvx���TC�PU������	$|b���|rЊ���c�e� P��ܢ�>�x\�ì�^�+ Ϙ"��b���V�/�Kl��7\�p)R�����Onkŉ�G\��3):�j���7��J��\��/-�^Ƈߎ��u���N@���]D����l��r��X\�T,�Xj�QE���M*f�>/������_!��_�U����Zm��͊�WԹ�/��b���F/�s�ds)�fL��|���\>=#���Q!�<�=���>���h`bM×g�f�jf���,&��~��c�=+���Ą>�6.�h�c>�&���$8#���X~���+p���z�Py�g�1�\���|j�'Ծg��� ?�Nx�'��	.���1N�Ax���d��a��6�)�u�d�?^�x\�V҉ӄ5�{�,ik�=r�����չ��m�}Dq t�*�W4�Al����κ��Dں��k�2qľU%��6φ-��yѓL����ý�Ck�P�R�HC=c�TP���̣-lT�
�Òת�5oe��N�X7NJVI�o��F� X�n�%�@��R���s4p�S��H��1�)���> -H��W���2��j��u�{#�&����;�����v���5)%�s;�|�*����=�v�d�ts_���G�ux��Ү��qLw,��U��Yt��%�VX����"����������Va���6��adߵwN?#���\.��Z�
H��4�T޺��=I�=�yu5aڣYxu.0�u��p7vre0����B�!�2@kuc[��F������fނ�����D+?�o"�b��PjX��jG�hw���z���i������Zl�L��l�ᰢ/A�M����F��!|}\�7�s�{���.5�6U�iE��߄L�����-�g��3���j�X=$V�Gy�[��Q>�!�ӟ7x��}h��A�u���9�2���b�l������?�����wUGFņ����Tb%Z�u����C�s�(|�s/z0o�5b�|+h�d�s4��0U&ֿ�L���:��Ǆ;�b���we.��W�M�S8~�g�j3��x���;�����Xdz7���f~M��*�ōF�f��'`o��^�H��	�F�py`�\�o�<���IG�Lc���(46^~���n>�.��E�[!1�A'�ji�ɢ1��V��NNJ���C!�� VpMvI~D����H���=�ӨCx)�ɠSTe����4T���t���]ߚ�z�3L(,ml���fZUr,�HA=;_t�68o�?q�l��I0`�9)�Lk�8[������ "t�wr��~qcK���p<�P�������O>)��"�Ў6Ӟ�9H�*tS𚯵�ڔ�Ԉ�Vn��n[�B������a|���`n��.y�|rU3�����̩��������t�w?���h�ܮ>�����#f�yJ���&ʤ�������a�M�1�
����x1,�`ӒAY�^u��ͥU�Ԧ�:P�.�d�b˃�l���tи�m7c;�AB]a1�;�a	��
6	Q�6�C�E Z:_Ʌ COF��b�c��gk�r�Ǐ��L	dU�O�E]��!-j(^��W!+����7rΌ����?���Z��a���icMޣ������S�\E�M$�M �bO|�nVa��� �Y_����l"����D�D��dD7�቗�@�Sǚv p���������P����6i���}� "E�騳�l~�k��W���d/�$�Y|z&�f��������R�-v��-7t��Z��|mQ�_��u�>%�4�u�C>=#d�;���CZ��WW�'KJ�<�J�gQn\=-�c�
 E)�H�5ym0�p���`�&Dm�zX_�|��y�1iL��]�B��U6��v:h�lk2�#��L3�v5gXrv����?s��k���"R,���f���2�2����#�p�5�LZX��=��H��e[лR5;b��Ig#����#݇��3Q ��;k~�s��� c�Ap�%>���j���nƕ,�l�J.?�[�t.�I����֦4�~T`��	�Ewo3'-���� r�;����� �Ze@���S@a{< ��� ȳ1�#r(U���[X4k�"J�D��$>qDq����9�e�K��ՠ�M���$E������.����G>e�@S���Ji�sl@怮�k�z��h2Ť4G~��5���� �7���z@���͑1�~��0M�	8NԷC;R��	��1�Q�" �:m~u{GWF���:��枯�0�j���8�\S�����(W��l��R�!X��f���[����t���i�th�<��}C:�?X�%G�z�<^S��	�J!kH8i斳�s�n?E�&V^�XN��zi�i�Vؤ�M��}���u���!�>GVJW� á1����uH��Ew� �he�:2h��(K�OJ=�a?�]f�_�k�Kw�7d'�lS陹A���٤�����@c�����$f�9HM^�1Q��1	�1��!�\�5���6�ن��F��O1J���|��S��3���#u��/	���C�=;ށ�~�j�D-��%G�M�JW���-����W�*�=P��#���N���I��2)	�Z�x�]���#\�/��dbZ �����o�/n�e�S�Gn�I��g���n�At����Ԕ�w�BX�_��
"���W���U�!��]�,á�n���u����o����z��/��蚸�m|ϐ234��k|���4�$%��Y�ȮFӂ������(��Kff�tB\c��R!5��q�-��~;�'����鐰*��>��~,����E�H���y��,��r�$KTT��������ؒ����bB�͗�����;���Cأ��mm���kwc��N"�F�i�g�KM��Pf��)W�f�򠖲!"��yw�K�&p)�_N��Ѥ������?W��`){b��Ƃ4������LW��(Q�������`N�ŝxm���v�!��{�Qt�l6v�!= �Gޖˌb�n�tſsu�d���ꮠ���Q�/a�+��={�s<�T���	ș�6�  Jh�L+-�.qOG��������w3��֠��iP�'������ �y�0T��ڱe���l)~����g��w��cc��ȶZ𕖲�����-Ty��b������&*
�Ќ:�r%�f����>Q���V�7V#�2��6]eA9M�U7`�QVOxG^ -�􎹧8S�"|�DI�hȕ��ï��������I�vZ(�f+��¤$�3�9�>k��:+@���<�*�P	�doZWf*q���l
	=9��W�+�_q�6��#@�@����(w��h�����ۅ�x��͛hU����z��/�+>�kce��;*�P��\�i��/'�K)>����d*+�Y2�([ʃ�_<��)K�֬dq�����	��I�}'��=%!X8QSS�27�^�U��=�X��5�{�-i�w
�^�xA#��@��g�c���r̾M37iͶ�M�>'�*J����(�k�<YE@�"SzZ듵rP�RcИ��b�r�{�Wb��D}��Wg�J���F!�VF�x�� �;����V�v��wfػ�|�sW�@��B�`ƛ}|�K�r4�RȨ)��UI���(���������GC��9)**�A�%��w�#2��_`���w����9z���/�{;҃S^ptFG�@�@�2�Z�����Y0��dU׳Q���+i֜Q>�Co��K�?�({�jҗ����U8�D��9���FzϴG��3ɢ�Z�N!�
W��.54�<�I�`�E����{[�
&�&��ܻ�/'�ݬk�q�%�Q�!	�7��*KJdI�m��6z�@�y�I�f��)R8 ����įzܐBsCY:����n,'}�5?�h�_w�H4�/�9=�]��CG�M�nt@��)/��r~����͸M��ĴK뮁V^ ����Z&�(�.�mh�,}A����-�+¯�e$"6sL���%��s�«W�2(�t+��n�v
�����W�uI?�f�pb9���O(�C3�(�m�e
��jl���M�e|���ߛ��X.���a_�\Ӓ@��"d���G��oI�f��Si�ּ�SPFY�+m&"��ak]�����T
�]�p�ׂ>��g��
�y����a�ejat�S�'��Ή浿�� է��w����=�ȏ+9��㢊�o��-�<����hl\_qStz�-�Fԯ]�,� �F1�qn�4���%ci�f�������F.�<���JT��NŮ��k��,�iE�����[���}u��Ϫ}6��1k�s����s���e����i�ÚN��CXp��HN㐽��d�U�a��И�1�$}�XD,2�
���p�4�
�@<�����m� (����T��P�VB��� �N��n��V-{�x�I���r����I1��t:p=]!&V��2!p�='���g�i���Y����v����1��iv�"���|N�u��V������[@�u;p�����VP<{��d�@�� ���*qQ�(9tݎ��PϺԽ�VVu(+��ǜقtB��4�c������=�zY����Uu%�qR-��N�Y���yX�P��"�{G6�C*�ס�Ֆ�~97�c�a
Z
]Ӟ��jZ�P���*�����I)6��7��`��T~�T�2����K�$b\Q����Nm� ,� ���;٬�,��a`}1B�<��5ˎ	-��E��	���~1_=ty2F�lj̢W�&��W@�-�Ӥ���xmt+6���y�(��2[z�œ�C�ZLaU"�/�'�je�D"9���b��m6�V��h�����m�o�RI���� ���k���?Sm���ъ��� T@A���� ��%�e���>ɛI?B+�JVI_~���aƕ��z�F֢��������?��B݀UY�Jhs�[�ۗno���7�ҭ�dP�!������9oL0mƨVtWe�럪����&?&�&�?Y�&J	;C�
�?��J{)�`B�#h��LÈ�6�S~L.}A�7nU��W�klf�)�]oJ�
�#]��Ų ({�?�w��1y�b7�	�7:b��Q2XHN��YԿ@Ar ��"^ �k�@H��\@g���?=cX�>���k!�5�8�@(i�' x~��2O_h�������Ԁ91/)g��{�<�l� $�K4�Pǧ3�(�s`�`߽AnH���D"���T�0��\}�\� �KH忛8�˽R�.��0�i�8��=��l��T�[��!M%^r��KSE:�e�������!
 X�����x� �&$����{r"�a�h[���2Q*���7�����1{��Z
[�:4(8��a�.�ihR��P�һ�d��p�?�կP[8=A�j�X<g��*�NV��{F��<�L��?�7sz�=˲�F۔���x;'^����D�C������f�vV�� �'���j��s �P?��	} gP'����'
�T"U_Õ�����t���)���r>��k���o���]�=6�S%��4�d����Ĺ!�"�����HrŹ����ۊ�Ŋ���z��&�d��w0���gI�j�( �1g����[�h��4�8N�͆^���޸�A�Fτa��~��[	�Y)�Ex닺+'��l��v^��D����#��V�ɳʠ���/1��f�]���m��R��B��(� 5�Z6C����aM�[9a������G�176�qW�t��7I����JaD@� �I�e�z[��LO_:w("��J���bJ����V��2�^�|�C��ߔ��Ň{�՚ƙ+�����EMʝ1�,J����ʌ����,:���mi?}V�D������&�pЬo$%�;���B��k�8պ�gG-�C��7ܯ�B/��H��C��(�i�gQ�9��/�ϠZ�Ǵ|�Q����������Ґ���%��Y�l
��b�]Y�{0y,ٙz��h�*toǈ%�`�JX���TqE���)�Ҕ���߲�I��.�{�>�9�7~?���V����i���^�l;�M��(��ة�ft��.S$X��M�b�̝1�^K�db�J#���J��/�wƸ3�$�O9.��͐���f�d?,�3c��N��ZuӜ�/�V��+��ή����t53�oq�]�~Ӷ2��@Y�N+�W�]��6�5���UE�J�U�Jq�����[�>��t�Y�Ѓy��0�ei�H�^4�ӊ���J&.������_\���m��^��@TD)q�nM^���N�R�W���A��Ӆ��ˡ\��yz��h�%"��� ��ǵ�Ac���v�3��y��Nx�-�T��_fс�w����<�,�Y�R$L�|�Q��[�2��A��#�;���G����|ٳ9�0��gԯuK�%M+���8	�X�_�hLzWm8$N��V$�Y/��|��w4�Np)�~Q����%(�^���܅>�{Vr���%������iL�0��]?�3�L���W����p���!u�{�w�-��I5����&��YT����F��
G�3�8�|�,`�r���G�r�����V��m<2�{*��X�p���g�P�a�f��w�5�4k�~tH�,@��@R􇿹m	8�2]n\|^Fl��޻�	@fv�LO����Q���W�y�X���Lg>���~F�Ô�WJ��и(x�� Xi񿜒��=8�|�@�]Q>N6O�
S�����GM���a�'����"dL�\��?�֝--����|�]���ԅ����m��Y�2m���=��P�r�OLǾ4�vQȊ�y#R��~����@M��@��g�C�1d�9���9kq�6������L��O���yS�5A���6>���@��G�5㽩�������;g^���c�c�u�8�av�8�|&ze㑀�ې����[�Bo����r�q���}V)��j*pN��Lx}���|�+�����n:C�ϓ��I�tF�Bh��ְ΍�le�V(�?h���3^�coʍ7�ؗ:V��eI+/����@[�����'N�8X{�C�SB�������������}9�`��?,>zs8���'FAus�hvE���ÎC���sn�-&��R:��G3�I�%��h玿g��nV<�ڮ�E�+��&۴ZMva��~p�n����ĺֿjR�E�1ʹ0v/X�ӷq��ح�L�5�[�l64L~�3fچ�}K~�����%�|	��?b�aHe�R����}t �B��[H^{����Ӏ�!zH���t{��i�A��s��yo�[�7�s�����x�Z�^���0� Z�&��R�-���䂌�W���ͷ��mg?�h�#���=�C�{�Ƒ������:�/�*��N�#7�I]��I���9�*�X�a��AT~5�*� �㿵���<�%�q����Q$\[>�Ê�
M����e�ݮ/�~"�'
'9h����Xd�Px�L�-}�p�����zj�� �\|�o�V�7d��>c3y���9��S
-�Fx�*��t��>)hyQlt�s}`S״��O9ΐZd|ѵajX(��(�C~*?���{*kZv���9��~�~k��U�����/���`�b�ې0��G����/�K_@d�CT��GS�B���%ƫ�/��^>G!�K�>��1��w���E��P�C�2:5w�V�{?N�������.d~E����ljY\9z`Ԥl�U�of�`n������u� ���^��fЩyl���k^�\��,H����ջ~��[M����	��+��[��:BP���[5����wuI�vc]҄�E��M�C�g=���?��R��3H���L��2u?�3'u����A�ep�	*n3�CLwI�v3t�/��h�Q�vM
q�J��yT�,�)8E^,�p��/��)��7����������ՙIBw�eb��'̼U�RC�ӆe�˼4�р ��l�
)�h�\��)���t
�41a������!�E'�(°ҟ(-u���U��%���i^�j.�����Hz�̍呂:YgD��?��̚��7�+Ϻ�9=��)���V�u`hx�G��Wb����{=�'K[3��_�� �������=z78ީ����Π���V$�ŻE?�Q"�U��?�N��k��WC�l�$eR��o�	���|�@BYW.^��I+��tK�nB��a�G�%#�=3�g��8��CF�*v�����u�P�ČE�9̄b']U�䄝��#3���u�gDJ�s[�ĺ
Z�|����[*E����f��+�������Y22��ƥ�yX�$�P�%m�i��N{���ғ!�*�����Ͱ�����݊�����P-h����Fidg�ݿ�>���F�Ϥ�6X�FNES��Ig��bW0�v ���𶢁�������Q��{6 �,.$Z5�͏5��k��NS}��1w�s���M֨g'B��!�vs��ݏ�
��.�����q���@.�N�j`W���t|5�*��yQ�����~��@?i>��^�lTd�}��6��Ҹ%��j��ϯ�~|淽���0�11��M),���r�����bT�()	���Rm�y+��Ӭ�������Sg6 \4�&�Fs��}�,I��a��՝�vs�;/��Ϝ�d(�>���_�뢁����m���')��@���fN���#�[
�G���b�M��NH&la`W_G�@%����<<_ro��"ˇ��L2xF�\O� ��﭂��z�S�[�_�]�K��c�����$�]��O�(֌���8�]=�����e؅���K�ȷօɯk4t�͜}x�d��:���u��������6v(S����V��M������ù��'�mp����f+9Έ� ;�ee�!D��ffUּ��22��F������������zk���(j-���ʞ�/��Zͅ&������J��M�CУ��jmw�KK�y��X�����h��������f�Y�{{�::��EEt�����-�EǻE|v3͜!.$w���@r��t��I-Dffflg+M��<������������*�h�U{���k}��4_gCEM�y�D�����u����i�@G�5�5-�8���j<��C��|�[�Xd|=:�c�1���Ղ2�r�]N��7�n��>�_����4С�����#G���ֶ��~턾<�JK������r?�4~{H�� �p�EHkkk����k5�k�������+r���
�XO[=v~�DQ$��1�����!���Km�v]!D��9Ӈ痀�f tT��[/��[��wf�;.�s5�����jYYv�����U����l���:dS#fM�E
T-��RI@`+�q�Ĭ�:��a�J謀P �B���� ܂�jUv�S�ɣ�e��C��>�%.�WZV��C�αk�`H����u4�X�U�4"�:���u�W-jj�fKM4�1�t��ΐ�(�9R%f���(����c�g|��9����}wϲr���]�:<-��zEU����])VK�Ik ��<�`�[3;��׍�lqcJ׷.���^�yW���ol�,H�� ���3YDG`Fր��UTj�d����An��}�9ꢸn�V�"H^E�~��k̕��@�$���QK����Ş��CO����Mv>j��R����Gww��{��tta��D@Is̀�b�@U����Q�HH�
���fJ��/�=��4�H���J��y���ʋ@���o�Vu{�]�gYi9�Ʌno�/Ɗ�&�+�-��#�he�s�NtO���,���#��Qﳞ�p\,	�A4^��u�g�G��Bz{>Q.�(�"��ӕP��i��#|5c��8|�0e��M Z���w��T�!\:�x�г�]��a�tvƈB�5n�R)�Y���1T]��r�������Пy���6���:	�	k����������-��E��iu�t?{�W�F8�2PE�����,�iz��!��4�h�����:�֋����D�WF��t���������!r�| #Y>��Zl�wPD�ɢ��F�i�s/�	��܎C�*k讃i�Q�JӲd����\`����V`��kk��#AW�EEV{X&2��ߎ�����J�Q��(�\	"�(0�|�"1_v�ٜ���0�������j0��H:Q���G�D.2��I��t�:+�HO�;g�"K��sRóp�I��@�[j���Z���NO�@�7�
�L�	�ȍ�H�����.��\M�5�"� ����>HJ�����l��Q�RJ�����)��=�Ԓ��Â���.�$[ޫ�����s��,������9�b�}�a��|�9����O�� �GK�`�(��W�|�{��:���.�#�c��v�Ň7�֫�\�/���ږi-�H�[���5|�K��N���ƪ�^����9��Y���mU&kl�=�뜙���~{�r{��itpn�w����	C`tW�3SS	�RN�pP�Ѷ���TuoJ�LjZ��ZҨm�Mp����Я���Y��eÇ��=ۙ4���R325�y���QJXD��$����Wm��q:76,.\:V]�	�����PɮRw�bN�B�R�n%7	����&!��:<��=��c�a�������>c�&��2�I��������=�=Gb��(@�̰�<+
��]����<�J}�K��5�S����~��7�O߱�IVU�����2�|���e�\��;bOظ�n
��
�-q)��:s ���^�7�q�p������E&6���.�*��xJ�	vvs�a= i���s�Z�S��j�f}�?�S���K�L�;����et�g.IV�C���6�
��2~��r�_"�lՇ(��6���u%3���Q��l����P��q�_n�]Z�B�w�+ C����Q�qE"Lˆ� �V|��'�����D�����w~���D��a w�y6x�L�NM�a��J�jn)w�[������cN�M��51s��S�h�9 ��z0��o"-�_I,J�!��@����c�����]X�i������� sy�LJ��w�f���3�z���O�]��b��r}�R71,���%O/m�+���Œ�*��p��!�5��������^�ĹgE��'�B���I[[cC���_otZ���N�����3{�|0c���o�ϴ�̟�#Eŉ�y\��Hr�����000�A5bˤ���F&X	���i�m~�|[3o�\8[ov�r��5O̫QZ�$�-	^��[1��a��	T^�P8f��>	����2�M�۲�^���r��Y_��XD�.ya��2q��L���]����U=�^�P��5Bd��X�a��.f��,ƞf�B{�׮h�D������Q)���_3����g]�tI��ZVt�et�����%zd������R�Ԟ;��o.�m� �S%T@f3���̎~���_�V���#�hx�z���ޖ���~�;[��{�ڻz�
�yk$���������GJ~P�)z���n%��W� ��qe@_����%�
���3���p`/���o���5���q��Y"�R�t��l�j��w�p/�քSP��b���	W����wf���q<�x���m�IU}�ƑoU|������:H��ҏ���2���9���ŭX�ۨ��.��D��N��N�Ғ��G�Yy��8]B7su_0r�C�3�'p�z6
�����/�O��Z
�n<B� 0"? 7���z��1�\���%��1Ά�\�lO~a?�W+��r����]��6�����^K��v/`,�&)��~������~|1C��̼:T�Fl�Qr�Û����j����V=0{T����Ȃ���� ��Q�E�����A˻�N��t2E�g���?O�����I��oz8VZl#���]��:Yl������C���>M9ʂ�::#��5��m8]�l!7V�w�m=�t�aJo*-'z|�6�����!��	AhQ��H`���cO��QJKK��ٍ����������7�Z"&��ߍ�yh|U�Yr��.���r�ӯ]��#���x�|��޽{4��M~�%(--}��]u�G��;a��d�>N�~�� kbbR��xG��K�Wlʖ�?5P�]�IK����Ib_�FRFߛ���;�v-y������r���j��f�W�_�����K\��fff��г��ٚ�޵�G/��M%�������}o����i�Z�IVzz������Z
^��dլR����_5Y ���`F��S�@3i���;s�E��ܣ�
�}��f3���~P�kkOm�++)u��|�����We�^*�Y`\�U���}�OP4�]����W�/��%�I����;��1�c8]\]�W��ؠ!Du�ll�Sp��}8����$��̃XL��!���F��U2��o��D2�Y�5���RL�үܕ�r����=n�3����{�}o��叏4��q�[m����a)<Vnͦ��amK�n´���ʪ:B�:P�З�m��oZ�l���~p]�L�/��-��8�%qx]��}��ߡ�e*TI	�����Z�	%3��X����3�$&,���b7sW%M����������e��1"�� __���ѯZ�]\���:�׼�adaY����|u}?�}�Bă}mm�b��~�m��!�8�0��}��� 凕�1y�ʲ鯩��Ŀ�p���>�|΋(W듖��������\\\�!.���N w��&o�F|Ğt�fx��qv]_�G����"`|00w8Z�ͪ��{w�7��|�S�۹��*y�c�݆��A��w��g&���8�v3��G����N�ڲ��✖�g�F|�5�%3jrЪ�������R����ᖴt��XA��^����$F�p�H_�~�����h``�n���+Q���Z)����o-AG�<�u�*��,õ�<V�pcD_Tv�X����ᝓjQ�GXy[�EEuJ�}���Hz����{���������	/���2 ���E�2���R��Cv�Nl�W���zv~�iF�	y��Y��n׏�E����LP����]IFGcI�]��za���H��yL���|��"����׋�+ ��i0��Ù`�aEo��Q�^`�'7�؄���'tLIɐ���-z��>X��J�Fu�]��.9u���Vᩩ��y�fq@ �C���<��~��򜅥�T��n��)�>ڦ��1 
�e��~AC[ۭ����O��J�g�k�;B�����G��:.���}�s�o{#a��gg8��C\5����zMS��������C�x���}��K34�MXykk��}s�v$��\������rB�22]��Ɯ�?F�}����G
qQ쮐��]��t��\\}m�E[�c|�㏁u�+o��r��(+�j��}�9�i� Qj��4�>��zk���$�u=Υ����o��U�]K��황X���|J#�3e��DpzKR���b��G����o����e�����?PE�^�c�*�x��G���i�n{[X0�]�w}yҌ�.sᛕ�0r����=gc;�N��;μ �эG��&~V/5�A�etqq�9���������)�d���O��/J��b�����i�\���������3����ᱠ�np���ݛ �����ʊ���c_������,n4�U5�3�k{���0%���u|�2�'�xÄ�/���������˶�P�NsXh�nf��GG���gMb�M}�á�{������C&S�M���������)q��-E�x�x�un���)�ʔ��}bxI4�����x2[o�<^0O� Pqz�������l,�s�˼099��v滶1��'��	9=�Z�G�ͪ�y/�}	���'�_x�����Bs	>q�mO
��L۾��YNr~�y�3:����$������Y��,�Ot	5l�	O 8�;53�[Z��^��������{��i�i�C��;�����.ARB@iiI���j��������ݏ�p-���������}�Y�� �@t�
��T;���6�:�\�c-��еaU��+>��d]��c����x�1�%*Q��.93T�n�S�-�Z�f~k�d�5�l���0֓y塎���:���>xmW�DJ�k�8?�� ��x*uKiY���-J.�����y�pQ$O�.�{�(z��8�1�ʁ�JM�IMs�O<��B�&8�Dy �R���᡺�6�׾��)��E�M��vU�+ZƊ�Ѐ�G
i>d�_k7���+��ը%��Ë��OӬ��א1���?C;L��w�+;�_k����>-���ZrC��#7��(��w{Ey�Α���:���x�gU����KL��U���5�'<���%Ixg܆���-���\�*�,G<�>��φk���̗�4ҙ�y���}�+P:�:hWwF({n ��P�!�!���E��?�n��=���x�y=�*�a����~��ҝ���[�wh9��v�6A]��:� !�|7�\<��y�QL�R2�˺ 8����Gy����-o��=�&ӚE5��ţ�s��[`9-��+�(�z�sr� Kt8;;3��wa�r�W��E>��ҮN_)��$�h &z;�FC֎���4@��U�����	y�kB�?t����cU���K�Gx8���Э�|�<Yj���s�6O����X>�lrrs㲵�5���7`RZY�&`���*\�	�\���e��Cc(��9��J���isG=::�ŀ�ORہ݆���Oh'����$^")���U��BZ�(�k1-j���z2��Vp�S���*�ݷ��\�~�I<�V---X.f��b�@�]���v
[��ns�7�1Ο�E�E���vU�����L��˽I�y���+b��gD��rm����
��Y.�	�hO�&h��@���������Yj�8��O3�EɊ��:k)L$��g���}Ȅ��,.-�27���~A��
H���J��b��u��@*��&B,j(x�@ wf(&������330�Kʲ�S��[�iN)�]�ƾgz(L�SvR�8����C"N��,&Po?a�)nS�}d��P)P���-�����W�����X� ��,�mCw�C����xxV	�^�IR�VnZ�Ӻ^�_�
9�r�oe���<J7�S�@_�~}8=_0�RG$�+�ta�\+��S4 ��E� ���k2*�;����e�1�3�Idw��AFb�*@*uuu������|E*�v X�S�_~TV��W�����"��o؞7��Y���@�љ|�jjT�?~��/�)��O�? ������e�Dqtfwww�7
/�$"�X���:�%RX�Ϲ�r������ߨ�o.�V�����2$:`Fl�J�n�$�k��_��&��Ȅ�4���f�fiߩ(}��֍�WcN,�bz �9�_�*:�h-�dp�w8�9g,kllq�_N�3�ck��/�U"L��V� h�p3�����Љ�l^?�!�\�1"#:��Zf�������P')�Џ\�pj�Ƭ>F����o�N��!�wP�ڽ=X���bY|Z��~�bnRPX��7��B(S�~�v��o{Lz|d�Ӌ�F�#Ugs_H�#V\̭P�J�:�@>�s��
F4��# ��Sޥ�hi}��.���b�
R5!��Ԓf��H3�����T.븭C^��H�� �I?k������ ��+,^�Ü�M�<j�p�u�}t@&d�Y@�#|��Rs��l��'�:dM�����,D��ɥm4���}Kyee/��H�<)���b�H�`p���g�E�:�3ps+D��ƕ��g�������nA���A6�b~�;̓�3���0�|��e�)���]���� �tc�99M8�U:�ʧ*��b��ZRQ���> �kY��E�b�����咶���5���T^^��ۦ��٪�	A	���4E@*f�߇"��0��WϤ�c�fr��������(����y�qe�B����F������o_���p���w��x
<\�DP���R&�Q����0!T���\��]��C��p;�Iw��A�Ug��c�����ݪ��o1ė,Y��pX{�D1=ȱ��Q���b
k��ϩ5?t�ӳ����e���7���D��{�KF~n5�8������r"s#+;�H;�O���Nÿ؅cj�<��+�~贂BVK_���҇
����\Vj�t����Z�iP���U�!h�F=J2����� ��M��� y��o�/qrr�[�-�1��^���*�W[���(��?r�3)��X��f'^�d�`$e�AJ\�_K� �A��������"sF_�r�Drss-k����oP���5h���	�#-���K�	z�����e�E=~���i^��nBy+��yx;�1>[���6D�4L�c/�������PB��0����_iy-��Z������{)u�����c	]߷�+ќZ������+�-�ɀn^v���I��k�����3ӵ�;dY �CHAq�y�/n����6�l~�����FF��Q���o�X��?L��;���w�%m�d�Or2��t7�j���"�������CLV ����ПB�g}DBME��3���L�++��h�IB� ��y���/�a���n��Mm�����A��c�%��~�����Ȃ=��ىM��^��~�
E�feU��ɛ��4"�1�\�]I\�*R�ջl�TR"<\N��y1�-h|q�}���x/=3�a䑐�j̀#?�����0�}9a.c�UC���x���c����d���G�B7���� ��=�J��)�@B��d���v6�\y@Y:��c�Ob�U����\o$��,�R�s'�00?�Xc�,h�pcc��nN�a��	����M@?�%��nϯm_^�c��΁�����c����y(9�v�gK��4�~�,z��3�V�xL�g�4Ɗ,���[�/լ����8ӆj�*q���t�t�,a���b�s�H��~-#��$BV����3 ���X�F���&��������%e���-��Λ*))9��-u94l�7�&fveszU���$�|+�xsj��Ǐ���B�t�����B �{�D�B4s6$�Kg����o��6��{F�G�"q��p�8��)�dF����5�Ym]��Ӕ��=a�r����w�q@u���T.($�i"q�Dl6��������M�=�z�z�D�w�8[2~��?(�����-
ő�`&v��x��E!�rӷ�$��z�ϗ��44_|M�I	E����C'�W��3d�uF
��4�8��|g@h�f��ܯ�$A dm�J4A5�>���;;���P�0������'�z���"�T�)%���&��ױCq\�bM����{/����@H�S)�3'�D�T��5����ɾ��l��ڟ.��'�)�)������J4Y�zĽ`$�/�XI*Xn5x���~���>̐�E� 7�c�8:�K}&�(FZF�-{u�ֵJsHkKA�gt���y� ���~ԉ��o�,A���TFZz��u�lG�#����x���3Ϳ$|-�����B�+)}k

�;q���fx��[�?ޫ��O�~�c�KuvD��K�>dK����8��%]k�/��4�I�K��]��Tl��ޑ��*e�*�v��^Y�9 {4��s6��~����l+(v<Z�����n,��{`B��{\�b���4��,��jI���fz�6;3ޒ���eِ��g�:�o��FP+��BW���$�!u�O$@6U��"e��@;5\Z�O�Un��ȸN���v�M������(UlYؤM���HTm-��uH���߼?z�P�>��r22E�ou�ۗ����d��ihh, ��b��F�$<�<�qd�WZ��˺?��ǐ�.��^�<lRA}22GF,�hs>�Ւ�VQ�k�J /���YZ�f"=*����H͋U��c-s�;��E��]K���ֲ�T"�3��tIXT��:e��U���WnM�-��lѴ�{�ê�5&�X�f�FO~ӠU[�W�tw�[f�F:o�J�K��z��b�[]͉Fk�"LU�njz����q6!��j�ÄջD����n}�f����l{��t�q�z��qJ��uXK�А�殯�5�±��TD��׮��FB�l,i�֖E��	\�+-�t�^����<;�ΜO�o�u~O�iķ'|μ�]�(�Rc��θц=��'ח�1+1�Ĳ\��Vuh�6�v��r4�a>�Bs_��B�]֧۶�ۆ�驫��B���N�I��G�0�b�kU�:�+"�Vo������y�ؠ���f%�P����l�R}""�M �^�e[���/�UX����VGX2�5���W���n���v���p&��SȪE�����k�H�;���6�@����;i#��x�Fw���2�.���K��o�ڻ����e�6�5�+�����S�-]֪Zd������3�@�������:�Bn��B�r��y�G�F�ݽʩ���^hdI|.��jTQR���tbJ�]�CcJ:���E����C�����VV�Nk�F�m��Y�y��a�@���B��T��������Y/�e\)�}��d���ѢBs����'n��Y��D?�������E�S5�u[��׍�r�!^j����)��^,�d��^���uʧؽ���}�aF*��,򵑥���$��k+��γ\��F�:����跓���Ι;��	�
+e���qv-�|�>"As�G�8��S�p��p"�|W��u���
 ���i��5��єUچ��@sA��ﶏւ��	��6����>�*��zD�֕W��^ �y� �,?H+I�Ni�f�Xx�y��Gr2X��Ĉw��4||��]����M�����c���uʦ���2������v1p��������'��t2��x���^_� �P�Q ��Z-2RR6�j�� ��N�K�����r��
�Ʌ�d�ƋaC{�S{��i /ZI�GJ��h7N�+Qz�5{�	N�s%�<�@�Ș��|�n�r��f`t���2���)8�$$=Uv�}��z�,���^��h���,?���T�R,	@ъL���S�-�����%J;<�����b"���9Jh���Y�l�V<ħ�#$��
��y-�/z+���H�M�ч�>^��I�|IDİ���'i0��t�����[[����y�`�q��.���gn��1ښ0=�{\9bm�#��.��mЇ�ߒ�ڰ(�������������=�	/s��Q0s�rݴf�"��B�Ņ�����pS�������	�Է>mMM$�,u/�E� ��h��+�����˰�w{��-�y]=8b1Qx
��::�x�l�nҸ>E �Y��Q����t��C�����ɼ����������56��@58ԡC6�%���bZ�JnM����^��ԫ��T���6	z�z*7h0��Q�����F�M���1�Ӄ��b[J����S]�BLJ=���5&/})Ah~R�L\�=y Ţ'�:~U�s�`=��'��π�r�oY�Z���]��V����'mPz��T���e�XR�K�B%���f�vŖ����ͦj�Q�dǝ���[����-�q����jJuJ-�/�gre��U�no��x&��*��g	���;bH��*x?�Z���{�rB����DE6�9�O����WX��O�˖���wT�0Ɍ��m���L�L�/��EӐ��az	�9]8Z���➔�x�Լ/���븜�����_�q��,�У <��j�^�J&Ӣ���W���hG[�]��������`.n|�|����u�jq�9d��ť�(Lȿ���j���mW���JEv����0��ggf�{��2�9L;�#�>�-����%�I/i����Yܲ?�׽H���͘�,�n�8k*+�?��N2���ME!���E���ċ�{�0a(E��~*��i��-,Dt�H2 3��¼��î��/Q�H^T�F�����v�x�s���h:P�P��eiӚ����f�N��K<� ������f1���}(=P��_;]6�^l��$S=j�k��{��<hqՅ�#LՂt��B1���b˙��㐷��rz>%6	'"*�w{Z��fqU���+�� d��Y���!�G�I�T-JƤ��3LqB}_��S�l�v�k�pG��2n I��C�f����#b�����cf����c��c�T-�Լ�:	~h!���]�Ջ��@|�<< �@v㛛�>��T�������8��n��R��Q����@��[����؞Ƅ��~�{�Rv�:���=w<\1���	11)Y��~��7 �����fѱ�e��xټ��&7:, ���ۨų����^_p�U��	���P9)�4iٹW#�CI��k֕L,�1~��nf����#�)���'L�%���������Y[~�%�"<���+N>��HdBy���Y۳������9ʀ�!�qՑȸ�~]�8z��"���K<��m>�({���LE�+$x�� ���li¯��w�rÉ-C�%"ܬ�|�>TÝ����;?�8@��nz(��<OnK+�w.�֞G�T�l4ky߀#�6���|�4o[�$p˔��b֌�B}��\�A������[ff�1(�7�\HMwwq�ӡ�� ��qG@Ȣ�w�z�̬�ut�u񒜜e�_K9]�Je�2��W1�1�����yj�G�;-R���Ű�?6�dH�b=7e�ʑq\L��e>�ֹ��?[p*2ϮR����s�������J�P������g�y�J����UM[{�1�J�T�А ר*�pFa�9ha!���Ơ<H԰��ئ�K�Faۃ��+?���A��\VJ��'���#�b��+�����g���P�`Z�8�Gѯ��7���$�*���1���S�n�S:K�c���v��P�P�S.�Xa�7�eamm~�T׸��U�v�]P�f=��z��� n8BO�m�?.�b8�n����hWMG��.V&3�֑�1��y�e7ӋJL��Ae+/��RF��Ɔ=�WWH�,F�>yL? 6͈�M�P��z�&�,�G@�ާT:�G�M������Z� N�W��bȠz?l�+�L�˧I���@:���K�B��E�����9��tY+R:�f�薿'�sjk1UE��TEo��1Q�m��G2jVέ�J�ee\p���zq�"�)��O�Ȑ}��Ed�¨��6C�A	3=���0���'�17?�P��җ<1)I�Q����O��1u��9���F���J?9�uJ	,--m멅��lmm�tX�%�{�5��P���wU��3��� ��.g����G�OSt���B^Cs�j�**�%���	V�������|6H��<��;�U�$C������G��t��`�4
�A��w~��<���FZ�����F�9W��X:_8Ya[��A���}�%E������f���x��-���� ��oϋ�����3Wi��vy�_���]���M�W�0�E9¬�.�m{u�)��n6�7Zg����0�f'N�r�����7�`>^n��=�V���B�vFә�_���)؉���v�� :��7���)��(Y��=���*����J�OU�����Xr��):2�Q+O+��b�F!A;6u�b�L��� I��vLi/�{-�6n�	��7l�`���>�67m�<C�\�gV�	(?i)�4��m��P)#�hX�S��z�Ƣ��'��C�g�Vo3))ħ�10��y���Y���������F�3@���Z���p����I��wB������`V4`��b���R��
�(��o�o���	��E�"L
RH7��m^��h� `~��a�� ��f�LՆ@��ݑsY(�S؂H`�e�xon�ޭm�R30�f6+ԣ�UW�2	��am9��P���;���_[v~�9�l,���xQ�lZ���6n~8�ps��$	$�]'۞mW3(D���j^M_��1��i�>&�����Ѿ�>�+�BU2�P��=�]%ك�=J7�>���xI"3;ỿ�%ڥ�[~\��WFOy[^�[����<�pέ��k��j�:�Z7�P�og�J+��ѧw�*��c�ᡣ�|���.�bơk��e+����9�!�=�*ֆ����m�35Ģ�xq���X��v�{����ۇ'QQQ�9 ��K*��W�.c�`�o))ee��4��<��gYf�Z�}|�z̰�#+��ɩ��Y�,W7Ut%��11��sg�Sww7�ߵ=��N˹��ЈY,�/��>�ԍ L�A!}?X�8�=;�
�P��Fb5�u�9�H��Й1+-P�3�{����]�|jz:!!�sL�J_��	�{��6���//omo�=?=j�SrZ��c�3-"3���R��n�X�����J
�� �L�tk�)�m����> �G����"89��`�� ���t�8���z>^���N�-��Ef?�\��!�э4���!q�'�|���F��sI;IG��ˡ�z�3q]D�Gq�w[�x��ӿh{�hO x�[�a���+�;0@+(H�&�l䪿����쯒��?2[�����4LL肙�*Eh5�1SS�qؘ��إc�JHK�!I ���|�O@��
�R	��������aƕ�������@�����mn^�lۖ�^!@l�^T�r�c2�]��˨_��~��UIhurө�H��?�:X�+���rq���[4��4)�_y�z��r��������HI]��*���Uqe%�5{����D��@��S7Uiq���i���!����8a�B�f/η?����r�m�!㴳����W,Z��p��eC9�d�!�L�	�ߩ�%������^�y��&cB[�DPf9�|�|�j��\�̈3k<R̼������s�h�Q���yX=JDi��A����1�w�#�.���&����^O@��[�N�/АP����oϷ�_�˃��_�x@�9���z�4AzS K�V2�&�M&��m9vF�]��G.O��͢���l����ѣ#��ݩw�I���Mj����a��PJK�Z ������$��ڧh�y�����'�8�'�-�KSM������p�\��� �l��>��miGi�V�sz�Z�;��5R���뾸� <�~qc��z���5B�o�4:�#�C{��)U��,���(�w�J�I�(�ex�d�w�K���`�kS�e�տ��^�����+ȳ��:3�@cZ+�tLO�T��4!�>b��g-�r��y�����g/=���9t�Dħ�lT'��@��m�d����@�}��zODEµ�X�譈ˑ�+�c^e�]��WY�p�x��~-p������h�(I��K���������ؖ�\����([fV.T6Cn��~��M}���,\�i��:Jr,�g�-�6c�� P�� ��k/���6i:�M�s*M��D��A��-��������Z}�M1"���k{���H4��������F�+�K���� 2�:QJ}C���>)ҟ��[r{ O�ntcd��;;문�����Am��-������is;��'��ɰ�2�Y��Mlb�K�>��� #�o#��VD���@9���)J^ D_�ۻ�$ (��o�6}����Hv��鑣�Ģ�N��O���&i~�d����E��"�����n�E��,��z���u@~�g㔊jN�޹j�h4�4�tJ!_�AQ�:"���W�⅊��f7��s�"Y˄���&��$c��e�-�p������J��b�@�/"���&x��g!��6���ΩT�6tD�/���%M��Z� ��
�g���G�t�ZX��),N�t}������\�O� M0�\�^�c9f������K��ځ�L"��7�~��Sќ����D	��%�F��7��z�ly�k��1���l�A�^C1�|Y�cIW��My|{��A_~39�NF������"ܛ�����7���2����w�n�ro �fq�ݼ'P��Y`u�3��<�
m��j"�k���s,�ߠn����nB:���~Zl�XeL=~"�N���Ӊ�'�Ӂ��]�������ga[�� ��۹:�U��p[���Ż\�Y���JD� �X�r�rl�r٪���W�4�:�����=�76c�ܹ/Uz��J����v�}�[��NFaA'8�7?��*mk7�2n�!�4Pt^��n.E� ee�
�^�;����TLo�����A���u�do�(U�P�cXOLx�S����%X&���)�$\�2���Z=5�t��9�p�.?�I��.�������;�~��ý�_�Ka,����:zٗu�AǗU���FlE�^��b��w�pd���%�0�,����~s��}FU ={5�<�]�6
��]'J�d�h()/G�D�f��_�d-�,8�9ی�MƘ�-|��z���z)��s����aɨL�7���漼�d�Oo����^ۧ�B��v1�Ӵ�`(�������u
o��g���ג�تb��B�9y<����b�y�H���LEwX�-־`f�����}o�XϚ�(��f#�JQ�x%Np�Z���# DE�>�a���G�Ov_w~��O@%�zDQw��ͫ�Z����8�-YS�S��_Tæ��)_Ս	�4d�6Z�J�$�#c9+-�߿s�k�ob��[���2��J���xQ\�����'q�=����4�TV2�_���k�Z���X���ē��OJ*�\�F���nn��D��V���K��7ׁ4��tQ5|�3�E�D��K����U廋EYJ��ka��1+�G����'�k��/�,����l[��>L�G�1
�B��M�����Wb�c�Vgtٴ^��~u���?1E�g� ��������`~�72��L�g~��/WM�z��"2Vΐ�b���*�B.��V}֛��B�N���t�a5����
�н\?�Vʜ=������Φ w7�h �Z���1{����vW�l��k�nG��,7~e߽۱���.W��:�k^�G��K����wGM3�W�|��]�c�^v���{=a
�'1]>@ ���IG-���H*|Ƕ�UP�o�1n����Ù��V�\�T��,�6PV�����+�_0���`M;�s��<�����trl�x7:u��a����E��b(���!uI�p��L�wgC�7�)11r�=~	����ya�m�L~z:�$�J�2��A`��{U���<m=�2�+��T�bA�!����$)���"$�:O�2��݅Y��p�v�V���݄�i��y��SJ���C^a�)��C A�n����TKA�c��'x�4��ZӀ�1e�r����a�Դn���{�j���癏O��!@c=9z�p��f��H������!��t�y��7:e2�K��/��'�U�������b���8�K/W�3X�<�~V�����͒������AhcL�J>���K��$F�g3��~����PW(���OG�q'2�Q��)NhȈ�:�̙������WD%0��}j��נ� "�'�zvj�?#�s/=�_�n�j=�0x�v!c,�w��C!����m���5��_�>.��Đ�:JP���7���,�A-d @!U���8���&%��ze���g@cd�3�?��H\�����5��+c_�6&�^�f~��s�cC��:1�$��	�p�M9m���b���B\0�q-ψ�O�¯�����xr���EC�Y,��V����;���!�	���9-�͆�v�zϙ�%ڍ������]ztr����]�/�RX-��>�H5���4Ѹ�� b�H���i�+�mWE��
��0��WfBd6�2>�n=]&8R!��(���W��_8t-AE��c��䣎�IKK[w�	�Ig�����"�'��G�$�����Ւ\X�^;@ˡ�s����\�:�S�_���v4���=	kbb.o��ɿU����R]O�h��S;=ϙ?l�_��vΩ�R?�pB��+����ľ��/j�cؖ�"�����'�⇳�5���9��P˲ݏ�b�=x*E\T�V��Y�d����M���F��~�wƚ�+s�n�	�eT[GϏ&U$-�g�T���~�AX�/M��ܵ	�b�� �m�`�_�&d�A�re��x����ϴE,���;�����> -s�9s[���p݃i���4�p�CwY�6�y���R�"onnq��8h[�m���3|���뉎f�ڃN�K@�n������ڼ@g�0X%���.���v憘\p�?�ެR�*!�x�Ɩ_��/r�q��ú3�C��Pā�54�P�)jz!���t:����hZj�J�Ԭ=���Ŀ������(��\��� ����&�ͭ�N�`|s߃�f�$�����y���r�wa�	6ʤ	�!i�U�n8�:S�X[��2�,nM����ީ��3b���=0k')،K�f6F(�.vD�\���(Fm�0&��Tf���l���cQ���X>J�
��PN������>���YD�(Ks)� ��8M��͈���tK��߄#�=A����m�u��؀z�ě뵋�t�qf�Ӛz�� �^e��S�U��ۇc������{~�ɪq��=��Y|W�C���yq(G3��5q�n���Ki�ym#�؂�(xu�o-ꟉO���#?d�z��Þ��"{�X��դ�d�>��m��-A��er��	C�fs�k~�0�%��X}��Pސ���{��Sg+���#{)����a�HS�v(���sM 2���]K~��������y|�����K׷	�>�k�7��_�ir��n�	��s���Eڥc�Hj��9�+B�&B��ů�/�_R	L2;V���U�c-��/��|��^)-qu���_��I���sr���)T
��A�[��^�IQ»�� ���M��u�]�#y�O�|�3�"чi�&�	�_�-���:�IEZ�:?�z�ty�G&��E�˩��]{��������?*�0b$��w���[#�Fq����S��oG?�e{�Ʌ����K򓮣6�WJ�=��y�\++"�s�4���h*���ȡT_d�c�H�m��(��ݭ�K}� �F�-� ��Wn��F��Œ�'B;!D1A����1�7��;�Ɂc��"�vDB��B\�c�MY2�fz���7)�L��q�-�+�'P
�X��z��ɰCw�P�̷c�Lv�jI�_M�1=�z���7AK�~.���a�A�x5vQ��pPYv�ӿ$y9HT�ϲ��u���D�$�f�P?��yp�
�2H�L��u<�`��k{��t�>�Vup�z�]��H���� ���@u�&H���.�;1����_��C�*��K^���d4�����y	$��D���H� ��������l�=��d����۰t+�C24���|�L�<�_�7ڻ��<���SV��AuTqvˉ�~�LlH�j_[������ �u� sq���c��U}Ľ��y��kCˈ˓��Y?D����EFYr�9�|�@9U��t0��� �g /��Y-df���y;NR-�o�Աako��#_��3�T^�V�"-��؈4�=�!MʎzI�oҖ["�=!<v"kJǡwk��oSnҖ����v�=�֪ϙD�c�莔����<�t����U����n�w�����%�l���]P� �z��q�g��d���6�bͷ��m,�����N�œ�~��4�u�a��@������ׄ���$��beZ�_^�{_��М���T|�������Cyz.Wh�_�~l(�/{�;
�!{a������Y��ޛ�Ğ�1���M.�
b�KwY��#x�c܎�j._��h��פͺ���ɲn{ƿRPF�)�_4�Tii~1^G�TkK�f&��6BL��,��C>��G����(YF	4�$�	����]�K�!K*t����ٙ���2�9���+�s��4ж��k���k��mܾ�,�q�Y61����v
KF�~9�!���5m<]v�@#���<e���*,��ms0���Ĵ�L��6���Ϡх��J���ʶ��)��
��u��S}u��5��S9��̂�!D�Z�t�ۆ�]����t���������F:���{Ʉ-�m��V��e�֨��8�nP�Å&l��*T�U[ݢP 	���x��˱���b�f���ذ���� �B�Ԍ�'�#M��Sh�4Ȑ1�xǹ֡���S�L��[	�.4*�}�̚y����
V�@��hƳ�P��w3*E���B�K���,�Q����k �\v��:�r}����ٹA~��CE���e>`����Ub[�3%�tJÀ�ǈp0���紙�IGB�;z#��p�ʌ����>���w	�Q�a^�����^R
B���{#E�9�O@(dՑ��l����R��9	M,3��=)T�&�#��ͥ��`
��p��{�t����1'���@�����i%��+�(����޼�_��ݬ� w;���݈�~�Ϻ�;|��ߋHWDs���*��'2_��x��@�4�+�6C��癩N������ �Ğ��s�G�^B#J:s�
"\�67�,��Q�\��B����#WD>�-pZT� ܼ/�-�����0+��(]̎;+6t�'o���+r����b:�B���q� ��]�T���
��ki�6��Y��Biq��p��޳e���!��C�ڤ����K�D���7`GD�F(���0�8�w�r��ފ�QbC` ��Y�����}VS$�;NGR�}��r��\�dVa��8���G���AK��n(6��L�"4����@ʠ�
�}�����"�.��^�֓AJ���&)����om~�r��~qb�o�ZS�Տ�3�þ���M��g��/�L�L�u���@� t耭g��Ƹ��n���ل���գ��R[i��c�Q�rk�
T�0�dj<�-�9�������'�H�טo5�Ԭwd�Y����S�!#�U�5�7+u͋�W!r�bȮXxz�|b�^�����>�����N�s{��9ϷO�����KSg���՝/����WT�e��(Y������z�=��=,��c�gh�B"v�_0�%G�����G��J`��	����]{��?&z!���'��������$8'����	S�����ZD��q�"I�vp6��Jo�^s{��_��[��ǲ+����T���Q��n�-��H�w+�y�y��������m@�`��$�ʮǱ��f�#�h?4`۵)gv�W��m��x҇8���Hr���Yz�s�^��c�p.�O��U��T��:fc�T����mۨ����Ku����OK:u�W�&M����g����]>���~1�Ϯø���O��E�֠�Z��U�?��m.+y�'�Ef����ڲQ_�z��,�wc�9d���eSq;e|w���yXɜ��v�|@c��)��i����q��b��`������Ds�I�픡ưq4�Tu\��7�0�nkf���=9��׫�(+>���6IIIw��ꓼ���|�sN�6�%ON��F״jc������옗d'T2��@�6EN|�+�J��qk{"pM�4d@�k��E�lm��HǷ������u��gO���|�e��A5���7`ෟq���D�~�~�/���I�w@�����`陠l�);D�n�����*d�R�����.Q�����Բ���Ϯ�#�M���a3k�^�&�3GX��:A>o�Mj�_@`�I�ݚt5L:O=�����^l'��>�'~���z���z��L�?Gym"�~'w�F�������,�ͻ��d��<��V�����ϒ4�(�3]�R$�ga���ӊr�F/&��wW�z�@�ɸ��������l����WF�Ҟ�(v�Yw������A�E�����|���̔���e�\19&6��o�.|�$1���qm���y���8Ux�Y��$����:��V�P�D����]@N�;�$�91_͗o��
ߟ�.�?~��-�·���U���4�����f�=_���1����fH��S�����Puu|�.,�%�pp�|@��W���1��g&�ɫb�h��⣻�>1�a�5_>϶����%l�|z�M�l�m�%�̰��x�%j��O��J8o��;���.-�xJ�U�����C�<ʝ)�z~�>��,IZ^�c�U�Vt�;����غ��z��MşG睴�P{����p�̋<>�>����W8Q��Koo�]��n�$�:r�T�?�Q���-��Uj�(}!�R� �,6S���P<A��Zǒ:����U$���/]��V�oJq_��ٞj�������y?@��}-���ęs�W��]�����9Ѯ����F˱+r��~u��������պ�����C�T��￥&/Ɵ�0��F��܃���p�G�(?h�Ѱ�>W�A��d��A��r���wVO᳅����r�?�-e^5��L�b��'P��,�iok0���4z�繲��|�_��6�����%����uptT��7�]��Ouo@�ɥt7�۞���uXrԔ����j1d?l1�U0��u�Ȭ��4o�0�.O� 6>��j�b:K�x������i��9�@�K�� ��Ò��QUO�����|��GC�1w�>zF���� H�B���%�Ӊ:�|Y��k"�棕4���cj��w����+��~���2^��۱�`�7I�NA�s�͏� �E��cW�gQ���7�=q�B��^6�?X�Z��w���?��;(���D�$�A�I2��$q�F%�!y�� �H�4���<�H�Yr��!Ð���m��>����U[Us�=�����t����no���%��TO��\��V+��4Ⱦ���ia��a<�v�`�c�q���\w�������]j�W�=圦P�(���۷��RW�0����~&Z��J�q�&�t�@�͓WW~gȬ�Lϣ���Y����hAo��%��Z��13�ѫ�]��1�'��U�g�����k�%�]}��I��@�n�"�A���{�:%M!�uﶪ|3g
AwM��B\�DsU��Ӏ��fr�n3>��c��I��64�������V�+�#��&�D�S+�?]L�l<t�[l�~%h���Z�I����.��5�:j���(R+ޢ�m�L�)���kQ���y`(D�-h��<��W.!�ZɆTO�o�k;�ް���r�1���(ƨ�Y�^ĭsR���\tbVK�Y2j_��h !�V�&ɀ&[�8���7i�'{d>c�y�N 5�������Ɂ xe(�����r�]Z�޽i��ŧ�T�����l5=/��9x
܃�wN�5�Uz���G�]�����Kt���=[Cf�%�^U�`�6����[�5m���u�|��#߶���ޏ%+mU��	j����Z L���R��UD\��L[��1j�ܴX�D�G��I��eg�0CQ�R�?��*��^%�_��4�|��"��s��QP}�FO����)��TAF�0��[ ��J���L~�諨*/ܾoAN�0�1�~}JL�t@Cu��s�y*�֭Q:kٙ���[	�j[�z��ߢ9�jk頟$E�;���ҳ�
iP{��^�CL�"7B�ܩ~�U���<��7���)��*���!41u"��q7*Qp�ۂiFc^ǎ�f��.X�F����G�|Fק�0�����6X�qK��%�2�tۦ��t~&X��5�}�N�&�Y��Df8������G1�t3�P�� �Y9����r�>�.ߊ}� |f��D���Zьa���0�Bf���?�6���|�1U+�0��b��-��gN?-/>����Kԫ��.�BF}��Ъ��"�ԧ��~��3U>��#]h�joyn���+x�9ժ|���TO��6Jm����u�y�v�Ww��g���D~!�o"t�LDv���u���Ԯ�N��`�NZ�눛X���(:aV��j�f���H�i�hd����ۮᜱZR�m&���Q��Cu�N��j]�_O�Zt��0��IL�A�og#���{r<:�9az��ae�$�oc�T�e�� W?�g]�T�������#�ظ�ޝ�{��x�Ta��bòF��C#D��cC��K���x�9h�C�%�%|�/��.f�ǂV$�)��V�����n������>{�A�YN��������Un�o@�ki`�Z�P�/ᇄ�{���Y*0vH���n�7@����2�����a�?�u�sHA=.R�ifB�ٍ%z��ck��xrۇ�3�O�JĿ ^ꌝi>��t֓�%���k
g&�ߕ�+��3��qؗ1�����{q)����_D�o5�$If��#jxI1Pɐ�o�n��/�փݰ��In��	��aI�n'�(^�]���
0�#|:�o�Bw�mk�����SN��?��ejKO�����WO\����?f�g�.]�wGg)X
�o�
ctqa��G�{�ش�4�}��K���.�E.����r������`�� ���u	���p�F �ϴ��e�;�����{�b��><ɒYԲ
}״����v��_Fz�&�s()m��Fp뱒Փ�|f�*(�R٢M�I�r��I �N�c&�H��bn�
0IId �W��W��wM���Ϸ�9�~F2	�q8�3��ov�;�L��DL�׷A�N} '�U��c6�Ǭ�����)��_g��>��X膘�s���[�Q�����ԟ���V�{���r+az@�"!��]ˮA���L��K��B��é���7�]w�+�Y:O����f{p��'&P���a�>,����w�ن��-��� #�Ԡ�]Q'�|�Q�/��Rt���Θ+lO��	�n����fuL�2�񳜉8��m9��nYJu�2�$�eWoQߺ	�����d��#� U���5��}��"�t�<���U����r�H���yj�|&��+{ +L�W���Y� ?�f;�����f3��Nkww|^���wd�B�^��I�� ��R���Е�{�h��_��c�v����0�TMא��e{G�,�O��SB�O���Q��:u����ዎغt�$k.���7�e�Zj޴%�	yW�qUM�jH5{��f��u|oY�ְ�+ġ��W<�������_�ɏVph�r����WG�U:	% �f_��Y�l� � Z�|�3��t	m�B����"Ԝ�
�*U.S��>�j"�HxV����BU�����~�)}pLk��N�tӜ���G*���UTT =�N/�026^�����4�Z��{K��E`�?zf�O���� ����?�[�Y��" (HfSyݎnF�"�
�$���pʋ���Ő;�k2�sa,�����%����(Ȧ���'�j�-�,����m&��P�����e��\&~�8
��pf�'L�/޾i���x��Rn!o��s�D]�y�'?���4���|cZ��k�UŁ�d�rg�Zt*�^�y��2��*�{e����[�2^����Ey"W�0O_�|�qS�Ԙ�ld�3]Ű��������vZ�Z�sH�}l�� ��Nb�����#�����+K��jǩ�`*� Q4�/���\��}�1�T�������Z��I��8��cZ�~��.3���43��Yx|7*!5�A)��,	��B,��H�@�u���s�y�˪N�7[��	f>'��͓2�ٶG찧��Uÿ�o,G���8���s(�b��j~�bT�ZC.Q)�Qu�D�ߋ፛��3���{�2��`l�>�Y�j* *D���M�t�;��̄���^d
%j�$P �6��WسŌ�܈�m��YR	�Ǉ8�
�'�*���6�2�P��;��O�JZ��G�ɻKw�EV���D��:?�{���4�z40�R'v��g�8���d���G!���2-A�)��)�䪃.�i�8l'KYiE�]d�����p.�)��+�����-�X3�Av�����^���^auF�WI%U������:Hz��f����"�\��'*,kh�	�9���$V�
O�MW�T�	��v:\$�`<���=�:v�m����u�榅@��!������u�n��XˤrN�xKvj�N��1��0�V2Q
ê��
.�k*Qk�.�W��@jw]i(R`�xV�)ϯb�Q&���_��N|�;��`�9Y_�E�c+��?]����Y$*{6�oޔp}�����%+�A%�T{�PY����q���(���Ӈ�#{-�6 ���6Ocvέ����
T�M�E���t��y�I	�]�?�����v�7`������z&(�W�Zx�	"j���|���۷}>A���vW��s��ͱ5R?�[��$�p��^��O X�+��u�LL�H��g����p�ɀ��@<A=���4�����B7W���L��Yl�F�[�R����9��}�k��5j�f���7B�JG�AZMN�ȧ#��8k���Q����w,O"O����?���?S�� #�*Z71�HɂH�솽΁b	<�}&���@�d8�:��eQ����˴�I��U#_��H.U����LC�i�O)�	҈�ȭe�,�s�^E��ڋ'~��y�143�����u3�>f�Ѓ��h�ҭ!9���J�j����?2��sT�� ݚ���s�6��#uG��$��$a���̫�?a���\?��$W��7�ʗ�VB����J��%aWoW��A�V�?R�7�I3���j
xN6LM��+10 ��Ql��LԠ��<8qq-����\�1���sGG��Je|�d�yeڿ3/�_�����[�>��#l5z�P��Ԥ�֬����ݭ�\*���Ϛ�@y�8�����8K�D(������A\R�-{�0��G�?W�q	���fԂ*d1�Ⱥ�ټ�Flo�X��C�c}e��~��G�y Ӝ�铔��t�ƹ%O��[6=�<�J���Oy�)�O6�e̟�ǧfs��r��O�bxdKW'7�./�s�ˠ�uɌ��{���<���*풵+��}��(@�B��'3ZQC�p�2d�J��JһEP��O?zlOS��T�As��������+��:����L�����hq$_�YC�X�Q;�/~sj����Z����!]|��dqa�Mb ��o�@��R�K�c_kJ7�t�yc�dA���׆P1�o|*[�~tl��lCy��|=L2���~Գk�\�Z"Y:Gϔ\���q�.M&>���2^dC��'v?5p�|4�b��^�PY��|~G〙�����3��0Ir0~7��H~)t�^&�el�j{g�RZ
zVK��I���E[T�d�{�d]�
��P�U�;��x~��?�:G}���8�D#@��-�ӗ�Lq�o�#�}�G󬵠��-�y��]_JhB6S�xѹG�"�n�K�a/�ǅca�?�C�9�T*XOr	�{�vߤWaUE�M�Fz��a�+t.�����qɀ.׶K���'u�{�P�������Y�$�M�~&w���QR~Hɦ����mF{_�ý�� ��㝭���d
B�m��+�=ZS��Mb��I����Te��]O����*���[���B���8�Ql��R��ψ��5�o~^mf5�#x��u}��sB���3^�^�����T�`_���F�U T^�wy�rW�˥K�y�Р����S�g}���~����`
QS��@"Q6.�8��.��0;� ���7��k�B�uh�p��+ǡ{��)Q�ʽh�*,�L���^d���wƹ7Wuid02\:�xX΀J�. ��&����X�T,O<0W��~�5��Qi%o�HQ�%/�����&~�I�)������P2WJ?��P��d�4�=_�l@ ����er�,���sB�v��	��;:�"S�쳎����t��-^�(Խ>;Ɇ2��G^�w5v�Y���h�3ezs�>^�Qߴ��Z�� ���H�w6����Y�<�
[h�KN�߭��������Q�fx�oPu8�"��RbFp�s�� T$�]~����Uˎ��,I�)�//Տ�,U����� �S���u�K"/E�xnR���	Uh&f��h���oVa��S^[|c*Jׯo�g�6��Me�)���C�) ��b��qf�K>ݢQ~A�t?t�K6>�u�[����`��2}��U�ο�x�����u����>@������^>�;�!x�1t�+��y��ً�ȈZqތ4c����;
�Y�o}Ȉ4o����F'� �>�N�&��NZ|#��
Q���F��e�%%t��]�~x2���C��<
� ,��9/�\�о<FHT+G��g�s�����M�M��M]|�l1>�o��K����n�R�Fq��X�}M��^E�fm��v����!��O�@Dx�'t�������ZO�ӟ�J���f�u�GU�z3]�7`�)#�06x���j����`�`j�[9y����]l�DłmeuBS�Ѱ��Yԭ����T�:G'i:.c9zS��s� ��dhV�P�r�%�čX�{hH���w
kn\zC\�[�H5m�a��Oiwk��U�}�|�7����}0���ݰ�E�1��r��GUݱy��<���m�+��ʫ���o�C�$�⪢����s��/�
�+7�Yb]�'yX�'��ҳ�}�T���?��|{H�����eG�2J�e�S��w�=�g3tۜ��テ�v�T�9^� �jU�ͪut1-��Q���ژ%d�m������b�_��F��!O��4r�X���6�`9�&R���C7L���o&�,7�`�9�f���w�5n�ϒC����+��[%����k<����@����4�9�''�	��8Y�ɕ[_���3�c,�I	�% �Ԭ�B��T4�)?~�׿l9��E��I����uȈ����jJ�y���ӎo�����_f|�v���RP�S�ii�����I�ճ�/��*��8�86����e�������H.�>I,��sy�͑��h-�8�x=�z=���IK(al>?I2��D��	�e�`�7�M�iZK�rԴN���Pf�֧.�m����h���9ި�k��f%wԮ�1<�
ww�ˮd�y���4�ē����p��u����Y��"|ٍN>��Ds5UbC�i1��33ֿ�����_�h!�S֖0J�b�Q�|�e�����|r0��_?�@��8r_�0%/=<L>ޞr~�^y�F�K��:�(�'�����?unf��{�g����.F9rg�"
�`:v!��*B]C�&L�p�r����'	fS�q.@�24�'�6Mr!v�Hsᴯ�y�����fxw��-s4����5�I���|լ1���}�{D/���&-���4J�Iϳ`9�f�z���	j��ox0JЁ�i>��8D�c��ǵ�!�: �]n��B�Nf�=�^�N�%�:2�u��}�4u�y(�*X2	,�,��h�Dy2� >�[\[��'/��U�̾:�Nl9�<m��%�nvh�7x�w�ɹ�z ��f�V��A���kf����M@���zRl}���)\q�P�=���c�VS�O��1>O���΀�`ӄ�l��~Sn}���:��%N����_��\�T���GtI���Ȑ�i�u�c��9�l/��=��w������p�)@�������Z��U��qѾKd����GX�DM�6t"B�!(*�wL��J@�(F�k��ŉ$��=0�f��-�}d>�Q`�W���YP��y�Hm��G��ğpߜL��E�Þ	�bAHu��M %��8U��MG�0]��Ä$�ϩ����k7�|����V�II�Qж,4j||ąs.��7O�_c����|{�n�N�S�����3����M�f3�;M��;�3�sP��|6Q�8��m,�b���
�����ሰ{�_��wQ؃����P+�c�#�ыL�{�U�-)��Nuޖ!Pq}�+��/3�{�{��6k�3�߃�?c��ǋ;`�mYm���UiC�{�׊�_�V�hi���7��
�p�8�A����Gzy�="�qӤ��MU*�oy�\����]��mX�;�����@>����A|H@T��?�?�v[�Zy�%�n1��Ylk���߹9�l�՘r@���Kt@ ͧj���nN^��?�����o4zy
�u�,(M"���+�x4�(T����]Dļ��L���96<XMM���+��zuՍZ
Ro�h�&ז�"� �317��E��@��a�5W��B�|mE��AN�d��,��.�
Z�*%�H�]��O;^9�YSA�t�_���B�:��V ��А�+�w�a ��DY-�n�7���d�L`ơ�GXW����j�N�%>s���\�n>��\�a���JG �v�d*yJ��j��b�L#Yi``��@�RV�+�T���	�7�+���@��v��x�o���M/�u6f��5 r�ԵB����f��y��Bep�࿳��'�}>�*#ñu'���,�=����!P`����1_0l��[� �_�L��&��^�H�h3ʉgb���j��4l=ւ���8}
��1XC�T��;���Ֆ7��dԛz�=�WQy�K��6�����y�z�
�.��
7k���
�$��	����+��������5I4㳥�X*�WUy~Z;�n0|�	Ҟc�����Rg��Z��k�e%v�Uq�pG�C�B������ޮ��=��Y�����hQFY�B۰����Ag��؋�K��Q�Ȱ���5%hc𫶹�z�v.�<��ޏ�?���哾��,J[`��b9-uW����	}����*���Lېw�)��L���b�V�.mc����s���[����96�-߾)��� -Q0*�8>浿Y�.�@��ܼ�}��X<�e]��4Ԃ*�u|�GKV�l��΂
|�4�;�3����Ib�sf���.z�����:��m�x\��`�6�o5�󱎳ɫ�g�y�E�H�ɵV��ȸ��RA�T��z�ـ^���5��fr����tp�8j&?��0XH~�:�����@��8�9Uӳ{�%��m1��>6-���W*��̲2�J�@��Q�榖��g`$�t���Rtj�b�S\�	��i�t�|��1�&2������?��`����}6�	u��뮜P��/��m̓��e�l�aWi�-��{��Ѥ�C�ga�����5,�8�m�Z�Θ3g�����W�s�(�U�`5��Xwg�@r�PԖ尔��wPA�8Vo�HK�~	�;N�%���OA>��vo�C����������c��?��c��}�w��l�i$�|��v�ič+Mմ�"��?k>�?���*����W:r����BS�q�V��j��wL_�*� �I�p������E�ys�o���}6�&����^S����0<E ���~C�4'�LrҕNb2�	B^��r&�n|K��Н�Yz:��*橗�KC�-���'��0]�{gI�x��*�@Q�>T���?r��r���fC���6&��C�r��v3�W*_Q}��ε��k��o��� �q2ҥ�Z��]�؃�0n�6�>��|7��7��0ߺEOb���=4�4#mp	��Y�<M�1��eͦ��K�~�Eܨd��������u�j�(L�>�a�T�`N��:H8���vm�~HT�C�����|���@�qJm����>*��=�jY��4d�:�hh���T���7>V�O&��^z�&�v�}>�|�=���kP��ډ�Yi�]��m�*x����6��j�|���h�Ӄ6lu}�ħg*ŭ���5eq7�n}}�yʫ
,#o6'wMy5.�rV��xTGm�(�b9��ݱ����� UJ��$� �D�䄝�򁛷?]U�N.q{�3�`�ț���A��ln�T�3m$*�ӐĽ��Ԋ���a���ДO*��8^��xH0����	1�3��є�c�y��C��˭��C�W_�nW�٩{(��{$,y{�j^���h�u]!���sX�V_�SV�Y.[?{S�gOW��
�o�<�\��}�U�ba�&�S2��Qe�"�d>�F,J�.��I����nh#��(����o8Q;}�;k}v��a�scXP�#q�cp�B&a-U�Y�D'�l�gY����d��7~^v����씣tϽ�ߋi|�r��3�j{�MBy�	�����W
�xnѩN��e�:�ᘽ?�p�$�W���M�	[�"$��3꽪+�K�m�Y�W|J�ben1���{N���}d�&�[�ͦĹ���-X���e���2!yR�'u�?NW7�4P߃
�x���x;R\���tԠ�M�s�L���h�v�۽�t'd��;�D�R�����Vhn��<���	2ސrou�	6�� �[�&��Ҏį;	�gM��q*t�F���]�.,0�ͽ�_���u�����ѓ�/�mx[��󔚊��+�*,�FP�Z�S9�� �S�.C�;�a�s�����׾���峷�~W�������yv�������n�m������TQ�+���fgp���)�;q8�~�r������1�/#�N�K,H��PvV'��b��Iu���Z�Ӿ,ȴ�X]�~o�]�i�#��f��}L
�="5r�����ɾ	T.��i�3�k�������ee]Ly��8��s�<Ĩ�"�@x67���|�&t��e�w°��Q���%AH �^��,�\I�����f��ՀNM�K�W��r�������|���,E}�O%����IqUT�!��1/�
�#�^�
La��P)_"�4&[jč��޵\���������9��90�A���g��3��@��}�)��;�w��!����j0�8�k*�Ũ[꒡O<�;$7�_��t��I�i� �Z��T��X���V�k�C���=j��~f+�3;͢ ����,ϣp��Ad���2���"�8�aX��\�07��E6�`��@�s{L��F_{�d�X��B�1�|"Q,���M�f���@X�������_������5:�;�(�$h+�n����`�^j��!�a�+��ŅX�{?��A����������ϲ�������pu	$�u�N9�;�*���(K2c7��}�ʗ��`�Y�f����+c\��ω�>�؊Ԙ����}�YY64wIW����R(%n��Z�h�,AM�]���"-�=fo&���aoǆc�}�`;��B�?-�!)Uhىr�+�vG>�5���$e���^��"_{�O^r\eߩd|a��$J\|c��#��Y|�~��i���<e��*g*A��'<r�0Z=Eдk�r��H��H�cK��u.<�������Qʟ����dF�X�(���N�W�֘5�� n��������G5��Jeښ>S�1��N�擙�jE%��f��t���x�!�{�Je��>Ԗ=ut���e����=�P��Q�ŏ�r��z7Ƭs����gD��e1A{U�p���wڟ��ز�L�F�f�I��l��0��g��(DsZ�������O>N�-Y��u��w�?�m�N��uV���5ƄԴ�md����ݛ��g��3�i� r���V����4�R�~��nvn^7a.:B&�_ʖ?�e����G�S��S�hm@��5^��`�?��Gh&�zz�ɭ��1�e�����B&ſ�,�����]�^r3�?	\B&q�FywNҡ�{/c���pd�hޭ�_�h�dJ�V6���b�כo��i.�F���,�c{�eG��ψ��{�\ �]B�G���Y)}H{��	�Ż�*s��u1���s�\�ZC���q�ǋ�OJ� 0���D�!���7�� �;*�� o:�R�w��.�N�e�����.yQ��rCŬ���1��gcT]���j��>-�0rOeю���G�~����>�ȗ/���3�
1�R�P?LE\ ��ܴzގS�K;f|`L����:7�d��q;�@�}��]����H����X���o�oD���~̺��x�l�ݟNb���}�@j�S�:ݒ��lv?gs��g�fr�vXמt#<,���g�'OD��`~��/s�����$J�^�&�'����y:	>f2����SPI�����% !;w/�A���{�5x�%����^�F��h�9�NÁ�~%�����n�T�����%��>IKض������m��Un�E��h���}:�?z�g�6�4�����~G��C��+�k����ǣ�Q�n�$�w���m�1FF���a��u��J�;������������ɦMhe���Ԍ�!,z���6��F�i�sQ�=��i2Z�A�K����ñ��	�@�6�����T�y��9<U����@���ay�wCs�K��t�gh��L&�v�LZ�%�L�����(_�(,c��!�^\�Ñ�rndU2G]v��-D	U�7{�%�2�7�� ���p�"��o�u���9-憎;�<�]���s�7�Ӆ�,N� ������8I}b<;�,�e���<��i�ö[[ �alI��e���ܞߜ`����\8U[,���{�\����{�g�6�?΂]���ѓ5Ż;$�����Y�Y��\Ue�~���4�~�1�võ%�#`����Y
��:�&�~)޿Y"�;��}~��U��h�gu���PK�`;�����!��n�6젙���Ƶ��
{�����ˬ���I_Q��+�_ !k��,��0��e�Yi��a��Y�u��������М�a�+fy��b$8�8��+R�8O,�G%�K�i���/PEg�����GcoN#d[�O�]9>�~G=$ƃ��\�	��|e�����M�O#Vu{��xR��~���!���6�s<לO�w����F7��PN���+��D��wO��ѥ<���)6�ק�ţ����I��7m�+�:�G�2���<_����L4�n�b���Ň�@�B�R�PFF��B���F��`1k6z���;n��R��W{���zc-K��g���\�/.�k���b[0R��h�u|�L��Z�W����S�[��1w�l��'���K�����#�l�d�*!�8Ze>{=/S_�� y[����t"��P}�����U�?I˪Pp��]Pj����Զ�dZR��̩}��~,=�!Q���h@��A�x��Q��d����I�3]F�}���E��p��|�;���ix�IJ��h O�ƥp�D�fP�q)1.�S݊���|�Ad4�ڌ�b�o���� �n���_��@/[K?�4���O>	~����	�K���H7�*�C�$�����y:1jn�����x�o}5��.��B�K8۰4�C0���h�6���}g��B?����%b��3x��z�+�%��(���/�쟵���ܯL�2!G�jڻ�N�f�\��n-�u���y��X�ثC����I�5Ʊ��a�|�_���0�_0!K�ڜ�~�fF��tj�F���/���̀�2��-�nZ��ݰ����v^�df������#�+�g�	�Z�͈�U�m]F��w?�!R����!��o[ i�^L�	�r��B�/X�R~�Ȧ�/����	I�$��i��"E3*�#��d]��Q�����ggg~w���cb���G�Z� �[�_z���'��8��"y���*e2]��:������y}���黤l���(���+�|��Ds�"�K3omO�	�Z�k�'�쵓D-�I��b����%Ļ���F߈�Rw�ٿ$�,su��gG`���뿋��!E��8ݻ�2�T�I�9?�ا1U�v�X����&�+3Y���+�W,>��')j��v��"�E'�EO�pV,;O���t.�f))v%�! �(|l��j�
�ؽ��4Fh�pc{$��q��gS��ݚ��i{Kx8�ej*ޗn��6�:��,��V�M�`z��^��
M��6h�N5�V]���a:O{�M�d\��ީ�w���ƬW�g����-���M:]��J��A`5o�;q�;qг������Myf��e/-�q�K	}����[?�[���	����Hl���� �ʳgR�Rn�e<N7ȫ�z-�9�bak�r6�;&�r���W�n?WT_x�0kPoH�����Y ?�]3v/0�v!���6-�RG�����{�6�l�"	���v��G��R��Hg��IX�{>v�@���F:{j8 ��;���������i\��y���C'����'eˋ��맙�>ȩ����,��M"�=F��Y��A���LY���13�����P����ݪ�[>���#N�D�x� %�'�i~w��I�p�͚rf� ��)�1+Ic������]Z�/:��wM��W��""��Ҍ\.-�.Z9��@��RY/�>��mh��㨖�J'\صyZ�o1���Z]O�O��~�H� E�@�x�Zs����{�<��ѿ�j��.�.��W�M�n���7.�?��x)]����oG��$��=��[|T8���{�{.��5K=��{�'�z-;[����#l�1"$�J�G�Y�qk4��������d]�k5�ζD�^Gvw׃�(���G�����������z�S���f�~>b�ѧ�fߘ_���QK�<�y<�Ѕ
azC���2��<Z.��0/�%�{��Ki����n�7�j��RE�O��.U��/�~�� ���{����F�3���ל��ɣW����a%�;�,���<$�ck|�|q��g���AD,�����sED���4�0Y��Q�P}��:��%)��q�|#������y�o��(�}�i.t��60)ߟ8��	�طa���^����U��Iz 	�+�_��iH)�G��ߚݾ� �Ө{Y^�OZ�WD�^	��?敞��>@�l>�Up��/��[��oPk���~r���A�z�`�Jhԃ�~��If)�h���x�J�����k&��s+:�Z�kj7����L�'U�Y���ͰZ�'�������i�J��ly�(�{�lr+���w�Mex7$T1&��W4,oU���I���<,��$�8�aͶ�$	 ճ)nG�{����c[�;9�Vz�$*�w��o&&F�b�~9vj�rM�LJy���GKy$���g?�^���LE���V"ǋ����9�H�~�J��@�u�~��0���!��m�10\���q�l}���0O�*B��Q�^ �Bz}�̘;Q��y��f�^?���Y�>�%��`+���mqw���K�={��_F�܈^�`	�������=ߋ7}tk$\���h��8z�D��>X�_4T�՚����q¾�~����k�o��
O��#��M�Z����^/���Kq{1I�=���^�pa�E�CR,�`�߁A�)rqc���㤪�A��u���/����U"�[����ޙr����|��{T% ��/�g���i	}DkD� y��qg���Z����|ז&��:��>�H�W���Y�O�MV��MM��b�'��O�M�̤��D���C_�lmʞǅ'�(�ƅ��D�E$�CSQ*����^::G������My�K��[u��f���'�Ψ�8J�c0��;�޵H��L=������Y+**r� $%vtOD؝�������4���u|���|<?^�:��F/w��j߹����A}��=�W��>�h)�[��d�����ۈ$L��'[�/O�^�쵟l�8�om�ז5�tbWA����V��{����z���GZn�{3l�x;M�k���$������bQ;���_����M�¢�������I�w:����!�i��sb�Z���	�P+���3�����z��m'W/�xY��I9�G�-$F���5��B����}.��wKX&�O�kfYX6�M�� 3�c���\�r�٠}���؅�7M;�4qG���a-��� �a�ֿ�,�o�5\���q��}��U,��W�>�߁O���Tf�N�����B0��s��ƹ}ak�H�S%Q����spݾ�s�6��6EB�V��~T���e�p[�2S��_�������Qj8Ϟ���1��b��`%�Cgo%�q��d��t�A�5z���h�`O3���&ׇ�G�.7�w�B�N4tU�8[/�t���A/�ɷs@����_((��p����;��#�f?/+� ����_Ӆ��r%ђ�g��.��������[~���ss�bW�d'�=�¹�m�ur�]YG�K��SK%9�X��|���n9�W�Ƀ���QM����R���R��8��
?�Z%ɭ�^s������?��)�bN���l��b���蕱;j0���݃�%������������Z�Szi-��%�J����=�}��keZ"�������\�K}��F�־��qa����A@_wM��"Od����`g��~�?V�Kz���j塙/ث՚��^t/y� �d8��$��k�,�ձ�y^���op��-�h�Ud�enw苫���P�вj�"�����I��W)�~)�9����y��V�4e�Mnl������t=�%�"�����t���-�}�R
h��&��'sI�?�k��K!2�S{��O��^3�`ӹHn�H�:{,�b2����P3i��\�8c&ԊN4�|�k|W�\�h:�:j�%9y�#��`7���Z&�M�5" �Ƀ���Z���C���I�Y��k����|�r|��P�(����쌓`�|��3�:"��]j�O�%���ۊ�V��v>$U��D�`k����e���bލ�/��9.xR�fu��_�,��*F�D�p��~n�x������d$�}��޵~�d�q"O��v4���m�ga�g���6r/9��7k:�5=LtعM���T�`�����i\컸Vni)߼�{�9���n��l!8�F�/�Y�C���Һ6����	�2Ȇ�K����O@,[�I�3�GW��A�v��T֡��\	0��=>�h;�����Rҁ���+D�/nw�����4����jЅ}w%���tӧtÜm2��=򖚺����^�b%$�L�Bz^�SX��O�l��w����O��42�C�XZJ@ZJ$��Kx,�H��Rt,;�2���3�@T�_�`o"�jn�a�;c�� :�V��ysk�'��d��+M����x�����6������q��e�z܍���Jҝ �0��t�ߐLs�M� �Z�߄^��/DEo����%�@�l�A~|����z�}���)%�'ao9�{K�������r#S���O=D���n1�bk��s��������Gϥ��T�SƆJ����lk�:�����-6'k�� u9c����{�k]�C���<����o�uZ��C�<B4\�� ��^��Tn��~l���[�$hA��[��k��O�c�W ����wM���5ɨX>����*���8D��hq1����̴�ƻ�&G�\F睲'f�,���W�ө�	��j��f�ÿ;�# �1��%�7�~�Dh��T����WƟ����#-���o����X���ȋ$i�'��)�ݪ�	�9u4�|Qs�$$���1�Ѐ;8Z3��p`txz?�!���TW���ǿ���D���"�(� �J߿�-�����"�G�`;Y>��E��4�������w�qj]�r��lR4�Z����������_��]ca�:&�k��!����\���0��ږ���G�\�.d��wH�X>@���2(�&�.�{����n	�����<�{pw� �!آy���U���?[s{�{�i�魻8�;:�q���Wz��ZE	�S�{m!U�ݒ0T���.�JWg�N̾���l���ZTs�B�S�|�b 90@�|�o�Ny(m�W#y���u���!TX�u���{M�#3Ӣ�ۉ��m,�	�;vE�yG�h�8~�~�Hj{�[.��H"y:�jĥ�գ*ޭy�g�B6�oI0`�
:�y/<X�	�}ݬh%{T�z����j�<'��>,�Đ�[]��mr��!�LeR���G�[~	3"q���-A^�v�̀g;�@��D���_��?��>~߷;��O�R��~���L����#	LS�(HA�G>M]S���7f.g���	��ri�p��g�=���S^Ə�D�{I�6h�6���W�9M�O�u�+d��,W�G��t��;�Ð�Ϟd#���v�
}5�P��%��p�qL��ۤZ�"�5���W�B°|ZT-��z��D�B���_��uWq�Ҙ@�x�5�j�+�m:�G"�� ��r��L*�r觿yV�A��$	�2|W=�-4w��
�}�Ӧ ���L�Y�NMቷ���_y�E�����j0=�,�O[� J�G*T����f,}tUmћ�)��q&N��W;y�{�Q~�kGx#�ҙ�մbj�-o� ��:oW���˚`�P�ö*�sH-�����Ą��%@��?2[���D��_��H�w�T���B��+KI����
�����o`��ޘ�>07�By��I�7n�ΐ2��L�#Uގ-���l��}�o�}Y}�"�����^�2�&2N�b��9ug $�o!z��l�����2Z�z��}(���u�:��%ڀ,�ʒ.-l~�AX�C2s�&_s���U���թ������'ɲ=J���6w7l���+\��D�	�zќ	�Dspk�8R;�)0��^��_'�!�n���!g����?Ȏ���	z��sx��q>�����;��^�5a,�˝�r�M��|�O.��\i���F�f������>���������䵋�~�&������`V!�����[��~��n$Xwނ�r��;���Q���}�C��Kp��$����@�׌��M����]�g����ex�m)J�n//)���ְ��q�����G_�f�a�t�wꢈ�Z�z�#V�n:�H�ݿ�qE��vT�	��Q�c?{��r��dE����!�W��1��Ls�ş�A�����˰� ����ۻ��^�:6��_�F�I�A��hzȴ_���t*>2�%�7!q<��t��1����1XL��f�:��vA�@e���X�	���>ڧ�˾��r�����Â�Djt��HӺm�7��[��~P㗗�"�t��b􅹘`��xS��v�O����h:����� s���yz(��Q����M2d�_ l�-7),�{��	v��4"�dײ��J�񖞛}5�x���z�C����!Ӣ���e�*b�*��(��u��-���L}$!!��<��
���?R�3Q��C��W%�;�J�"u(CQ�g�2đJ�ɻ`���r�]e�l�!5�i�������?�--,D$Ȅq���:�H�A^C�on�� � �w���4/E��C��{sf��(p��
�u%l�;4�t�uBڕmx�v$���Qb���p*e�i���p�	�[�����k�@�d�;0Fp9o��5�|d}�����<����5�@8 �����ܟ��Q^�/���8��)�eǂ�x�ز�l�Ftj�Kt����+�����\�m�fJjrΡ\�Rl��Rf�L�{���(M�E5��eE`�{��0�w�-$��W�>��7B!��C��J�������n>��;ګ��//�|G��?�$]q/ۙ���Z���۾E��zE�vk_��A�MҾu����!!�D���Y�� 7Kx<W�����h�n�8��Y(
یH��U��3����-ɉ�PV�U���\���m�vQp�2��!)�n���������/=�D� i���H]'�=��::��q���aDu�{2�a˓%�1��.�]������!�Ra�ǁ`���Xf=Xg��HX�����QށST�}�%�&,-URv �R�©�	�[=KQ[�;�J#�.L���G$��MB�S��T�����YJ��t����������]n?��If�m���k$θ�6ɲl8�FW�CcA/EW�
!�5-~�DЎ�5}z+�WRr��>��`G�1�#��;+n��κ.���$C�*5J�U�p�j7�s6��}�xHqv�F(KD��d/E�蕹 � a�_�갶څ�z���|����]��Mơ�+l8��p��e"h\e_�Gs�*���Y�&���dF���r��%s䉲�߸�W21�9���}
�`~���b^F�3�5H(�D���� ;r�mߢ�˦��j��ߢ��{�Fl�l��r�LR�g�R3΂�3A2�j,T0�b�Jc�z��Z��i�ãۇ���l�COSńp�R�uIa�?Q_��A�����#qh2֣:a����@Vz�����z|&+�2	��[S\��3\����Q�p�g�q9��`?��.�&-����/Θ�B�qF	�F�|Q#�a�OJb�ðI�X�A��)� �|����9z�#�z�[Lt^m�u9���J�gR�YA
�*�z�F����a_��[a���g�}����ד�_�7���߫Yɬ�;�=�!2�&�C�&J�s�%M|�G*�ŭt��~�M<GqD������UT�uj��w������6ǶJk/��E�����-�w��N���V��[s��"�c��q%��`_�J�|�+8ǟn}���k��Y����&�a~���Ri��/���ʕ�n�K�:Ip~eK\����$K��]*Ȁ|HĪ'��ի,�2{�ƥjݻ#���\�|\T/�܍��l�Ý�@����_C�i�%=p
�Dq/�n&���*_�U�` �?,�b��Ĥ�1�MwK� ��Փ=su tTd�悴�-��c!3x��H��yu�T;i���Y�hj�8�
%u���i�P�� �yS��}���Y�����<+����P��
�+�����'�r�>[��
O�U�� ��5p�E�s�p��-��)�g+�#��j�7�CѢ�C��h�$Y	7��AS'<�L��F�����Ϋ�%NA�d�1�'�\������D^{��������֦�q�支+��
z�e?/�9����8�� /x�\��j!��s8в�T�d���f5k��qep9�hu{�UN t;`T6��We!��Ch� ޲
�4�fP�G(�pG_��HM�+�j�I�k�-¡)���{T�^X$����3w��[@�[s뙩zX_ɳ��)�򿈖ܱ>�,4f���K8cy4��׫|ٖ� ���������ӓ�T�l�u��\(L;��^�3�U+1ж������A����qg�ډ�����[��)��R
!B��߰�J߸���h�2F=����Kf�W�-���yJ.��{���܎���nG����zM�)�c���ۀ�!X�]U�� @�#�a(O���6;�`�*�Օܩթ4L(��x�/L�����6�H�e���#~i�Z�.�ȇ:jd��d!E.���xNȠ�4A���cW�Sǃ�u��n�لC���#+y���i�RE(^jB�b٘�Q�O��яJ=U�C��]��QVp�?T��#�s]ڗ���^����	vd�ݫ�F��}B\�B7$��b��p�*,]�&�jb��-8%ރ��g��%2�
�;bm%Xf2��<��df�nt�%	�:RP){+�=
M3 v��n6�c,?�`Ox~U���=��+P���h���~ш�o�҇�Y��9�L�����ttXk�u�挥\�]Q�og��܇�Y��r�9�Y�?��Rk0���W��1OG�*A8�].�$:��- �6Lm.Ah!��ꛤnB��RJI��8!�n�l�<�܏e�gIh���Y� ���L�o���n᨝�'�;���5&dV��$���P�����PI�㡥��a�&	��R#ޯ;i5&NS�\�A��v8Zu%��	�l����m�>j�b���/�T�<�VL���yևȲ�*'ɟ��R;|�$A��(iX5GK�q���S�*k�oٵ�+�
#S5�^s��4Rz?C�2%�i
9����έ+�8͛�o�SJ�[�9�e�_��M���/"-W�V��X��󰮄FW�}\�8�D�������;���V�V��tj��,1Z�5l�Ǚѿ����K�x�A����r��;�[9�*[���pz;�XJd�7~���M������K��ƴ)�>���+s�-<�24���=z���0��ϐ�B�m�Պ�J�g�})_#S{�Ӷ�|ƧO��[���Yt�+JZ&�;�,���*P ,(��lm�D���P���$4%�M5VV+iBܟV;�֒<�>���gd�@f�0L���o2<g)�v�����k���ٸ�|�Aˤ�{'�&Py}ǽ��d�q�0���)�bpSCv�2��^!Tùx�ḤuC�Ɓv�(����5�j#� �f�:���dH�>���#hC�$�Q,Qٛ�Rg�!�5}W!�RC���%�lͥ�+QΜ:���̞*2�WOe�3���Z܀,�3i�x$w�=����i��~`��li���
� ͅ�/��̉��*YH+m:W$�|���w��X�t������6�^�yJ�@��,����S �(���O��ƫ�Q��.�FQ[�x�O����a6!�~�l��4��s�t'�	V��E�i�v�Sv���z�d�x��x�%o��������6�S�3�](Ć0-p�:_5�ڒ�j� �q�uFD>� ��!:O�_\�����B�ju���b��zS�������/ty�K�,�`�X[�l�d�qw���ZgV��]��$�O.�B�|�?0�	^j�`3^RJ����5�w^���ɱ�C��2c!
l_�E�/J���wG�)�AJ�	��_x��܋��"մ�'n��4$���H��أ������
��&FE����<���F�.���G �z��\ӚG�x�F�5
W����e�q��-;�1l'I}��.J�@hR�p�8�H��0�{n�{/y����9�� ���F�۪W��Yu_@��.���]>��Q��:N���y��_j�-\��E�� �ˌs,�3�h�/�=��n���f,�I��0�m������6�nS�B���ێ��z�!��I4����E�LU�K
H҅��B�h�P�9�y�[0�c��lO샕s�"���hIuR��
�x����0�5�9��N�!P���
�8���M�%�Ϊ8�WS��o�
w�oULȅP�yV��>�n��R����ԟ4lS>y<'����u)2h��5X�0U�FYX�}��Z�
�R��hJ嫻�Uh��AC�3����2�	���1m�:�p{�h��M!�/��Lx�w�zӡO50���	O�~?86�jH�b.�ԧ3S��b�P�����<�=f��ԃ���P\�k*������|���1�s`ք}���3M;��B�Ic�]X�9�l�~�JO��D���|�k��u�Ĝ�Z�_޾��*��x^�u��\?I��CT�
�MH��Et9.��وN��Qˏ�%��G>�ك�������@ޕ��yPߪ��B��1�v(���hr��y��\D�/N�]�=����u=W�%D�Ё�s�)k�؅Kz��˧=�>��#���8Ӻ��?�#�������N]��	�7�'LE�FԻ[��n���i�#�����K8���E�pQ���������eܹXx
��j�jB�3�+A�vnʋC��3�](�![�Н�>O��T����դn��_�J�xۖ������UJ*���)���u�s�BaZQ��t�b�J�n��I[\b>CC_�^�Mi"z.R^>���\ �C���2��7��[U�6�ͬ_�u�t��SN?�'�+&�5O�Z��v@���j���՜m�?��<)��?jˍ�8�0t|~TB��(� ��b4=3�U�a!O{��xs�mD{;�)�{ҕ�s����{��6��mB�[��[�@s-sYj��J�X�"h�
�y��׍�!��:�.�_�$��Q�&�4�Exu���$�J{'���*8����ڪw�����;��NQ��*�`�t�!vی�〼��`�{���<ԋ/��uml�"�K�+�X�l���;tTL�j��>Iv~�M�N�<����xfSw(t����-����̤,ӝ�	�AL5k�����c�,�Y�5d���+���Y�V�mh�"|?{��iқG_�Y��3���ߓ��l��B^��1Z�[�I���,��.�TA� �ȶ��L��3&YRw��:��1��ws�I�@�5#)9�L w���$Ql.�@u�)J⒐J���ߋ���S��9p!��{@
��9_J��%X��h�U���n%29����ޝ� ��/q'N����:�a�������FڭG���L�I�x7a�?cu�<fi��Rߡ���YX�G�<��͚�'�Nk2�h�F�NB���M9	C�g&������6�
u�晭z*���ްٟ�{�c��ԎU�݃�53�(
�����Lw���>T�ͤ{�Ÿ�ew����b�&�M}��CB�
��r}��BV�߇a*�?�������c�)�=D>!���YP?w�/�=ce�>�}bn�A:]�ob�2B6�Y/���hΞ�|�H�S��r�K	�W��� ٜ�5BB��x�.���5)�E��a�uO'� n���wb��������G��ۺ��%��EA�k���NcH�/�p��;ٱKk~V��w������B6l�:�@m�9���33�6x�}������q������ ���=m ��?�d��u���ד\>�'(J�v�da�h5��[b,#)'����)U65Z�������&[]��&X��vz�^���s׸QJD ~��i��3Ԕ�.mA���}��-ðӯ�YlL5�Q�v����:��E}���6�Y]�	�V��'�F�������3��IA���P��^Ņxd����q))�������u��@�z�o�ʷTк�����!;Cݹ�ן���/M��oѝ
*j�ۘ�4�Z�֐��zN]%�$�7���������7Q[]�ϵ}�,� 2��+y���U���#���VB3�eJ�rȕ��= ���u,�A��V��<�����Q�����l[ߕ*��,fC�������d$�4�n����l�u��<����XD�~�m��U@2�̫�6~?].g?��H�B�a%|���{��״ѭ�+̒�����6�{�Ie����ZAR�H�������
�֕�;�0�\mS�+��:��lk�ҫ��f�o!���`���
ټ�K5��UѪи	 �S�[��y���x�L��������R���*���!��l��N�nc2fm��V���,TnG��v����k�_�<�I��弍 �eˑG$))�/wU篷v�^{&ۋѤ$��y&�a��IB	�}ZZ�)J�k��ݮ*[ɲ��z�����E��}������	#�Ƨw�c(�"���GVvFq�9�����;��u����[���$	�i�J2��Ol�6���G蘚�*d�(�ڔ-~�1��(���Ti���/�^�Pn����(��;^E��as�)Sj�ڪ�ٚ5|�s�*�zƺ�]�?�8
 �����	p��\�s��if#�h��J;w�ⵦ��owh�s�jd�n6A��7L�:w����Y<��fpu�ؕ�)�q�I��ot;=]�vB��^���+#��>�����{p���;1���9 �
U�Tơ"�9pOH0���+��G��[����j��bO�����4lGX���+q*n�j,>���D�V�X�� ��G�/{�����j�$0���ƿO[X3��|���zs�J���E���@���8ea�Qn!.Hbͺ�?e`Y9���#�a��I�[ھ�K�rW���U�3��J���W��Yi\�98���*�����
%��C�W�,���o�	��(����u<l|�/̥�#|���;1,C����c��!��X-�u�ծ�Ϯ�G�)��n��`S���|��&^��[�����  '�[�6fu�!����������͕��w�e/���ߍ3��̱;���n�z(���4G�?	�;�1�Q���A<4�	.W�ߥ[�4�H�zaV2u]��'�翆b�r��L��'K'6���&F�(����O$Dz:9�3����UWdƃ=��������d��>��
�KX@�ukU�q I�-wI/��){yY�����),�$�ʏ,�{��͚��uJ��-�@bA���O[ح������$�yʽ))$5q;���/�9�
+��$Cm�e�ϗ+�U�����3�$��f[�������_��ql�=�����'Ę�La��Cn������Xc޻c�򲂩4�w-7��t���4�p߈��/�u���;�y� ֓�'/)yT"ڔN,OE��j*��3Q�W�3=�E�l��E`�	����9�򇞗�;f(��ޏ���%b��ra��v6�R������6	T08� ����zW\ 0��Ž���J _�#��Q�
��&����s,}����o������&k Vh�߿�z��<S�~�f�ί~�0��e�m�*�\�Un���Y��@��QSk������B�[A*��i `�E��i"�N�H'�d����/����]�.h��
�d`��g<�s��)�$�.�$���n�jb�a%�I�!fo����U��l��_�;�Y��sI"pˌ|��8Q��D��j@�C�]��" &i�e:�{�5��U��C;f�Ĭ��hR�2�;�Zu�Ƌo�XqUG-<��&2���S��?H�+�J+O��ɇ��Ng����$>1�R�>eT���H��Td���<���(Rs78A/%�vA�q!UM���?=�h�$|���]$uGL�}w���~�bYuL� �����D��Vԃy�F�[�G��)w}T-�tT� W�L�ò�� ��Z�/�ꩨ��|
����壬tIz��)��^�e�/�<���p� 8oF��	��`��7��f�E����B��q�K�pG��I�݇qW��+i_����3��K����9�*�oZ�(p{�ۊ�W˧"�A��8��xկ{a>\�{�w���Cge�٭j�RJ��x%��CІ�'o�@������g.�Z��zRL�ڹ���"!�m�o��Mn^�phۯG(��+���!r�!z�n>?��nSw��~)������gu�I{2r�BR��>�,��vQ�]@��
��g���%����e݆8}`��֙�d'��ML�ϔ�"�Eg���y�i�.ǚ�j�r<xQ��cR=pA7��D�q)��X�3�1����[8����3�b*���Tk���Pm��������"}.]ę���%��'���k��T�>x�3W���Լ�9�좿";��x~�&޾��y����p��,F��B��[�%���J5L���V�����#�տ�h��e��;���|y*q^�9"�ם*V�l���Ʉ@k��*�o���c��&KUn��$'�e�.1�ߥ*��Ćc;�R�������TN�Q��0�����?Lݑ�l�]�*k�?pNA��.�M�	�������rN�����з:�,&*��ⷑU��������7π��y�'�;���_���{r+Q�yf廏(�ܰ�ww#��Ɩ���Z���Ú]��m@�)���ƾ8��'Q�HX�[' ��q�}��.�w��eA$�<��x��}G�p�nӮ&Q��)D�C��׌0�
�ke�B(����a־5�u����:3�t7�8�r#\�1q�=l�p�1����(�$�ƻ���n� �"ٯ��Z�ܓ$|�9�7(��d.DX��4d�
�@5N��h;K���E,�+E�p��`J���:0�� e������D�V|ƒ�Wٜ�����O������s&���I޼l����4n��d�̬�SM����G�C�\8�?�7w�mB*��a@�.�ou�v��<_F1K!�]_/g	������[��ퟰ"	6�qi������[�|�푹3�N��B�k�3�iu�r�&���R� rpldC
�^F��,�F�H6���b��2���]�V��Ǡh�\�!V	�����L�@�,�I�sE�{��C�5n)����;��Y�~�&+��<�y�P�܃�E�-tbCq����93���F���n�L����_���y��O?�(�	�ͯD�8�/_E�3��8ZQ��`�d��x�mI�L5��
뷾Qǝ!.����K�ѕYS��2�������Bo����=��a�2�-�)Ub��I���.�$26I�����dŪ��9L%�(��h��_4qG�>�Le��$�Z�;�����Q�05'�ᲀ�[G\z�dfX�\�T_���%#�)������H���q�.�v�8�~
��x�о�)$b��:G㣐�|���.��_���z�e��ZB%f$Z\�|S��g�L&��� m�ߔ8%����E�J����<�<X�H���8���:g$j�T�j���j� `�s1 �9�[�	)q��@!���;9�����+wT�v��"���>e��(4�@(�zL�r�*��U҄�F�FTn�>YՐ����Q��TeC���Q��`F��8�$�yK���ؗ����	�PU㑓2���_+�#�[e?�7*C�Vid���fF"����!����c�k�+*����\���z��X����ɦ�^�8mx��ʳ�]D��c.�vG?����ۨ�xnnîg(X��K1�,��0.a��m���օô�;>>���Nd�K|_,�z��6�gA�A6�8i�ŝ�وO	l�U�&"Y$niݗ`�3Q�L���9������ �r0b�ׄ򧿄2�՚�YҦ�?�2\)1ɕ͜���8$�M��J���y����ԑaާKr:D[����;_���-��Ah�E�����g< "mA%B�����ծ��N/��}����ʢ"U�-�@Յ����m�(8w�S%�TT�Gxy�D�Ԟ��I"�|,	V�8�I�!�8��%ҿ�m-q2��0��@̝��������W�{[A�2�!�-�,'r��t[^��[���(��k�	����ܮ���E^�Pa���
��Ϥ�Ptkԥ	Ի�E�%(;[�V~�	=�x8�R��b�Y��1����Ǎ;eZ
��̩3��hn�"c�Q�k|*�"�7���%*ר3��uf�*���
ε�ے�{�����k�=H9�D�at9c���_�PKl���9i[�f�)��ۦQJ:�4\�p[�c�K�A��!��˥5i�g�:�XFS�5I�;f��eh7"uy�ïЋ׈R�h�̘n�m�2�Nݻn�,�����~�?�T��9Pni9+� �tX]&��v���^�D��d�t�.7D6:�I��v�pJZF��L�HkznV�1�<(S��=�)�S���R�+��ŧ�Co���KW�\�a� ��0�⯷;����g�������_�Fg�7�GU�P�N �|B�M��z��ˢt���Y5v�9#��6�0>������;�]%$��6=���QQ�o;>���	!)n$����X/#S��y�_RV�6>��r�;���y���8?�����t5B�#���G���j�g��^A�_F�Ť29Qi�}�r����6��g�%Bu�Eb}�ܰ��Q[y�k"��Xʔ�����7zPu�"��&Dxy~4�E[����;�X�e�̞����ި.�I�E��"Bʕ�����¸�S>��R�>�ir �h�۝��U�]�"c�b��8��t�ՙ8�4k��r�z�!�Q �*ڀ	�$�p�q9�/@BL���:�Ԏ���NJ����Q�pK��Jy�fTVaL�Z�%ZG�▊I׾2�_L�/�*n@��}�)��ID�Ȏp4L��%�L<9$)P��ܕ$J	�6�[ì���o/�y�+���`�D������%�����\j��,�����������N���!5���X��������0�4��u���R���I�g��}Z�W�mᜁ[VF�3�pGS��3���M�Xɵ�?��W��	D����d���|�p�v*'d�w[��x����M\����l�ѣ�?]��mg F�h	�����^�b�'�1����#�_�e��XW��9~���YLQf�Z:�jS�rC=��آ�BG@YA{~��-'<3(��(��p1�e5����۹��
ǀ���6y�� ��?����gq%;��� l�	��}���7�BߢV�ޞ��#��׷�ω�X����c�3�#
 	)��㆏/��~��$��#N����]D�K'����ȟ'�&�@�$?���8߾uE�u��/��d����G�f<>�-�%IH6��t���KZ��u|/(�(s�8W���y����,�����aU��sv������"
r�*�ڼs�iR}�9[L̫=�l�\��^ko�\���>��(]���&�O�6.k�qO��6}\�S�{��5;�y�U�-@�>�_�'�� 6D]z���\�UB=|^i��E���zY�)�y^�x��
����o�k� ��L;p���e��5���;�њn����h��i[/r{͸6u3.�D��đ��#Ω���1a ���rU�+��B�IsA֗��4>`X2?^U���GM�)��T�A!�1bTV5c�ˢ��e��z��X����N��:J�@{����GCOؖKS����L��X�[�vL�v�]��.}C昛ߧL�RaTE�I s�1&e�ń켐4���Z��߳|�������&�-�H��9k�%�{�@��λw>��҉e4Ĉ��� �o���~X)6.c��[E�����6�A�;f@mjC���DxN5�<-#�)�d{5m�������g�Z�������I�V�e���0�.��[L�:�G���VO�Q�hT]���7$�GY
��K���w��b�~3c3�ξ,�
-���s���\��3h�� R M�����|���*J��rl&�jJ�?�)4$�Q��+ڥ�,nf�"�'��!|,U�h��I�N���2�������a�1���{���f��#\�^*��e�m�g2����pz��7�Z!Z#܄w�e�IV��(e���������t���1��Y��\p"N`壜�H������������,��q�|���,�)�u���s
�rw�ѵzT����N6��B񴦝Α�Ď�X
���L��K�8$k�����X �۱.pv�R�yZ�� +y bσ�����s���<O�\��=Y�+�Z��eR���ٻ�"��8�9��qD =]��5�J��3M���w~6�Ne(G~��9�����N�NIV2� �໺m<�zօ��6dHN=�ꅡ@�|	�4{�F]�D7�����e6�ޟ)��x�tֹ���VA���q9��-��;j|d�p�����ϟs�jP��j\���W��2f�B���2�WƨÃ�l�w�.�üj����v�i��+ˀ��͓ɵ}��Z�	
Z� >�	���d4tǢQ�'Y�%29]�(�#�]�׎xLA�ć0�ġD߱c�vyK���b�R��)��	qQB�hg_�|�=��yR���ƙx�ߌj1�YZX��;�ݸ��ؿI�t�)��eR�s �O'��V석�@���<;԰&s��~+;r��{�D�Mpre�M󂛒Y��A�M��1�{/"k���A��Db�W�p��=��
}��F�ȭ�����G��h���oW%�Z���z���}Ώ<Sx�k���	�\�&���3���B���p?%�\S%�o��Uy��������|4�i w=��A,�U�)���<Vo��8jA"m|�������e+������K它�mr����Sϯ��VS9\���^�^p".���ς3ߑ��0����<km�-8m'̚�o���E6��38dq�3y��յ�B{e�@#e��G����_���W>1`���m��R���w�C��*�t7K�	�ฺ�}5� �ԿV���t�!��re�|�aZ}}Q'�_����!<)�ʣ�)X7�����1��`�����dִ��������� }���M��B^��Y������Γ"n�v�d}hk8��8�s��� ]@���3�������~�fw���B�=�;[[����]��4Z8責�X�U��K��J��⛞�'j�<�+��M&���!�
�^�IO���X=\��v�i@+�պ�`m�h��?��(�����r�`�0B�,�粸11^��̩Ș�T�j��Ď�����Bw��ROt����x:_a��ϳ�P�Pcw~U���O>3���珄�h���VO �2�NK���B�P]3cWԨ�U-���U�e_b�\���_�!���;k����2ױCN�gs_\�*O̔����o���&�7H0��0 6k����!@�k�I0c�!��"�o�$c)���R%; �D�}�3>�C�[�IԨ������5C��D1F�Vc$e��G��_���/Ӽ$�/H�r�3�<�ίަ\֜�ֆ?����W,p����=S	C*�P�c����X���N�r�b�,��"�ktꡫ͇G0S��<>k��pL���yD���Ln��ӽV�����2)�Ev^ө�CVE��'���G���촙#�,n���扼�ϑ�Y�+h�{̮UȣEd �U��
y ��?�o'���8�0ee��'�Pda�x��H�Y�G�6�Ӿ��č\R�VÍKr\�U����2XW��w��Vcɍ�՟g�WT�8ί�T9q�¬�X���N��ڧ|v�j4���L�;���6�}�U@�OԨ��Dky�A�0��N�d|KX���ů�i�ֺ�`�mj�+p���O#��x_z���0L}W����I/U���7�79�ms����p��W]���~�sb�,x?p��u��i�M���������
�2��Aѡ��bP��7�I�=nl��'��3"�E��E�Ș����J��gkpUj�X��b�2�x>^�)�_b�E������8��{B�qZ��~v��� ҨD�X��NE�K��������S��׬��u��}{�d��󂦞����@�l�K��Z�����>��?�.?r��H��$��o��.�|�`q�j���X<pբ���qǍь9���U�Mw�(UOAlP�ER��+ol�
�����iiZ�MX"Ԧ�e�F帯�pQD�q�G짒��=���,Qӛ�d�8,��=�?��~������8|�vhݖ٥��ł&�����.�A��!�qK�F_&�B}�c��%��D�'R�3�;|���uu��p̺3��v������Ox��%�s�ҳ�/�J��w�_\���ek�e�#Bݪ��o�#_l�16�F���X9�ݮ�:v�6#�?�_�� ���Jݖ��K�����rr�ª��-r���N]�e@��Ւ�LexR����I���. ?���$]�E5�^����;(k�U`m��i�8n1��V�L�9A����J8M�#�H��������ʊ��+g5)dgp�qe׿����1��j�Q���8��=.�,u? �cPK����r���#��� ~�S�r��G�(��� !P������g�=�r�d�1�,!o�Co�/|��'���3�@L~@y�B:��&�fr��d��	��v9��Yx@j�����`����9��*�y)G�֜lg��̧N�2�6�T����{^�Q�w(~.��[�i�V����1������B�Tʨ�U#�D5�~������g�Y��>�bz�R�!�6U?K;d��~�5�#I�bf�~ژ����b3�j��o�E[$3�
�^���q���v6㥌+�m�N�ٔ�u".�k�/J�H�zO��wh
��H�
N�?�^��.��	�ܥ�k6fΪ���Q��7^�a��6��BS�4�����?�p�y@Cp� �� A�sf4�.��O(ם�� �D�����7<i�̏s���E[��Q@3�N�����T�?�x�Z{���[��3���Œ+1��{��ij�B\8c�L
�.�%�2��j�V��[߽�~Dx�P��)xF*������i �}~��=21~�=�˹+��5"ѭ������;��"����>��y'�DZ��A�D�M�q�1Be` n�/W���R�5�J�М�X!���T�Ra�4Ѻx��ꓥŬ�,�����F�/�E�!��w��[�u��a�x<�N���a3�Q�AE����{�t����w#��w����ko�G�.��� ����������!xX�-��ͽ�����;g��9�3�U�UO=5�{�wz9ƀ5'�
�+�zR�`{Y�v�<�4��7�*^O�&# E����j"�}NSQf�Th|I��1q!�z��}X�j��%���H�u_89yP>��ф��Z'��n;���
"���ï�c��D�xx?F�~����p߬�����ګ0�ɕ5|�cڎ/������G��^�H��Gߡ��YR��qc�F�)�a@�@=c1�8E���A.I5�����J	DD>�Τ�^��ly��xJ�;)���n��h�=�D�6J�s��@�lW���'&eeT��+T��#{��	��a�V�M��.�Մ�����j�~���-b}��GH�0�xv󙽦��I��h����O�t[x�&���9��,�%��x�®�"�~���{��H��o#�ѣ�,4�z�"]k�D%e!�7�_��^
5��)��SOR���J�C��p�7j�.~��Aɠι���8V���_Á^]u�������b��<v�3I���9�#���\w1n�0��vj��t��~
���u��c�tj%��TH7��c4E�/�M@�&���E��a�V5{�9ts���3H�քb��I
`�Ĥ�7k��*�5НV�)+(��k�*ѱ��t�ҽ���֛�w�׏K�RTt�u �y1S�\*��v6�@���&դ�c�~�漕�/��*c��v9*%�*�p̋�mQh|��	���3~�Z���`��Q�⒗��G�W�����D� �cHh0����0�^�;���I�y6�C5�dL�����Y�����I����y��7�}[Тj|<޶��;M5�a��~�Ѓ"���o���.+ "~��&�ξ����NF3v��]R��0�n�H.��Nl�}�����{q�Y�%�ycJձF	$L�v��]}�ԥ�����,�-[D4V��	�j��E����ku�\��n��hf[ڞ���:������]��<�\�)<n��B2}�d�#�2��/�$eH�u��ȡ�����r&8��ʖd��������Q�Q@_�f"�".�Z��$(!���2�H�N�ܣ��|}b���s����K^��
J�t��Ũ��,B���pXo1� ��SNѵU���{��]洝��hV ��~������k��c�r=F������.z��,az�|��'�k�Z���'l���
���	�Eq�:j�	�.�l����-=����� F�����>���fF�w�2�d��M��[� =��Z� ����V�K/e��IPd-���z�좕�N�\ű*ш&�̘N�ܓ���o��"I��N�'��NKe�Y���FkWb��F�������ܷz��9�����߇}�(P+2�9��4:pe�a�|r�]���;b=�X)���&�;T\
���E	R�;qt�	"�K��B?/ ��!���-9|s�\���'dK^�vآ�Y9�A��2͵�dtFN%H��^̝�|�����.�IhT=��/"+�F��r���x}h����2sZo���N�ϦfO��EU]ŴuĸŽ��1p��HZ����.�R�9�=�giA�jC��~!Ti�Gf;���fw�Ǽ�Á�	ϐB�!��'�:r��gH�L���G�X!3 �ct�s�2�Έ��k��~7I�8��-
��De��t��k�S�}�&I ��ɩ�V8��d�ЁI�s�Υ1�x�\ J�Ó�Mŋ�*"�hc㢟�	t i|+��"-&�;b�v#�d�x�`�*�\���5umw���_��WŊc8�H�h.f���>��ަ�ҝ�Dn�c ~."�������L@����%t��V����Y��i�3mtϼL2�&7`y�%NlS�����S�ei���j&��-1��i5!kTZ��Kz���[�"��^Yף�]�S�M�^��E��#�Ǌ>X��<	��Ϫ=�!�6��"�!�n@��m��,�6ROW�&�8�'����3l�yˊI�}]�2A!��+�[�e�54��[%�q������-�+��[�lg�5��(ew'�Ѱ`�qF,��l�l&���[�L�Q�����d�귗 ���IӉP�'�TX8�&ކȥ=�p��"�X� ʬnUE	�cl��m��B�L�l�(� ���wP��}e	�9WJu�֟��?�~{q�C��Y5��V�H��$f�?�gD����3��Mߥ6��&�Յ͎�܏m��b5��y"���h�8A��;���������u��x����-�i��WI�I�"*�3�P�(`-��g"�;��@3���\�=X�>���cB�U��X�3��N�9Nb�,��(�/��z� [ط7=���I�U�vrq1h.㸵��(����w0�d�]�/1I�;]wW������Jp��1A;&�زN谳����j�"�V~I+V���X�2��������X�ҙ @�s/2c�����6zh�&Q��(JƐw���7x��F��Z��]{I���sfxQ��)�s�G1zY	�ʉ˼���戔L�G�Z.cJ�[=+	u-N��L�A��ߞm�/ݝ����VZgJ*4���)�b��]�j�
me?tU��!B��C�B*&�O���H�x�� ����*��=ƀUӽy�<�w"5��&Q�a-r�`�I�vr����ɖœ�z��:�л)���!�w{�\AD�yq��/��
�U��^!9n�=wv���{�~���'�cMb���"j����(	},Tta�S�SĒ@��&#*F+J����e+~h�?�Z5\q95��¯�ە��:�q~]��O�~a��3�0����\��	2$x���+�R�U��X��V"*���u]>�
{�������3ZEr�@���kj�@��f�{c/���Q��K*�l��$Yʎ�����t�2�	��d�ȗ��͐w��:��z�	���ڿ0���s]�ڂ#������#�C%O6.�n؜���j닔c��o��;�+:mR�E�� ���8n����۶O���}G��#��Q!��ؽ�Q�����u�y��<��X@��T$cy륜�	�	����يz�����'u(Sڼ��a!�?FX[o�Li��h�X�9�%
���s�H����m=ӣ��6 qY�2��`ٷ����������h\��]
%&�J{�d��0ӯ���Z��~I*=-��!%� �y�qS$
�v�ƎP�ܲ�<�e~E:�~�P$(�٠�C(�R��g��d'���[��}*��ې%o:Q_z���|NH�����	����f�9�o7�M�����l�#�<J����5��֞1Ѩk��6�L��i7Ǽ�f�Dd���z�p�{cƅWQ�z6Y�t��?<)���2��^p��ڈ�*�N9N�M�C-�n��E��z�r��6�)!5�TYc�GՌ��B��x��ӗU���F��ĥ/�n[o��tD�#'#:�2�5�>8!*�O{}��ѭB�j������P�ɨl<yڜ k�L��N�TV�,�Niz^��x�_S .��n��7�q�V�V�>��,E�+��y�f�nZ?".d	P��^/�RH@�l� '��;�ʢ*Ey��}�-����Š���3Y�����n t6̐����Ҭj�IQ~e{X�^�g����k���
�tԧ���X*������;��wK;��A~�Jĥ!�k���xnA�@�5���iIǭM�1��Õlj9�[UR��z�s~�G{V&��O�d.�T�b�i�RE������߃�\�A�]Kx��SJ�wE:�l�W����[�X���Jd�'mmI�Z����; ���ZQbc\��I?���죑Ѧ���j�I����Ҳ4~��~�{$���<�_&�T�kw*<<��t�R�^���.n����<#< �?������\.�t����<o8�߻�l��Δ1OE�XN��R�9m�� qusl�蘭/V�;��a����S��z��*�Ё�l°�J�Q�aw�٦�?�y�u,�IԱ��6!C�_�s���M���}���No,������J7I&�}����)���������O�ך�z{{���uR����!J�[�Ҝy��z^�+|x�F9�^���yX�H�T�)$�s�S}"��b&p��)N��[��O[5��U�����A�!!q�7Β�$Yܐ��ntr�6�/~KNP��f�N�r��_at%BB84�ar-�h�s\h+	��� ���x�b� ULm�����5}o&�}�0���V���iQd����**��x�ՖD�D�)9�k�*���'���/\�a�DB��)D��a4ro@Cvd�)�=���k)� �LeL��)2�rȌtO෯	S�����^q���gb"/���0�����PV�w�I P��sӹ�͝�{b��*A���iWSj��c��������?���Q��9ƺ�;C��|E\R�?G�W��_?���`ö�P�J#�=�#V�x�n�Z0��A�B���e-|7�/�bz��s:�n�~1���gZ!��e��z����|�2絧����ԡ@���Ũ��*��⢤F���Ϯ-���)w�Y�d�pm��J�Y%�b�Y�����4_�d̸!�t�kf�.ۣ-������j����ķ� �X<X��W#��== ����%X@�d?t	]�"Ԓ�IcGȝ,M��A,�m#�Rfʅev��sPPl�PE�T�I�C��O�B%V��s���ӱ�/z��:����kX��kQ����c���ɹ����$������׭��{<h���G���yi�� 1I��~�F���䄔<UtK���?Z��r��fu����Т�_�S'�g��B����:*/o�l�r�0B��9"P�Q�N{)���?�l0�u��"�j~w����Xnnnbq��@��uA��"耞!�o�XN`�+0N�^\�hӄ2�`����)f����m_�S�I|8�椆�xԖ��@C�'8Xأńu��@�^Y��%|+��g[���3M�NU�jئ�t:{]�2i&�\Y�4�xK�ēf��I�@R��t
���ER��o0���|�e )� �C0�P|��G������$$<$o�Q�Ż�E��1ƅ��J�ot���T-���G�:�m[0��`��~I���vw;�ë�`K��W�6�$� ���q�tNӢ���ǉ*O��DS��2H+��q�Њs�a
p����-rQG}2)Џ��{ҷ�~���oΕ�t�Ǜs���:�\�qt(�_�~8�~�7�ě������c���G#� ��	H� ���K#������2�d�Uu�����B�/�?�ʣʫ��p߇\bY�9>�a�LF1�n�BhbSڄ>E�RQs3��Wt!ER�$�D����p�ˍ�$s����n̙�\�G�$��͠�#�Grɽ�P�!ִ�J��ѝFN��@�p�0�Ͽ*CϽ։�g�ނ���v��<��gP��	xs{����fo��Hl�A qsޑ9fٙ�仙
��׏�
��:�	���7����$t�~��KF>7�?����H�Zmre�_�0n���T�r�P!��XS�Tu|�ݵ2ͩ���P�><9��Ka$vb�!̯��.Jjj#���Z�A��D[�X�����j=���ƀ+�-�����U��
���Wdܨ}�6�5Bbb	�{9T4�8Kr����۹<5J���^�q�2�<�LЎ��Oc2-{��0�p)��'O\�(l(�i�N)7��Fyd��ۯ��OCeP'm�����[�	�dD�t�:
#: 2����/�p(�*�&^����x����� �R������IX���.Ѹ!���v2����I�/�!ſ��&�+u2�ϳ7]#PB��6߲�Tt-T�K{U?,to�L��P�����;׎�R��Ԡ\�r"�Pn�<��%�"���R���d& fRɫ�#�\��2��Nk��BGd�:�)8!���+IY.r�c�Ǿ��L���S����/e�*hI�H�U��b� B&;(ӳs��M�7���,�V�V�����b�h:!>���2���Ԋ�-���LpD��S�H
�r�H���V'<Sp\<ɣ�-� 9H��³dUck���
�W�M�p����<���9c�a�d0w!_�B�_)aB˖$��o^�(��E+ۙ<��I��IH����YwV~�K�@@5�	r�1gH!:�%�d���ʀ�^�L/�h)�
�� U��5UMj;N���e���Mo�}��Ao��]x���~
��	,���o�Hv4xy\ԡ�I79_B]8e4��`��D�G����,v,�B��������s+йu�[a6'|?�I&�����l���8=��5�܇s6��	�y^�b�U��Z4���
t���yytleb�-�
 ��=��̅�T���x���M8�~>�;.P�w��9u�]��ӵ4��7K���y[`Vx�f��Z//��Y?�E�N$j��m�y�!�!�FUMF��ݩ�KX����lĭ�00�7,��^()�<9�L���bJ͗6nbee�>���HŜ+F�tCl�q��rţ�KrV�X�ۙ�7O�Ã�]���^2(���LR��.'�����!N7&�Z��0��s+~f!��ވLi��M&'�����a\S�5�3++5]w�P@�@�T��z��&u�(_r�H�q��~w�u����sZ'C$r|mb���J�T�#��4r�<C�b����IQaIQ%f��rf"K�%���l�ħ�j+)�)aե�
gp��YB����dr$r2~�.���Z���� "��;�6����@��o<�u�61�~b��q8�s\����w]����G���@2�%�(��}��V;>G���;��m=Vc��{�?��J��W��ZPo�d\����,��m=i�d:(x
8uڱ��0�H����gʤ��耥�?�j����g��w�p����������<#\6�����{�Utr��V��J(��#H��l���^���N����4\ΫWd�p������26�MZ�b�oK䋭������9j��kf4��'�Ϛ�\ٟ�Ƨ]�ܓ���l��t�ʚʥ`��~y��K f�����Ï����W���>h4 �7ig���wz�>R���e�
a�K� ���;:ɲБ-��sN�-�Q��!)Tp8r2雜�Y���5yHk��f�{P���&6�-J���׶��
J����']T��!bO�!�()��o�epo[DH��頂���a����>��১�����<���<�e�j|��J���^hΐsw�jV�P_H���&�H� �=z �v���2�Đ5�R���/�^8�G9��>?�K'�``��.�n??�M��w��I��5�&o�*,�����.�����`I��@����/g���m��',T'�`��=��D@��#���+�L��hI����yޞKD�s~���'�x���@y�Cz@u����^-,�L+Ĵ�rm{s����;Ԅ�"��,�t�7���ű�|@^�v���5�t�Ci6������Ӂ�%Nv�	0�H�4z�e٫ /����8��"�E?�P¹�Aa����u+�L;�_�*��DI��D���W1�])2쭒�ESn���ěs�W7 �!�B5��M�H�2-��<ɦ�G"A�GH�����"T0��r4��ċe{Ъ�g�����/�e|�\Bԙ�-FUx��Z�A����tmĊ�G���/0C`Ǡ�7W��T�Zk�+�N}o�?�Z�0NIz���":_��D�<:}�Z�	��+:W>��_���+7`�}�ъt�"0�m���Ր�
n��^�{q�s��)�u����(�?s��^v�Q�W�w:���t��Np��"W�Pe�Ė�JU�p�nx<q�����ʛ�(�Ʃ���b�!qn�ǃVK�OJ:�� �8����bA2C4i��҉E��k�Կ}�J:m]����W|���;%��i���bN�5y���L9�/���qd�r��8P]�>�r��67P�V'�;|%rMv�)r��!-��"�!`Zj	k�r��1y��s}�b\�g��S�p��2
�>E�n�� Y]�p����I1y�A��8���]���⾻�~�����_��>���o�n���_z��.�5K@3i�+���iJn�bs�5����.��ʙ�	�)v��!��<���>�e��[�|f	I>��z�)��Bl/>���Y�GW����w����̓��%A��ia�H���8����kT�6t6}��sА7�,*6	���e2��$� e�����WL��c/���fgj�da���ͼrA�:=߾ȫ��/�|�L����G�����YB��2���5��
I0>6�f��MK $mӠ	��Hi�F�*&u���6��ʄ�Df3h0uV�CYJ&�!�9��i����2�m��a�'�\a���?�SSk$0�h,���hv�[u�3�P0s�˅3q[���d��k������x�2N���hLZ:*Ps�!δ�Q�9�Fm�/U!�^\�.n,9���	�kR�EԣW��vy�a����>~��Dn�]��'�n�x�``��޷����P?�=�In��kH@;�Itm�P����dT�_���O�<?܏� �Ǝ ��tن��>�����t�>�|���On�}����](��]�^�!���Ho���Y�Y�>��|�6ْroixO��4΋}��I���:"Qk�
�ti%�c�4�d�e]<�k���>Wc���$5ݐ7�B���?�R��K�WR%�8)#ƕG�/;�#W�[��/'
�hSWE0\*f�Fkl����jM�fr�c��8d7ʇȚ�RkH�]»N��!�����7#Q�aϑ����r����ՋV2��!��5�vq�޻���pOU`���h���������	}�$W��L��W��	�2���lO׬�ɞ�g�E�7F ��"W-,�f�/D\�������FyrE���Yl8.�>|ivݮ�	�������`��C�3,|������}��:���|(b<%�.��&"�0��_�.I&O�o�ު%W��­B���˕��Q8��z��A2���j��PP���(e����WDo��!�Aa���л�� �qi۶)/���	&<�QJg��Gu���UK���@��"�]�Ԏ��L����*T]�:�+!s�M�Z��O�����t�o�+7Z}w�yhp_̖�]7\�p��d�Nz����6Z�X��7��f��zN�Oǒ�DP�X�r�>+����c2����榧�ű��G���v�q��S���~<�ag��f&��
��V39ߣ1�Y�	�o.���N���r�;~� )밑��D��o.�:���g)5�֩f~�i��
���|�Y����uEB�|>%�Ҳ%����(�2<���	E��q�L�������q�S�v�ͱ�;��Q�rR���㢛=JR.�T�/�:�������!��c�>�ڗq�>a!�C����D"ޔ�ڌ��xJ�`�?B)�9�=��^
�]yɎX�u���Q��h�y��~'�7�����8oϠ_�I�jT^���{�o1���Ip4�����Ӑ��$>��u�[^wH�
;z/1RvL���"O�ЫC�0�L�r�'�r\w��8�<{$ĵ� :�|�}9��y؋�c]b�~5����_�G�Y�U�^�t^�"e�h��C�Z�������do��ŨW:;OT� ���G2�(��koJ�E�
��D��nw"��dP� F�P�j�?������pbF�g��a'���$����@H6%ca��⡅!r���M���߇�a��7�j�Ce7�;�!*�Ur�`�(�T�, ���ыjyvȈCxp����� ��������;�	X�K�<r�o�����7���n�ӓE������ˎ���`Zl>Ro)��[�',Uk��&�b�ܝ_��b�a�n�Gz��4�~-���W�Y�%Y�y���C:��c��}����x;������2Iw���E:�}��
������AWLC�,��C�����wU ^�*7.?,�%�/����9-��Ӛ=��vD4�;���ᘒ19���*N�C	�^m��Qé��vO�!�!S¶=G\��D\��M�f$o�^x-�{�|�L�l	������R����pщ�/8�Z�W��1k��/��qu�b�r#�9�&��SC�E�/�W�� �垤\�λ�s�f��1=���P^[6#rZH �J���?&T��lO�:H�&�,�cY�3��j=�"w��k̌�*h�=�4��>��Ӻ�I�G������Њ�f{J���eP�M��p�3^^�U�+:�Z��x8��l����9e���Y��� ͓g��W&�����4���+����-<�d���e)[P���'�+���)s��)����X _O�ayA���#��O���H�q�l�`f��u�q��L�����@�j�U�^y�-/q���J+k�<N��h����M��4l��B.0�%��bUz�~>'�=�]=��h7J)�za���N�A��
�t��U
;;��T5A� �=��$i��.��B�[K��2�&�u�s�P=2~z�<$;N��m��B�ݎ���	H��!76�w1$���?"�]�?�[�/a���.V6�y���� �;������ �4���D�M�p���_qe>��~P#Q��CE\`?Д�w��#����Mv��N��gc��Ƀo�i뵚bZ�_p�y&[�(�#5�:��}u��	�S�c3G��iW%M�7�H_���D.9]�;|~���M$ ��7���h���{"�}q���e�-�5��*�����$&�9+>ynq�2�BM-��mP�1����{��?�=�,�0���lXwl�T��������iҡ��<����z������V�p�j�#�=���<�MaޜA� ����az�i�i���i�3,�<�~q5�}�AZ��l���b��-iz�N���\�����G����sXÓ�S�Z����1�?iI�����}��}����j�*����L�ڊ���'E�/�-�P�"xY'��]���W��u.g�b��|R�ݨ����|��Cͦ�q��8�z�TL��_��"qt�pٖ4���^e��x��G1��(7S�R�{��{�jgv%��"�c=�b����SBʵ��b�:5�6�	�?��V��+L2{�=�X\�9��9�o���a�pr��+�~{���^����߰�1��Ѯθ�}�@�����N]��I�>�p��T?�_<��������fe�lU4����Y(6�a��5��/1u�\�1�~%�a��&}TmT�pڗ�Ğ�-8�:���1��'t�K� \P�'��3Ol>Ѥ�Q۳����r0��3��0V��������	�	��,�yqF�ɣ'��యm�.�����R�^Sk�3d2�GZ�
��`�#[��}�=�\�H ���,/�dD��ň�-�:5��:Uc�l���ǧy�2òi�����O1��[�X@i���̲��q2 �=���E��|�'�<1(���l����Rmy��'�^z��^�6�����:�r1��2��.�BN���p1��.>R}|�ک�9>n3�t3�K�]8��E�@��QB^��Dxpu�À<��8Y{3_��ft����cp.	o�C�'׃Ԕ�Ka���Z&�OԒUPR���&#�t�V��� T6Bg�VT1����-pmh�u�+��	p�"�A�3O�'���q���&_K�5\z�����B�cZ�6��eSLr?P�Q��4�6j����DƆ,�Y��}�#���������y�ޚ�:�̄�?�6���.�o���yt����ɲH8��|ln����W� �^�ij����� '~��x�7��*tqN�JfN _f��Ӭ(�	,�>��1����=�B�C�յ�<�tkH��p!C���.]ш<��?��$r���"F�a�$rS�d4��n��w����Sj1�������+�}��;Ш{�o��
�0U���s��x+RZ�XY,��5��i�T�xU�Pb�)�\�h�cTmj��6	m�i�8�|��c@~uD�J/�p�@�&�	����.���"� ԛlG��n��{N�" �`ʢޯ�"����#}_�H��&?wGU�>z��B�������SR��&XNr��ZR��p1}���~�)��&Г��G�C�)uJ�v�tI;�)�y�TP!�
*�¿?D3N"����v8�nۆ#�|��YEGG�yoT3������@�I�/���ˎn9w�_yF�:I ˁHF�ɲERc����I��8 ?���EV目�@�La���S��,(���v��J�!~��$���/
�;�K�l��l�N�@ٵ�(`�	Қ7���-֢t��]#6�oW�ψ��SN����g!�d[������,MD�8oCd��B	��x_�	��0���bU��'����=�Qߝ����Έ��2��)N''K��{n]��A6]�h��lqLXU.�?��P�>�zm�m6C��;�˓"q?�)]Tp�xP�p�.�@C�bF�>5�-��*<���x�� !$������I�������)m_�;���X��:>��~tnG���A������~=�1�ZL�p.{���S Lj܉�������J�e�S�*��a����D�Ad96�F8O������/֙�eN��w�$
�O��»#�[zK?�r�� B\���p��������nvx���>�"�ދ��c��'1���"9˖6yc������n���x���|4�,��g��UʯZ!W:GU�ںެf$�J@j9W˨���)�v�"=%��Ԗ3zL�x�;l��0wO�H�L[�S(�7�*���{N�i��+CD�ۊ���ㆃ����؞�Ż|x��������;,DDN�<�� *�	��BP�1S T4���e-E�-[b#?�1�6��(�#WR����^4���b@�C��Fm�d�[<�ĥթC-UKdH�KJ���'��Ճ,3l��!��co���C|��AW�*���1��뛒6��)R0�)�\�XK4�!j�<�$V$cQ��e;�;�-P��M�Y6	��	M��F�7O���
W���5�[�����k!�tB��������c�;��!��r�v�����V(F�>����uI*i�=1ک��>:g�g�?�ݟ�y����Ʉ�PD>�@,>�p�8��܇#�9��3e�a>r��.&�NP	ktw�#����%�\x)�ՙ]_���HA�O�}�!�@��Jk����8[�/��Kez�g��v��*Tx����9w��/�}����-ꇹ�,����:�FE�!�z�w�y�)�@�x:n ���܎���/������M^��oãG�����?g�����9���[o���#v�:aZ. d"�!�$:Z4ᓤ���(��N�ɠb���sPƐ`�4��_����+�z\<��~�y�9˖�wYvf�:������$��4K���p¥�!K{��T�!��+{#CL?�ps!
��<��o�]א���s)Q��c"��on��Ҙ��L����!A�!�?P�\�m�C�)J�#���2c�y=����C޾��
49�O�P��]S&�#.��
���*�>xM�O@�/)���u�\Xj�e�u~��.��l��\�!`�����>)N�|Z�ac5��=$e�gG����|o��7Rt������PX�-xp���xÚ���Ư��I���\��+`�bB��*V@��F����FS�����.��K���z��Q����',7���MC0� ���������'n6���×h7����j��� �'_>����"�L�N������(����Qf7ï�ߊ"Fu���sL�4��H�ơBfd?�.4<�N��M������D� )+'�Fp��N�� ���`4;f+;�L���l��C�݇{y-E|Ι�p�?�L�B����O$�s�ř�_�ۘF`�]�.�� *^(��c��hf��C�Bd� ���05 H����CC��6)<1��� x�}��U����_[$S ���R���!QzJ�U���Z��v��9�S|=9 ���F��it�Y|`����{�+�E�J�B2�i��	{!�
uVL[��W-��f���X�43U��0:�@m�S�m<�2[aE�?W!U�r�u�۩��"�?��,� ��Z��S�xl�Dm���@C���1S��طM���t�0�l��Z�R��Ц������uf��IU�~V��\J4?�����&U���fr�����2�9�.�[�k���B2�#�+�Y���E��rx (�޸�m��3��4
�i��q6�0a�6�\����[�B��*�P�����:)��[�!i>�ã��/����B�_��Xlf��b�Ji���`�<_,H� U��-6�&%�9��y��P�x�S�
�f�}�TRLcl,k�*�n����~8��H�_g$���x�� ';�Z'{��2<�H�;-2*���h�-����=v_p)���c`�u`<����m��p�K��@~���4A�����^J��4�U�~v�`Q��PxWbR�mK=�� ��9oRA,îJ(�,ܱ���W����FF�c��@K֨����ql�!o}�2)�Ps(��?�uqv���^���3���؈���@��wN����@+e�Zlvܳ!�
BIͧފz����}i��� �I��
 ��� ��}��$ι�Ko���	�J��[��W>1	I�����~ǩA�3U��z2KvE��F+�2Y�aǙ��	��f�u���y/��O�YKZ�����f�d��'��p�]�N�s3���v�ԞYՋ����N�vw��n	��n��=��u]�5>�i\��V^V����LŊ��WH$��ٝ�O�<��k�7�Ӗ��D��d0Е���.���o,���!�8���q��^u���x}�ﵿ����Ns����:�&�G��q�1e8(�6Q����^Q��[��i�>�I����'�ȑ܆s�QO���m�	�i1�mz$q�"��|�h=F��j��M<ᛯ�<(��rt �32$��Rx�WfQ��n���_�[:�Z�Hܕ��?�QW��\uz��-{������"�n��k(�߽�_p�|��O!��� �͐���3G��ei'^���S����l~�lEL���t��b�}�xna�lH��}�r�����d������\8�A�7,�`�j+����WRO�M�P�.d���Ɲ^3b�-Ư�ך�ڧ�zVr��$���ﶃ[��#^m��BN�;/�x��Z��a�x�:;�t�^4A/����1hD&��Y��ux����x��.�^\�N%yG�s�"J0�C���b��p��!������[\�#��j�r��e�=edB��;�	�T�ᑥ�XK��sWK3��웲l�����|�6�W�c4�P/�,���5t���woޗ9�ο��8���>�~U,{s��l���F���dO\8�����^oȸ=?���)�"^��k�f��L�'!���>�w]eo�K���N�P\�,���Pl�*;�kɧ�o�l� �}�${�Q���������Ex�s�ayW����u�Ũ������Z�<������1B�����5��|�͵��un�a���-��/��*=�͔�������אּ� ���|#p��Z�*cP�&Cs���/ٯ���3�����#�S�O�eؗ�E��#�t��������	~o�3��33Kj��A/�O��Ͱ�yt���v�8Z�.*�	0Ԉ��Pg�=j�^qd+�x
�n�G�V7:_\�\Z5�%5���O�@�6sh�\�f�nK���P�)Q)`�ۋ���y���x���J�8��t<��\����q}P4���*՚��u-��nH�~�A,��H��E�^�U���I�T����.���_��ӎ��ֺ/���I�=Mn�)7]�LJ��p���������q9�ƨ���?�]�+�j��=(�ê�V\����b&}�;hK��O�s�f�B:L��d0gX����,D'���3M֜?T3�UwTlx8U�� 7��E�8����yTʽZT1禍����[5�[x�f��,�K<7v͋3��)]�)%�U�u��<�B�}����o�o7=t�n��rs��0���^3|_�-���%͈<�>Ѡ^������H�`���e�ʘI��/��^%����R��>��,X����p��1��k5���?�#���ֵ�(���UhL�~�-�z2���a ��4q:����o��9i���ˤ�0��,�ȩMU}��D7(�<�U9�־Fx]w��L��Q2��/]��gf�/�~�6��c֖X�K\�SyQu�B(�yQ�q��t���2UZe��ƿ]��?�Z�WV�Z�e���,�ˣ6[j��bh�d����4W��)�2Q��,�rS|[�P�E��bB��$d*����������s���������Ց����NV}��\��_ّ�"79nZH�B6?h-��nIVݗW�q10_�� �H:�8�h����L_���C���Ӕ�\��wϞ���d�q���UT�������K~�R'�>Ǜ׭9A:;Ƀ�L�����4�`]ꬒ�7�]�v����Ndg�<*Z�-�'�����ּ ~W��f=0���lW$��D���(D��u��SIP���hX�E���IX
�y��6�F���n���;���oH�Y�v���	U���~��D�)�Ut��X����.�Wf�aߜ�p���e�v�{a�}�������GG�u���b�Gl4���)<d8/�}$�V\O��pO�Y���U,�ᨦ�H'�Rp�%1�����~?v���WC�y�3-4���<�v�Ea�ɸ,r\Vҳ��/{8Q��'�0�S��X��k!(�u���?�Yq�v�(s�Ax&���bӹ�B`��r�yK� �� X��R��9R���-���x2��G�B�}�h����<Mil��|:�)P=1�֛�<|ǛeWY/���=��iI?E� ��];�<�ܭ�C����DJ'[����s��K��)�yDoG���L��]Oei�9,7���̪h�7���Ԍ���F�!�C?4���Nd����a�ۏgyZ�aˆ'�˰�����Hu$���˓�0%5-ZH��E�t L����^��U�t1���&7��'7������ݫ�Ϳ�$d)���_2��\"z�l V�iMn����H�.D�:�5sӶ-�Y�� ���\�ы��B�u�*����)��a��V�r�5���1�?!L��)��dFIE��쒑k���ע�!zz������Ul'.f,���N0Cz��` �"����{�T���	'b��C.>�r�΃(}M�7n	6ظ�[����w�<3\goSEc��C��e1yo$��opk7�+�70،��d���>"��3�&k���6�W��o�O'����
�v�k�~�y������`������N��O��%�'�J!�:��;�bMk��Q��m� ӊ���w���ٺ���m��m,<_�ò�.�5������$u�l�T1A��FsoV�؉��\_0=�$���YL)L�2/v��k��g]Ƨ�`ҍ�����w�y���̙���q���ud���O�C��\{C����U�j�}@N�=�t�a11(\����	������ݹ���E��j��:MX����{�ȥ��[�d{*GD�w���%�-)�+�A�^j"(7��y�+!�j��W\���{�U� ��t'��m�2�5�݄��B4}y=�`�up:�a�N��J���U�#�jD�#7)en�6�e+s%�ǫ�}��cQ��Xh�z�S�_M!66�(��8�?1?&=�^�%��/C�7R�\��e�_j���9bZ�1TWP�Ȯ���qV�J�����4܊�AGG��r �k��~�M���ɍ���veko$W�xMH�}ɼu%�o�q��S��ۡu
�����~=j�>��!\L�[S���e(�NX0�^_3���+V��]{T�{׳���Sr�}�QF��C�+�^9 �'(7��1e`YP�W�A��/8��,�`�K G�n��'��ş&<�>�m��߬����M
\h�e�o�H��@h������PK   %��X�"�Q  �     jsons/user_defined.json�]�n#7�~��,2S����l��������`�x�֮-9��F#����3�|�b��V:HPF�֭�C���<d�z��t��n���t����/qq3���<�c�ܬ\�ӛ�g�����+{U]�f�1.FWn����]����'�����:�lP�L��(��%&�9��$˹��
g~u=�����mY�a]�[�g��*�lo�bz�\����o��K�^!mmD��,���S���z�����l}�LhE2�*�]���<9M����ۋ���x:����_��˟��"|{=�������_f�������~:�_��<�d��?���wg��w��}�[��M^A�f/��r1��F��7�����e}%S&�>$�����7G3�a���ooߥu���v؎N� =�˛�����f�鍟/>k������&���/�������o�ꆾXS��t��7�h1����&߻���wJ�<aދ�^�at2]��tY��}6E�9I�t*(�(���p��m�Fq�-��\K�:�"CISY��"�,GJIF�����M+16�_?b�-[�w�79��k^��W��x>��2��!�A�{+2g�I'x1�^-G�S�m�B�W�n#M���F�}5�A�{|�|сO�ݤ|k�#�Wk�m���.3���$���n};/��=�t�G	��]��tWNtXi	�{%iR���Ik�+-X�J��tG^ti2��%�ơ�Ch�wO#쯷��fm��:�^]�*il/W�.�q����_�N@���������}��?���UG���9{v�J�/W��x`�����/��2��b>���=���C�-)0��)
��L"G@�c�������T�[7���"�����e|oGTH�D�Ե��Ae//�Nt��M�!� @���d-�1b@W�r��!*R�DTqM@�pB���4`���.��]�`�5yfY<���l����E��d�^�l2/^�=����!��)e;a[�(�={~������E��m޹���"P�"!��ˡ71�ڔ��}�ΠE�G��������y��&%ʺ�Qǰ�M9��vD��P���:4N�B(��G�� (��G�� (��G*�$#e�:�$+��&�$+��yF�&�Xa�'#�&�Xa�'yR�&�Xa�'yV�&�X!H�V�I+V� ��m�t���P����i�ɮ�Ɋ���瓣<t�x!41_�����Z��J���]�-|���j�懗P���B<R
/k��x��@\
/��y°��fJ�9���%©Bh<:�1��XK�+e]t!�~K�S�c�%���u#7IKiû�[�d)kD7r��,%��Fn���\Q�ȼe��M��Fn��BdӍ�2n���wC���D)4�n��R�n�+���!o��2�ι�&		)�=���&	.�����?S��!hDK����e�Z�����֢E�V�� 5�D��Pe���nD��PUj~p'Z�g��P�*\�(�
��v�V���D��v4W��a��&���Z�fK`�&3�"��5a��~�������H�X��d�a��b4�d2C1R�1��d���ю&ː���v4Y�ea�cRV6I��gG��X�Z�!դX�Z��Z�dX�Z�S�I��$*�g�T�_5jIT�Ϣ�&�jԒ���ZMvq\:��ɮ5lIT�h�&�ְ%Q���2�*�
-��WQT�7���(*�LgV�M�3+�
�&��E�|��Ɋ�BG�eXV
�
� ��t�:F}�D����L?Z���9�A����ِ,:0h�̊����`�q1:�����y��̫>�d�^u'/�4w#|���"2D*�D"TQ����DѢ���+E<��;ĕ�HSP��x&��v%/n���X+&�&�����u��r�o��*=6��C�SY/3u������ǚ?ۊ�L������z�$1�a�{�xB���{���I�1�����lZ�������]������z���|���-�e)%D�5�3GQT!�d��j�]ԡ��)��L�Cpc"<���1��M�Dw{o6c�[G�w9t��M���#��=:��P�(+�sY,/7��3�����^�����|��KiX6i=���!�/faU]��<'mp�0l�ȫ1r�z��*9�������>�<]|����F_A����j�iP�@P�Q$^I�PJ8j���i�:�3��c(QSj�}� �F��|�ћ����~�fi�7�z��c�|��g!��8k���{���y��^��,��0�?ʗ�	��.̻��c¥j��|���!����*�uW������T=}��I{��� \�7S��hm�0%�"��� ML�	-I����)^^�?n%���R&$�JI����X*���T�>�NV�hr>$菑#�h����@T!��I��kA�!+!8q/�vk�H�&P��	�����c��_�8����Td$2䅰�1���&k�<`��ɶ�$�As����(J"��dc|�꟔��!H�Wu���h���"��>�qW06�d�����j�5��ZY�u�@�xB�j�t�L�<��;U�\I���	�*�����q���`��ҁ�J�+�~��x�l����BP{�2���T�D��`Σ��g�fz�lL��(��)���T��u�2�y:	+�+Iy�E�N.+��ހX��g5CN2�����t�~S�6r&I�-��@�w1>�)��c7K��EE齟�B�)�JNҏ�a����#Ǻ��Y=��P�Bao9�������� ���pfg����+��{�� �	�{��˸xl�@����W� �i���?���5���~��Vu��f=D�4�VW..F�������}����Cq(�l=�̛hBD8
�ax�-w�2&V���0x��#a��G<���0x��#�Ky�7��n�\�g}Sƴ�H��V1 �E���`8)%br��R?�cT.�Ӵ�5r�}��^z/�!������&�� ���1Ø�)V�.)+J2�I�x��)T6�j�Z��G�ͽ���'̯��-fZ� o�L�2�j:�[i��C]�����c�\�K.�OFtt���f�z�6���w��[��=O��hC���O�#�Q1!�x�K��	�0��A=���#|�
���&Sw��vRb�9��]�
�,Q�����i��XM�\�z/n�1���/AV8��b�,�aq�;�R�#�cLh�����}>8d�U(�`L���?��jB�s�N36V��U��ќl�X�����ud۔)�6@��0��ɀ���[tm�{Y�8�aA���W����ff�\[`��� �ܨ#�0�e�c?k��-H�zY����쭕B�94�����Q[�S xjL��������?:6�6w��_���`:}���o����
�����t�?��B�ɵ����Yl9�`:fJcr((���m{M�O�>�t{�N˩(��#��v޼x��;M꛵����������j�P�7~�6�Es_�Ӧ:;z��;�tj]#̊�=�l���j�	M%09��7��?u�w��a1�!p��"�5�)$c��x�K�G����!@;���&9o-~?YCTA�VJrF�F#�M����!z��`��-����`�UF8����ْ<�і��(34 r,�h��ea��5eH�?$��r�Q�6	���#-GZ%��+J�S�N&�Mc��"rt=��q{��P��m!�F*���F��J�a�Q��Y�VŌ%� K$C\P�Z����j� a�`ҏ��P��%mO�@;�_J3���a ;$���-J���y!]�-L;��N��O�h�TQP��^�PѲ?�Y�5#����~��mlFNݿ�{�gӿ�����8-�����㨅�����`�EC�],t��"�K��0��Ad2O�;�|n;�}�Zt �v��.&:��n;����o�mQ�dR��5���j����jߜE<�J�W�h���'���}�5�A�~��/f:�����P&�1!��E��4�4D���~)�J�"�J�X�сlQ1ʙ��Z��b�ʩ瘵i�Q�>n��CM�8�-������ό���(�ճǶ���H�C����J
�+�|(>����|�J���I#6�M�~s{DY�����wQ�H]���:H�cP�4hD�$�%pأ������amX�|��+_1���W�b������b��BF�\]AK�O#;��X-F۪�}N�|�"��Rz�"�E)��A�	c��İ�1e�"I�=��-�T�j9B#ǨrREG�l�a덦. �A��sQČ�X��#Q��"�:j����3���UfJ�J4��OV5:Z���t���iW���Wߟ�$l�!��@��5��҇4ۃ!Ͷ����f�Z��P����0x��#a��G<���0x��#t{���������2^W�?z$�?�lJTD�)���a�R�ѐ��~^Y�ψJ��q�T2��pHP�8���|���f�@o�L�1>�H��ę�t̵$�^�5˦��g_]_'���[����7#�ƭ�O���Ɨ3g��u0D��Xoy�Lh_g�wx���ĩ&u]��&C�� ���B;"]RGy����PK
   %��X�M��i  �;                  cirkitFile.jsonPK
   ���X`�/��1  �P  /             �i  images/05f650cb-cb4a-4256-a168-b327b67eb2f6.pngPK
   ���XG�~��  � /             �  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK
   ���XWC��)�  � /             �\ images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   ���Xw�'<�  �  /             .1 images/0ac982bd-8891-43e7-be61-3976077ece17.pngPK
   ���Xyɜ��  �  /             
N images/110f4c69-ce42-4daf-8800-65b9db14e3fe.pngPK
   0��X�r��}� �� /             �j images/1235872f-9927-4bec-a0e7-84fb82154d9a.pngPK
   ���X�䓶� � /             �R images/132fbcdf-34e4-44dc-827d-09a965026955.pngPK
   ���X��g  n  /             �
 images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK
   ���X����  �  /             n
 images/25cd0dd7-bebf-4a92-94a8-2c258b16bf7a.pngPK
   ���XhT���� ċ /             �7
 images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK
   ���X��НR5 �� /             �� images/52cc771c-8bcb-4758-820d-da79c3626c72.pngPK
   ���XT��"  T$  /             : images/53cc934f-9b11-4097-8823-694d19808ece.pngPK
   ���X��_8
  3
  /             �< images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   0��X��I� �� /             G images/60733dc7-8aae-4c8d-a308-d0d87ce42cc9.pngPK
   ���X�,Y�/  �/  /             �� images/6adb3134-3cc2-4380-b4ac-017fb4b87c19.pngPK
   ���X
=)�.� � /             � images/770fe9cc-a3ef-41fb-abe5-14f6fd7b0eeb.pngPK
   ���Xd��  �   /             � images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   ���X�IM��  � /             4� images/86917e2b-5e70-481a-b4c7-aed39e2d087b.pngPK
   ���X�1.:�  )  /             �� images/8d2526ea-6e7a-4b7c-a99b-0902daeefaab.pngPK
   ���X�Ƚ׌  �  /             �� images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK
   ���X?S��� 2� /             � images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   ���X	��#u } /             c� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   ���X$�8�l  �  /             �> images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   ���X+L$��� �� /             �\ images/aad47697-5cf4-402f-a095-abba84463b41.pngPK
   ���X����<  �  /             �.! images/bdd7c0cc-86d6-4eb9-abef-3fcf444ec41a.pngPK
   ���X���7z  �  /             7M! images/be8de2bb-09ef-440a-a2d8-19619bf9d0dd.pngPK
   ���Xp>r�  �  /             �h! images/c13bb491-011f-4ad1-adfa-58d33d2d83a5.pngPK
   ���X�GDU7� �� /             7�! images/d628d844-ce42-4e82-be63-f5fdfa438334.pngPK
   ���X������  ��  /             �j$ images/e758c5b4-10e9-4263-8b5b-5233ba63df2c.pngPK
   ���X��6�B  �  /             �1% images/ea05fd3c-afe5-4b36-b101-0986c4cae35e.pngPK
   ���X��@�/  �/  /             O7% images/ee535837-a8e5-4cdb-98a7-fed99fa44d94.pngPK
   ���X�T�|  �  /             0g% images/f1ab8fe3-f826-4bea-bba4-7763291602bf.pngPK
   ���XF���?� Q� /             �~% images/f590943e-678c-44eb-a174-3243ba5f3820.pngPK
   ���X�$&VAS }d /             ) images/f915906d-fb0f-4209-a242-05d71b94b060.pngPK
   %��X�"�Q  �               �c* jsons/user_defined.jsonPK    $ $ �  -v*   